* NGSPICE file created from sb_2__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxbp_1 abstract view
.subckt sky130_fd_sc_hd__dfxbp_1 D Q Q_N CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

.subckt sb_2__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11]
+ chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16]
+ chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_left_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11]
+ chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16]
+ chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2]
+ chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7]
+ chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11]
+ chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16]
+ chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] chany_top_out[9] left_bottom_grid_pin_1_ left_top_grid_pin_42_
+ left_top_grid_pin_43_ left_top_grid_pin_44_ left_top_grid_pin_45_ left_top_grid_pin_46_
+ left_top_grid_pin_47_ left_top_grid_pin_48_ left_top_grid_pin_49_ prog_clk top_left_grid_pin_34_
+ top_left_grid_pin_35_ top_left_grid_pin_36_ top_left_grid_pin_37_ top_left_grid_pin_38_
+ top_left_grid_pin_39_ top_left_grid_pin_40_ top_left_grid_pin_41_ top_right_grid_pin_1_
+ VPWR VGND
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_38.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_36.mux_l2_in_0__A0 _050_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 top_left_grid_pin_36_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_062_ _062_/HI _062_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_28.mux_l2_in_0__A1 mux_top_track_28.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.mux_l1_in_0__S mux_left_track_7.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_36.mux_l2_in_0__A1 mux_top_track_36.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A mux_left_track_1.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_34_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_061_ _061_/HI _061_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_30.mux_l2_in_0__S mux_top_track_30.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l2_in_0_/X _083_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.mux_l2_in_0_ _036_/HI mux_top_track_10.mux_l1_in_0_/X mux_top_track_10.mux_l2_in_0_/S
+ mux_top_track_10.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A mux_left_track_23.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_12.mux_l1_in_0_/S mux_top_track_12.mux_l2_in_0_/S
+ mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A mux_top_track_20.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l2_in_0_/X _075_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_21.mux_l1_in_0__S mux_left_track_21.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0__A0 _036_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_19.sky130_fd_sc_hd__buf_4_0_ mux_left_track_19.mux_l2_in_0_/X _078_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ mux_left_track_7.mux_l3_in_0_/S mux_left_track_7.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_060_ _060_/HI _060_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0__S mux_top_track_16.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_7.mux_l2_in_1_ _067_/HI left_top_grid_pin_49_ mux_left_track_7.mux_l2_in_0_/S
+ mux_left_track_7.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A mux_left_track_7.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_10.mux_l2_in_0_/S mux_top_track_12.mux_l1_in_0_/S
+ mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_13.mux_l2_in_0__S mux_left_track_13.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_10.mux_l1_in_0_ chanx_left_in[15] top_left_grid_pin_35_ mux_top_track_10.mux_l1_in_0_/S
+ mux_top_track_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 top_left_grid_pin_41_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_42_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_22.mux_l2_in_0_ _043_/HI mux_top_track_22.mux_l1_in_0_/X mux_top_track_22.mux_l2_in_0_/S
+ mux_top_track_22.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0__A1 mux_top_track_10.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A mux_top_track_0.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_15.mux_l2_in_0_ _058_/HI mux_left_track_15.mux_l1_in_0_/X mux_left_track_15.mux_l2_in_0_/S
+ mux_left_track_15.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_18.mux_l1_in_0_/S mux_top_track_18.mux_l2_in_0_/S
+ mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_2.mux_l2_in_0__A0 mux_top_track_2.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_26.sky130_fd_sc_hd__buf_4_0__A mux_top_track_26.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l2_in_0__S mux_top_track_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ mux_left_track_7.mux_l2_in_0_/S mux_left_track_7.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__072__A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_20.mux_l1_in_0__S mux_top_track_20.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_7.mux_l1_in_1_ left_top_grid_pin_47_ left_top_grid_pin_45_ mux_left_track_7.mux_l1_in_0_/S
+ mux_left_track_7.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_7.mux_l2_in_1__S mux_left_track_7.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l2_in_1_ _035_/HI mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 left_top_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0__A0 _056_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 top_left_grid_pin_39_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_22.sky130_fd_sc_hd__buf_4_0_ mux_top_track_22.mux_l2_in_0_/X _096_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__080__A _080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_2_ chanx_left_in[0] top_right_grid_pin_1_ mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0__A1 mux_top_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 mux_left_track_1.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_16.mux_l2_in_0_/S mux_top_track_18.mux_l1_in_0_/S
+ mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l2_in_0_/X _099_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmux_top_track_22.mux_l1_in_0_ chanx_left_in[9] top_left_grid_pin_41_ mux_top_track_22.mux_l1_in_0_/S
+ mux_top_track_22.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__075__A _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_34.mux_l2_in_0_ _049_/HI mux_top_track_34.mux_l1_in_0_/X mux_top_track_34.mux_l2_in_0_/S
+ mux_top_track_34.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_15.mux_l1_in_0_ left_top_grid_pin_45_ chany_top_in[13] mux_left_track_15.mux_l1_in_0_/S
+ mux_left_track_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A mux_top_track_6.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_27.mux_l2_in_0_ _064_/HI mux_left_track_27.mux_l1_in_0_/X ccff_tail
+ mux_left_track_27.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_30.mux_l1_in_0_/S mux_top_track_30.mux_l2_in_0_/S
+ mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_12.mux_l2_in_0__S mux_top_track_12.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_23.mux_l1_in_0_/S mux_left_track_23.mux_l2_in_0_/S
+ mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_7.mux_l1_in_0_ left_top_grid_pin_43_ chany_top_in[17] mux_left_track_7.mux_l1_in_0_/S
+ mux_left_track_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__083__A _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l3_in_0_/X _107_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 left_top_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0__A1 mux_left_track_11.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__078__A _078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_22.mux_l1_in_0__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l1_in_1_ top_left_grid_pin_40_ top_left_grid_pin_38_ mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0__A1 top_left_grid_pin_37_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__091__A _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_0__A0 top_left_grid_pin_37_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_38.sky130_fd_sc_hd__buf_4_0_ mux_top_track_38.mux_l2_in_0_/X _088_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__086__A _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_28.mux_l2_in_0_/S mux_top_track_30.mux_l1_in_0_/S
+ mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_2.mux_l2_in_0__S mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_21.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1__S mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_34.mux_l1_in_0_ chanx_left_in[3] top_left_grid_pin_39_ mux_top_track_34.mux_l1_in_0_/S
+ mux_top_track_34.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_21.mux_l2_in_0_/S mux_left_track_23.mux_l1_in_0_/S
+ mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_27.mux_l1_in_0_ left_top_grid_pin_43_ chany_top_in[7] mux_left_track_27.mux_l1_in_0_/S
+ mux_left_track_27.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_30.mux_l1_in_0__A0 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A0 _052_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_36.mux_l1_in_0_/S mux_top_track_36.mux_l2_in_0_/S
+ mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__094__A _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_22.mux_l1_in_0__A1 top_left_grid_pin_41_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l2_in_1__S mux_left_track_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0__A0 left_top_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_38.mux_l1_in_0__S mux_top_track_38.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A0 mux_top_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__089__A _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_36_ top_left_grid_pin_34_ mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0__A1 top_left_grid_pin_35_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 left_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_099_ _099_/A chany_top_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 top_right_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__097__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A mux_left_track_15.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A mux_top_track_12.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l3_in_0_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_30.mux_l1_in_0__A1 top_left_grid_pin_37_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_4.mux_l2_in_1__A1 mux_top_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 _065_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_34.mux_l2_in_0_/S mux_top_track_36.mux_l1_in_0_/S
+ mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_23.mux_l1_in_0__A0 left_top_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0__A1 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A1 mux_top_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l3_in_0__A0 mux_left_track_3.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A0 _039_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_27.mux_l2_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_098_ _098_/A chany_top_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_1__A0 _044_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_3.mux_l2_in_0_/S mux_left_track_3.mux_l3_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_0.mux_l1_in_1_/S mux_top_track_0.mux_l2_in_0_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_4.mux_l1_in_1__S mux_top_track_4.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 left_top_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_23.mux_l1_in_0__A1 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X _085_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 mux_top_track_24.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1__A0 _054_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A1 mux_left_track_3.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A mux_top_track_18.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l3_in_0_/S
+ mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_16.mux_l2_in_0__A1 mux_top_track_16.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 mux_top_track_8.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_34.mux_l1_in_0__S mux_top_track_34.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_21.sky130_fd_sc_hd__buf_4_0_ mux_left_track_21.mux_l2_in_0_/X _077_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_left_track_5.mux_l1_in_2__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_097_ _097_/A chany_top_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_15.sky130_fd_sc_hd__buf_4_0_ mux_left_track_15.mux_l2_in_0_/X _080_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_3.mux_l1_in_0_/S mux_left_track_3.mux_l2_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_32.mux_l2_in_0__A0 _048_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ ccff_head mux_top_track_0.mux_l1_in_1_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1__A1 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.mux_l1_in_1__A0 left_top_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 _059_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_6.mux_l1_in_0_/S mux_top_track_6.mux_l2_in_0_/S
+ mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_3.mux_l2_in_1_ _065_/HI left_top_grid_pin_49_ mux_left_track_3.mux_l2_in_0_/S
+ mux_left_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_26.mux_l2_in_0__S mux_top_track_26.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0__A0 mux_left_track_7.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__100__A _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_22.mux_l1_in_0_/S mux_top_track_22.mux_l2_in_0_/S
+ mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A mux_top_track_30.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_096_ _096_/A chany_top_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 _063_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l2_in_0_ _039_/HI mux_top_track_16.mux_l1_in_0_/X mux_top_track_16.mux_l2_in_0_/S
+ mux_top_track_16.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_15.mux_l1_in_0_/S mux_left_track_15.mux_l2_in_0_/S
+ mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_23.mux_l2_in_0__S mux_left_track_23.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_1.mux_l3_in_0_/S mux_left_track_3.mux_l1_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_079_ _079_/A chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_32.mux_l2_in_0__A1 mux_top_track_32.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_11.mux_l2_in_0_ _056_/HI mux_left_track_11.mux_l1_in_0_/X mux_left_track_11.mux_l2_in_0_/S
+ mux_left_track_11.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 mux_left_track_25.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1__S mux_top_track_0.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.mux_l1_in_1__A1 left_top_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A1 mux_left_track_17.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_28.mux_l1_in_0__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_4.mux_l3_in_0_/S mux_top_track_6.mux_l1_in_0_/S
+ mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_0_/S mux_left_track_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_7.mux_l2_in_0__A1 mux_left_track_7.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_20.mux_l2_in_0_/S mux_top_track_22.mux_l1_in_0_/S
+ mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l1_in_1_ left_top_grid_pin_47_ left_top_grid_pin_45_ mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_095_ _095_/A chany_top_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_30.mux_l1_in_0__S mux_top_track_30.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 left_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_13.mux_l2_in_0_/S mux_left_track_15.mux_l1_in_0_/S
+ mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_1.mux_l1_in_2__S mux_left_track_1.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__106__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_078_ _078_/A chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_12.sky130_fd_sc_hd__buf_4_0_ mux_top_track_12.mux_l2_in_0_/X _101_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_28.mux_l1_in_0_/S mux_top_track_28.mux_l2_in_0_/S
+ mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A mux_top_track_36.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l1_in_0_ chanx_left_in[12] top_left_grid_pin_38_ mux_top_track_16.mux_l1_in_0_/S
+ mux_top_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_36.mux_l1_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_28.mux_l2_in_0_ _046_/HI mux_top_track_28.mux_l1_in_0_/X mux_top_track_28.mux_l2_in_0_/S
+ mux_top_track_28.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_30.mux_l2_in_0_ _047_/HI mux_top_track_30.mux_l1_in_0_/X mux_top_track_30.mux_l2_in_0_/S
+ mux_top_track_30.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_7.mux_l3_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_11.mux_l1_in_0_ left_top_grid_pin_43_ chany_top_in[15] mux_left_track_11.mux_l1_in_0_/S
+ mux_left_track_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_28.mux_l1_in_0__A1 top_left_grid_pin_36_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_23.mux_l2_in_0_ _062_/HI mux_left_track_23.mux_l1_in_0_/X mux_left_track_23.mux_l2_in_0_/S
+ mux_left_track_23.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_22.mux_l2_in_0__S mux_top_track_22.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_0_ left_top_grid_pin_43_ chany_top_in[19] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_094_ _094_/A chany_top_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0__S mux_top_track_16.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ mux_top_track_6.mux_l3_in_0_/S mux_top_track_6.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_26.mux_l2_in_0_/S mux_top_track_28.mux_l1_in_0_/S
+ mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_1_ _053_/HI chanx_left_in[17] mux_top_track_6.mux_l2_in_0_/S
+ mux_top_track_6.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_36.mux_l1_in_0__A1 top_left_grid_pin_40_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_34.sky130_fd_sc_hd__buf_4_0_ mux_top_track_34.mux_l2_in_0_/X _090_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_25.mux_l1_in_1__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0__S mux_left_track_13.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_28.mux_l1_in_0_ chanx_left_in[6] top_left_grid_pin_36_ mux_top_track_28.mux_l1_in_0_/S
+ mux_top_track_28.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_28.sky130_fd_sc_hd__buf_4_0_ mux_top_track_28.mux_l2_in_0_/X _093_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_30.mux_l1_in_0_ chanx_left_in[5] top_left_grid_pin_37_ mux_top_track_30.mux_l1_in_0_/S
+ mux_top_track_30.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_7.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_23.mux_l1_in_0_ left_top_grid_pin_49_ chany_top_in[9] mux_left_track_23.mux_l1_in_0_/S
+ mux_left_track_23.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_6.mux_l1_in_0__S mux_top_track_6.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_093_ _093_/A chany_top_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_076_ _076_/A chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_059_ _059_/HI _059_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_6.sky130_fd_sc_hd__buf_4_0_ mux_top_track_6.mux_l3_in_0_/X _104_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_left_track_7.mux_l1_in_1__S mux_left_track_7.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_1_ top_left_grid_pin_41_ top_left_grid_pin_39_ mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_4.mux_l3_in_0__S mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_092_ _092_/A chany_top_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A mux_left_track_3.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_1__S mux_top_track_24.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_075_ _075_/A chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_12.mux_l1_in_0__S mux_top_track_12.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0__A1 top_left_grid_pin_35_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_38.mux_l2_in_0__A0 _051_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_058_ _058_/HI _058_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 top_left_grid_pin_37_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_6.mux_l1_in_0_ top_left_grid_pin_37_ top_left_grid_pin_35_ mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A mux_left_track_25.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_14.mux_l1_in_0_/S mux_top_track_14.mux_l2_in_0_/S
+ mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A mux_top_track_22.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X _087_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 _035_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_091_ _091_/A chany_top_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_7.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_11.mux_l1_in_0__A0 left_top_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_074_ _074_/A chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l3_in_0__A0 mux_top_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_19.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_38.mux_l2_in_0__A1 mux_top_track_38.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_057_ _057_/HI _057_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 top_left_grid_pin_35_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 left_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A mux_left_track_9.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_11.sky130_fd_sc_hd__buf_4_0_ mux_left_track_11.mux_l2_in_0_/X _082_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA__070__A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A1 top_right_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_12.mux_l2_in_0_/S mux_top_track_14.mux_l1_in_0_/S
+ mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_3.mux_l1_in_1__S mux_left_track_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_0.mux_l3_in_0__S mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_0.mux_l2_in_1__A1 mux_top_track_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_6.mux_l2_in_1__S mux_top_track_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_090_ _090_/A chany_top_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A mux_top_track_2.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_073_ chany_top_in[6] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_11.mux_l1_in_0__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_28.sky130_fd_sc_hd__buf_4_0__A mux_top_track_28.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A1 mux_top_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_12.mux_l2_in_0__A0 _037_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__073__A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_38.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_056_ _056_/HI _056_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__068__A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_36.mux_l2_in_0__S mux_top_track_36.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_12.mux_l2_in_0_ _037_/HI mux_top_track_12.mux_l1_in_0_/X mux_top_track_12.mux_l2_in_0_/S
+ mux_top_track_12.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__081__A _081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__076__A _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_20.mux_l2_in_0__A0 _042_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_27.sky130_fd_sc_hd__buf_4_0_ mux_left_track_27.mux_l2_in_0_/X _074_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 top_left_grid_pin_40_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_27.mux_l1_in_0__S mux_left_track_27.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_072_ chany_top_in[5] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_12.mux_l2_in_0__A1 mux_top_track_12.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 mux_top_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A mux_top_track_8.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_32.mux_l1_in_0_/S mux_top_track_32.mux_l2_in_0_/S
+ mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__084__A _084_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_107_ _107_/A chany_top_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA__079__A _079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_25.mux_l1_in_0_/S mux_left_track_25.mux_l2_in_0_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_19.mux_l2_in_0__S mux_left_track_19.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__092__A _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_20.mux_l2_in_0__A1 mux_top_track_20.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_12.mux_l1_in_0_ chanx_left_in[14] top_left_grid_pin_36_ mux_top_track_12.mux_l1_in_0_/S
+ mux_top_track_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 top_left_grid_pin_38_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 left_top_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_13.mux_l2_in_0__A0 _057_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__087__A _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_071_ chany_top_in[4] chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_2.mux_l2_in_1__S mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_23.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A mux_left_track_11.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_0_ _059_/HI mux_left_track_17.mux_l1_in_0_/X mux_left_track_17.mux_l2_in_0_/S
+ mux_left_track_17.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 mux_left_track_3.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l1_in_1_ _044_/HI chanx_left_in[8] mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_30.mux_l2_in_0_/S mux_top_track_32.mux_l1_in_0_/S
+ mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_106_ _106_/A chany_top_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__095__A _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_23.mux_l2_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_32.mux_l2_in_0__S mux_top_track_32.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_38.mux_l1_in_0_/S mux_top_track_38.mux_l2_in_0_/S
+ mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_26.mux_l1_in_0__S mux_top_track_26.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l1_in_1_ _034_/HI left_bottom_grid_pin_1_ mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_21.mux_l2_in_0__A0 _061_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.mux_l3_in_0__S mux_left_track_7.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_30.sky130_fd_sc_hd__buf_4_0_ mux_top_track_30.mux_l2_in_0_/X _092_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_2.mux_l2_in_1_ _041_/HI chanx_left_in[19] mux_top_track_2.mux_l2_in_0_/S
+ mux_top_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 left_top_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_13.mux_l2_in_0__A1 mux_left_track_13.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_070_ chany_top_in[3] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 top_right_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X _095_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__098__A _098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_23.mux_l1_in_0__S mux_left_track_23.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A1 mux_left_track_3.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 top_left_grid_pin_38_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l1_in_0_ top_right_grid_pin_1_ top_left_grid_pin_34_ mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_36.mux_l2_in_0_ _050_/HI mux_top_track_36.mux_l1_in_0_/X mux_top_track_36.mux_l2_in_0_/S
+ mux_top_track_36.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_18.sky130_fd_sc_hd__buf_4_0_ mux_top_track_18.mux_l2_in_0_/X _098_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_105_ _105_/A chany_top_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_17.mux_l1_in_0_ left_top_grid_pin_46_ chany_top_in[12] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 top_right_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A mux_left_track_17.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l2_in_0__S mux_top_track_18.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A mux_top_track_14.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l3_in_0_/S
+ mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_36.mux_l2_in_0_/S mux_top_track_38.mux_l1_in_0_/S
+ mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_9.mux_l1_in_0_ left_top_grid_pin_42_ chany_top_in[16] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_21.mux_l2_in_0__A1 mux_left_track_21.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_32.mux_l1_in_0__A0 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X _106_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_6.mux_l2_in_1__A0 _053_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_34_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_15.mux_l2_in_0__S mux_left_track_15.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l1_in_1_ top_left_grid_pin_41_ top_left_grid_pin_39_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 left_top_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__A0 mux_top_track_6.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_6.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_4.mux_l1_in_2__S mux_top_track_4.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_104_ _104_/A chany_top_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_7.mux_l1_in_0__A0 left_top_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_34_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l3_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_2.mux_l1_in_1_/S mux_top_track_2.mux_l2_in_0_/S
+ mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_36.mux_l1_in_0_ chanx_left_in[2] top_left_grid_pin_40_ mux_top_track_36.mux_l1_in_0_/S
+ mux_top_track_36.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_32.mux_l1_in_0__A1 top_left_grid_pin_38_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l2_in_1__A1 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 _066_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l1_in_0__S mux_top_track_22.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 left_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__S mux_left_track_3.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_11.mux_l1_in_0_/S mux_left_track_11.mux_l2_in_0_/S
+ mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_37_ top_left_grid_pin_35_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__A1 mux_top_track_6.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l2_in_0__A0 _040_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A0 mux_left_track_5.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_103_ _103_/A chany_top_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_034_ _034_/HI _034_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_7.mux_l1_in_0__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_15.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_5.mux_l1_in_0_/S mux_left_track_5.mux_l2_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_0.mux_l3_in_0_/S mux_top_track_2.mux_l1_in_1_/S
+ mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 left_top_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l2_in_0__S mux_top_track_14.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 mux_left_track_5.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__101__A _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_8.mux_l1_in_0_/S mux_top_track_8.mux_l2_in_0_/S
+ mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_26.mux_l2_in_0__A0 _045_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_9.mux_l2_in_0_/S mux_left_track_11.mux_l1_in_0_/S
+ mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_24.mux_l1_in_0_/S mux_top_track_24.mux_l2_in_0_/S
+ mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_18.mux_l2_in_0__A1 mux_top_track_18.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A1 mux_left_track_5.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A mux_top_track_32.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0__S mux_left_track_11.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_102_ _102_/A chany_top_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_17.mux_l1_in_0_/S mux_left_track_17.mux_l2_in_0_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_3.mux_l3_in_0_/S mux_left_track_5.mux_l1_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_6.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__104__A _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2__S mux_top_track_0.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_34.mux_l2_in_0__A0 _049_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_6.mux_l3_in_0_/S mux_top_track_8.mux_l1_in_0_/S
+ mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_26.mux_l2_in_0__A1 mux_top_track_26.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_7.sky130_fd_sc_hd__buf_4_0_ mux_left_track_7.mux_l3_in_0_/X _084_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_19.mux_l2_in_0__A0 _060_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l1_in_1__A0 _034_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_22.mux_l2_in_0_/S mux_top_track_24.mux_l1_in_0_/S
+ mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_25.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__107__A _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 mux_left_track_9.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ _101_/A chany_top_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_15.mux_l2_in_0_/S mux_left_track_17.mux_l1_in_0_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_23.sky130_fd_sc_hd__buf_4_0_ mux_left_track_23.mux_l2_in_0_/X _076_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A mux_top_track_38.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l2_in_0_/X _079_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_34.mux_l2_in_0__A1 mux_top_track_34.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_27.mux_l2_in_0__A0 _064_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_10.mux_l2_in_0__S mux_top_track_10.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_19.mux_l2_in_0__A1 mux_left_track_19.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l1_in_1__A1 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_36.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l2_in_1_ _066_/HI mux_left_track_5.mux_l1_in_2_/X mux_left_track_5.mux_l2_in_0_/S
+ mux_left_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_19.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_100_ _100_/A chany_top_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_2_ left_bottom_grid_pin_1_ left_top_grid_pin_48_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_18.mux_l2_in_0_ _040_/HI mux_top_track_18.mux_l1_in_0_/X mux_top_track_18.mux_l2_in_0_/S
+ mux_top_track_18.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_20.mux_l2_in_0_ _042_/HI mux_top_track_20.mux_l1_in_0_/X mux_top_track_20.mux_l2_in_0_/S
+ mux_top_track_20.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_13.mux_l2_in_0_ _057_/HI mux_left_track_13.mux_l1_in_0_/X mux_left_track_13.mux_l2_in_0_/S
+ mux_left_track_13.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_27.mux_l2_in_0__A1 mux_left_track_27.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_38.mux_l1_in_0__A0 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_6.mux_l1_in_1__S mux_top_track_6.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_1_ left_top_grid_pin_46_ left_top_grid_pin_44_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_20.sky130_fd_sc_hd__buf_4_0_ mux_top_track_20.mux_l2_in_0_/X _097_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1__A0 top_left_grid_pin_40_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_36.mux_l1_in_0__S mux_top_track_36.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A mux_left_track_21.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_10.mux_l1_in_0_/S mux_top_track_10.mux_l2_in_0_/S
+ mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_14.sky130_fd_sc_hd__buf_4_0_ mux_top_track_14.mux_l2_in_0_/X _100_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 mux_top_track_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_18.mux_l1_in_0_ chanx_left_in[11] top_left_grid_pin_39_ mux_top_track_18.mux_l1_in_0_/S
+ mux_top_track_18.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_20.mux_l1_in_0_ chanx_left_in[10] top_left_grid_pin_40_ mux_top_track_20.mux_l1_in_0_/S
+ mux_top_track_20.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_38.mux_l1_in_0__A1 top_left_grid_pin_41_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l2_in_0_ _048_/HI mux_top_track_32.mux_l1_in_0_/X mux_top_track_32.mux_l2_in_0_/S
+ mux_top_track_32.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_13.mux_l1_in_0_ left_top_grid_pin_44_ chany_top_in[14] mux_left_track_13.mux_l1_in_0_/S
+ mux_left_track_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_28.mux_l2_in_0__S mux_top_track_28.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A mux_left_track_5.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_0_ left_top_grid_pin_42_ chany_top_in[18] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_089_ _089_/A chany_top_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_1_ _063_/HI left_bottom_grid_pin_1_ mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1__A1 top_left_grid_pin_38_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_8.mux_l2_in_0_/S mux_top_track_10.mux_l1_in_0_/S
+ mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l2_in_0__S mux_left_track_25.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_19.mux_l1_in_0__S mux_left_track_19.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A mux_left_track_27.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_36.sky130_fd_sc_hd__buf_4_0_ mux_top_track_36.mux_l2_in_0_/X _089_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_41_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_16.mux_l1_in_0_/S mux_top_track_16.mux_l2_in_0_/S
+ mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A mux_top_track_24.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l1_in_0_ chanx_left_in[4] top_left_grid_pin_38_ mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_21.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_0_ left_top_grid_pin_42_ chany_top_in[8] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_088_ _088_/A chany_top_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_20.mux_l1_in_0__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__071__A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_32.mux_l1_in_0__S mux_top_track_32.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_0_/S mux_top_track_8.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_12.mux_l1_in_0__A1 top_left_grid_pin_36_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_7.mux_l2_in_0__S mux_left_track_7.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 top_left_grid_pin_36_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_14.mux_l2_in_0_/S mux_top_track_16.mux_l1_in_0_/S
+ mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_top_track_8.mux_l1_in_1_ _054_/HI chanx_left_in[16] mux_top_track_8.mux_l1_in_0_/S
+ mux_top_track_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l2_in_0_/X _103_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A mux_top_track_4.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__074__A _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ _087_/A chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 _041_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__069__A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_21.mux_l1_in_0_/S mux_left_track_21.mux_l2_in_0_/S
+ mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_20.mux_l1_in_0__A1 top_left_grid_pin_40_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_13.mux_l1_in_0__A0 left_top_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_18.mux_l1_in_0__S mux_top_track_18.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A0 mux_top_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__082__A _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 left_top_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_34_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__077__A _077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l1_in_0_ top_right_grid_pin_1_ top_left_grid_pin_34_ mux_top_track_8.mux_l1_in_0_/S
+ mux_top_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_21.mux_l2_in_0__S mux_left_track_21.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A0 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_15.mux_l1_in_0__S mux_left_track_15.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__090__A _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_086_ _086_/A chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 _055_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X _086_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_21.mux_l1_in_0__A0 left_top_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__085__A _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_19.mux_l2_in_0_/S mux_left_track_21.mux_l1_in_0_/S
+ mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_069_ chany_top_in[2] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_34.mux_l1_in_0_/S mux_top_track_34.mux_l2_in_0_/S
+ mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0__A0 _038_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l3_in_0__A1 mux_top_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A0 mux_left_track_1.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_27.mux_l1_in_0_/S ccff_tail
+ mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__093__A _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0__S mux_left_track_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__088__A _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 left_top_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_13.sky130_fd_sc_hd__buf_4_0_ mux_left_track_13.mux_l2_in_0_/X _081_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__S mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_085_ _085_/A chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l2_in_1__A1 mux_left_track_1.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_21.mux_l1_in_0__A1 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A mux_left_track_13.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_22.mux_l2_in_0__A0 _043_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A mux_top_track_10.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_068_ chany_top_in[1] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_6.mux_l1_in_1__A0 top_left_grid_pin_41_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__096__A _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_32.mux_l2_in_0_/S mux_top_track_34.mux_l1_in_0_/S
+ mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_1.mux_l3_in_0__A1 mux_left_track_1.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l2_in_0__A1 mux_top_track_14.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_20.mux_l2_in_0__S mux_top_track_20.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ _055_/HI mux_left_track_1.mux_l1_in_2_/X mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l2_in_0__A0 mux_top_track_6.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_14.mux_l1_in_0__S mux_top_track_14.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_25.mux_l2_in_0_/S mux_left_track_27.mux_l1_in_0_/S
+ mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l1_in_2_ left_bottom_grid_pin_1_ left_top_grid_pin_48_ mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_14.mux_l2_in_0_ _038_/HI mux_top_track_14.mux_l1_in_0_/X mux_top_track_14.mux_l2_in_0_/S
+ mux_top_track_14.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_3.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_30.mux_l2_in_0__A0 _047_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__099__A _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_084_ _084_/A chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_11.mux_l1_in_0__S mux_left_track_11.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l3_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_22.mux_l2_in_0__A1 mux_top_track_22.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_067_ _067_/HI _067_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_15.mux_l2_in_0__A0 _058_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 left_top_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_1__A1 top_left_grid_pin_39_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A mux_left_track_19.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l2_in_0__A1 mux_top_track_6.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 mux_left_track_5.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A mux_top_track_16.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_4.mux_l2_in_0_/S mux_top_track_4.mux_l3_in_0_/S
+ mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_1_ left_top_grid_pin_46_ left_top_grid_pin_44_ mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_10.sky130_fd_sc_hd__buf_4_0_ mux_top_track_10.mux_l2_in_0_/X _102_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_30.mux_l2_in_0__A1 mux_top_track_30.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_083_ _083_/A chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_23.mux_l2_in_0__A0 _062_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_1__S mux_left_track_5.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_23.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_1.mux_l1_in_0_/S mux_left_track_1.mux_l2_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_14.mux_l1_in_0_ chanx_left_in[13] top_left_grid_pin_37_ mux_top_track_14.mux_l1_in_0_/S
+ mux_top_track_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_26.mux_l2_in_0_ _045_/HI mux_top_track_26.mux_l1_in_0_/X mux_top_track_26.mux_l2_in_0_/S
+ mux_top_track_26.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l3_in_0__S mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_066_ _066_/HI _066_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_15.mux_l2_in_0__A1 mux_left_track_15.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 left_top_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_26.mux_l1_in_0__A0 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_19.mux_l2_in_0_ _060_/HI mux_left_track_19.mux_l1_in_0_/X mux_left_track_19.mux_l2_in_0_/S
+ mux_left_track_19.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_18.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_21.mux_l2_in_0_ _061_/HI mux_left_track_21.mux_l1_in_0_/X mux_left_track_21.mux_l2_in_0_/S
+ mux_left_track_21.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_7.mux_l2_in_0_/S mux_left_track_7.mux_l3_in_0_/S
+ mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A1 top_left_grid_pin_39_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_4.mux_l1_in_2_/S mux_top_track_4.mux_l2_in_0_/S
+ mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.mux_l1_in_0_ left_top_grid_pin_42_ chany_top_in[0] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0__S mux_top_track_10.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_38.mux_l2_in_0__S mux_top_track_38.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_20.mux_l1_in_0_/S mux_top_track_20.mux_l2_in_0_/S
+ mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_34.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_082_ _082_/A chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_23.mux_l2_in_0__A1 mux_left_track_23.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_13.mux_l1_in_0_/S mux_left_track_13.mux_l2_in_0_/S
+ mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_top_track_4.mux_l2_in_1_ _052_/HI mux_top_track_4.mux_l1_in_2_/X mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l2_in_0_/X _091_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_34.mux_l1_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_38.mux_l2_in_0_/S mux_left_track_1.mux_l1_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_065_ _065_/HI _065_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_26.mux_l1_in_0__A1 top_left_grid_pin_35_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_2_ chanx_left_in[18] top_right_grid_pin_1_ mux_top_track_4.mux_l1_in_2_/S
+ mux_top_track_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_26.sky130_fd_sc_hd__buf_4_0_ mux_top_track_26.mux_l2_in_0_/X _094_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_19.mux_l1_in_0__A0 left_top_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_26.mux_l1_in_0_ chanx_left_in[7] top_left_grid_pin_35_ mux_top_track_26.mux_l1_in_0_/S
+ mux_top_track_26.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_7.mux_l1_in_0_/S mux_left_track_7.mux_l2_in_0_/S
+ mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_38.mux_l2_in_0_ _051_/HI mux_top_track_38.mux_l1_in_0_/X mux_top_track_38.mux_l2_in_0_/S
+ mux_top_track_38.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_2.mux_l3_in_0_/S mux_top_track_4.mux_l1_in_2_/S
+ mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_19.mux_l1_in_0_ left_top_grid_pin_47_ chany_top_in[11] mux_left_track_19.mux_l1_in_0_/S
+ mux_left_track_19.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 left_top_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__102__A _102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_21.mux_l1_in_0_ left_top_grid_pin_48_ chany_top_in[10] mux_left_track_21.mux_l1_in_0_/S
+ mux_left_track_21.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_18.mux_l2_in_0_/S mux_top_track_20.mux_l1_in_0_/S
+ mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_081_ _081_/A chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_11.mux_l2_in_0_/S mux_left_track_13.mux_l1_in_0_/S
+ mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_0_/S mux_top_track_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_34.mux_l1_in_0__A1 top_left_grid_pin_39_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.mux_l2_in_1__A0 _067_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X _105_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
X_064_ _064_/HI _064_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_27.mux_l1_in_0__A0 left_top_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_26.mux_l1_in_0_/S mux_top_track_26.mux_l2_in_0_/S
+ mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A mux_top_track_34.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_40_ top_left_grid_pin_38_ mux_top_track_4.mux_l1_in_2_/S
+ mux_top_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_19.mux_l1_in_0__A1 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_19.mux_l1_in_0_/S mux_left_track_19.mux_l2_in_0_/S
+ mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_7.mux_l3_in_0__A0 mux_left_track_7.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_5.mux_l3_in_0_/S mux_left_track_7.mux_l1_in_0_/S
+ mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_4.mux_l2_in_1__S mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_38.mux_l1_in_0_ chanx_left_in[1] top_left_grid_pin_41_ mux_top_track_38.mux_l1_in_0_/S
+ mux_top_track_38.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_080_ _080_/A chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_27.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_34.mux_l2_in_0__S mux_top_track_34.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_7.mux_l2_in_1__A1 left_top_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_28.mux_l1_in_0__S mux_top_track_28.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_063_ _063_/HI _063_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_27.mux_l1_in_0__A1 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_24.mux_l2_in_0_/S mux_top_track_26.mux_l1_in_0_/S
+ mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_28.mux_l2_in_0__A0 _046_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_36_ top_left_grid_pin_34_ mux_top_track_4.mux_l1_in_2_/S
+ mux_top_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_20.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_7.mux_l3_in_0__A1 mux_left_track_7.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_17.mux_l2_in_0_/S mux_left_track_19.mux_l1_in_0_/S
+ mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

