* NGSPICE file created from sb_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

.subckt sb_0__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_11_ bottom_left_grid_pin_13_ bottom_left_grid_pin_15_
+ bottom_left_grid_pin_1_ bottom_left_grid_pin_3_ bottom_left_grid_pin_5_ bottom_left_grid_pin_7_
+ bottom_left_grid_pin_9_ bottom_right_grid_pin_11_ chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ right_bottom_grid_pin_12_ right_top_grid_pin_10_ top_left_grid_pin_11_ top_left_grid_pin_13_
+ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_ top_left_grid_pin_5_
+ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_ vpwr vgnd
Xmem_right_track_12.LATCH_1_.latch data_in _067_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_148 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_56 vgnd vpwr scs8hd_decap_3
XFILLER_3_45 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _116_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_203 vgnd vpwr scs8hd_decap_12
XFILLER_10_103 vpwr vgnd scs8hd_fill_2
XFILLER_10_114 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _067_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_87 vgnd vpwr scs8hd_decap_4
XFILLER_33_206 vgnd vpwr scs8hd_decap_8
XANTENNA__108__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_195 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _146_/HI _062_/Y mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _140_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_75 vpwr vgnd scs8hd_fill_2
X_131_ _130_/A address[6] _111_/C _083_/C _131_/Y vgnd vpwr scs8hd_nor4_4
X_062_ _062_/A _062_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_198 vgnd vpwr scs8hd_fill_1
XANTENNA__110__C _095_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_35 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _097_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _165_/A vgnd vpwr scs8hd_inv_1
XFILLER_12_209 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_20 vgnd vpwr scs8hd_decap_8
XFILLER_18_64 vpwr vgnd scs8hd_fill_2
XFILLER_18_97 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
X_114_ _099_/A _116_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__121__B _121_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_7_ mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_139 vpwr vgnd scs8hd_fill_2
XFILLER_4_205 vgnd vpwr scs8hd_decap_8
XFILLER_20_21 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_161 vgnd vpwr scs8hd_decap_8
XANTENNA__116__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_23 vgnd vpwr scs8hd_fill_1
XANTENNA__132__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.LATCH_1_.latch data_in _069_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_25_131 vgnd vpwr scs8hd_fill_1
XFILLER_31_31 vgnd vpwr scs8hd_decap_12
XFILLER_15_54 vpwr vgnd scs8hd_fill_2
XFILLER_15_98 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _064_/A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_134 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_131 vgnd vpwr scs8hd_decap_4
XFILLER_16_142 vpwr vgnd scs8hd_fill_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _066_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _140_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_101 vgnd vpwr scs8hd_fill_1
Xmux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _143_/HI _068_/Y mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_64 vgnd vpwr scs8hd_decap_8
XFILLER_13_112 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _147_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_171 vgnd vpwr scs8hd_decap_8
XFILLER_27_226 vgnd vpwr scs8hd_decap_6
XFILLER_6_108 vgnd vpwr scs8hd_decap_12
XFILLER_10_137 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vpwr vgnd scs8hd_fill_2
XFILLER_5_174 vpwr vgnd scs8hd_fill_2
XANTENNA__124__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
X_130_ _130_/A address[6] _130_/C address[0] _130_/Y vgnd vpwr scs8hd_nor4_4
X_061_ _061_/A _061_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_34 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_113_ _098_/A _116_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _068_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _072_/A mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_88 vgnd vpwr scs8hd_decap_4
XFILLER_29_86 vpwr vgnd scs8hd_fill_2
XANTENNA__132__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_34_121 vgnd vpwr scs8hd_fill_1
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_198 vpwr vgnd scs8hd_fill_2
XFILLER_15_11 vpwr vgnd scs8hd_fill_2
XFILLER_31_76 vpwr vgnd scs8hd_fill_2
XFILLER_31_43 vgnd vpwr scs8hd_decap_12
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XFILLER_22_113 vgnd vpwr scs8hd_decap_8
XFILLER_30_190 vgnd vpwr scs8hd_fill_1
XFILLER_22_146 vpwr vgnd scs8hd_fill_2
XANTENNA__053__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _059_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_168 vgnd vpwr scs8hd_decap_3
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _066_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _161_/A vgnd vpwr scs8hd_inv_1
XFILLER_3_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__138__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_8_194 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_149 vgnd vpwr scs8hd_decap_4
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XFILLER_33_219 vpwr vgnd scs8hd_fill_2
XFILLER_5_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_230 vgnd vpwr scs8hd_decap_3
XFILLER_24_208 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_230 vgnd vpwr scs8hd_decap_3
XFILLER_23_88 vpwr vgnd scs8hd_fill_2
XFILLER_23_55 vpwr vgnd scs8hd_fill_2
XFILLER_23_33 vpwr vgnd scs8hd_fill_2
XFILLER_23_22 vpwr vgnd scs8hd_fill_2
X_060_ _060_/A _060_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XFILLER_2_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_167 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__135__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__061__A _061_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_76 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_211 vgnd vpwr scs8hd_decap_4
XFILLER_11_222 vpwr vgnd scs8hd_fill_2
X_112_ _097_/A _116_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _061_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__056__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_29_10 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _059_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_67 vgnd vpwr scs8hd_decap_4
XFILLER_20_78 vgnd vpwr scs8hd_decap_3
XFILLER_28_185 vgnd vpwr scs8hd_fill_1
XANTENNA__132__C _111_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_130 vgnd vpwr scs8hd_decap_3
XFILLER_19_163 vpwr vgnd scs8hd_fill_2
XFILLER_19_174 vpwr vgnd scs8hd_fill_2
XFILLER_34_188 vgnd vpwr scs8hd_decap_12
XFILLER_15_34 vpwr vgnd scs8hd_fill_2
XFILLER_31_99 vgnd vpwr scs8hd_decap_4
XFILLER_31_55 vgnd vpwr scs8hd_decap_6
XFILLER_0_221 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_158 vgnd vpwr scs8hd_decap_3
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _075_/C vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_169 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _061_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XFILLER_13_147 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _063_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_3_26 vpwr vgnd scs8hd_fill_2
XANTENNA__138__B _134_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_140 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__064__A _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_35 vgnd vpwr scs8hd_decap_3
XFILLER_12_57 vgnd vpwr scs8hd_decap_4
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_132 vgnd vpwr scs8hd_decap_6
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _086_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_80 vpwr vgnd scs8hd_fill_2
XANTENNA__059__A _059_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_135 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_14_231 vpwr vgnd scs8hd_fill_2
XANTENNA__135__C _096_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _065_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _145_/HI _060_/Y mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_18_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
X_111_ address[5] _134_/B _111_/C _116_/B vgnd vpwr scs8hd_or3_4
XFILLER_7_205 vgnd vpwr scs8hd_decap_3
XFILLER_7_227 vgnd vpwr scs8hd_decap_6
XANTENNA__162__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__072__A _072_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_13 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _148_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__132__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_15 vpwr vgnd scs8hd_fill_2
XFILLER_6_26 vpwr vgnd scs8hd_fill_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_6
XANTENNA__157__A _157_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_197 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _144_/HI _071_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _091_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_156 vpwr vgnd scs8hd_fill_2
XFILLER_25_134 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_68 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_112 vgnd vpwr scs8hd_decap_8
XFILLER_16_189 vgnd vpwr scs8hd_decap_8
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_126 vpwr vgnd scs8hd_fill_2
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__D _083_/C vgnd vpwr scs8hd_diode_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__C _130_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _062_/A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__170__A _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _084_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _142_/HI _066_/Y mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_199 vpwr vgnd scs8hd_fill_2
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_46 vpwr vgnd scs8hd_fill_2
XANTENNA__075__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_39 vgnd vpwr scs8hd_decap_4
XANTENNA__135__D _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_1_191 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _070_/Y mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_202 vpwr vgnd scs8hd_fill_2
XFILLER_20_224 vgnd vpwr scs8hd_decap_8
XFILLER_18_68 vgnd vpwr scs8hd_decap_3
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _056_/Y _057_/Y _095_/C _111_/C vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _065_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_49 vgnd vpwr scs8hd_decap_6
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XANTENNA__173__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _068_/A mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_25 vgnd vpwr scs8hd_decap_3
XFILLER_15_47 vgnd vpwr scs8hd_decap_4
XFILLER_15_58 vgnd vpwr scs8hd_decap_3
XANTENNA__083__A address[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_190 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_135 vgnd vpwr scs8hd_fill_1
XFILLER_16_146 vgnd vpwr scs8hd_decap_6
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_90 vgnd vpwr scs8hd_decap_4
XANTENNA__168__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_182 vgnd vpwr scs8hd_decap_8
XFILLER_7_92 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_35 vgnd vpwr scs8hd_decap_12
XFILLER_13_116 vgnd vpwr scs8hd_decap_4
XANTENNA__078__A _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_160 vgnd vpwr scs8hd_decap_4
XANTENNA__138__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__080__B _099_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_101 vpwr vgnd scs8hd_fill_2
XFILLER_5_178 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _067_/A vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _093_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_222 vgnd vpwr scs8hd_decap_8
XANTENNA__075__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_104 vpwr vgnd scs8hd_fill_2
XFILLER_3_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_38 vpwr vgnd scs8hd_fill_2
XFILLER_1_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _062_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__176__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_5_ mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_58 vgnd vpwr scs8hd_decap_4
XFILLER_34_68 vgnd vpwr scs8hd_decap_8
XANTENNA__086__A _084_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ _169_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_122 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_188 vgnd vpwr scs8hd_decap_4
XFILLER_19_144 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vgnd vpwr scs8hd_fill_1
XANTENNA__083__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_139 vpwr vgnd scs8hd_fill_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_169 vgnd vpwr scs8hd_decap_12
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _060_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__078__B _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_58 vgnd vpwr scs8hd_decap_4
XANTENNA__094__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_194 vpwr vgnd scs8hd_fill_2
XFILLER_3_18 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _064_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _154_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_231 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _099_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A _097_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _061_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_26 vgnd vpwr scs8hd_decap_4
XANTENNA__075__C _075_/C vgnd vpwr scs8hd_diode_2
XANTENNA__091__B _092_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_127 vpwr vgnd scs8hd_fill_2
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_9_17 vpwr vgnd scs8hd_fill_2
XFILLER_14_201 vgnd vpwr scs8hd_fill_1
XFILLER_13_81 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_6 vpwr vgnd scs8hd_fill_2
XANTENNA__086__B _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_219 vpwr vgnd scs8hd_fill_2
XFILLER_11_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _062_/A vgnd vpwr
+ scs8hd_diode_2
X_168_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_099_ _099_/A _102_/B _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_6
XFILLER_1_73 vpwr vgnd scs8hd_fill_2
XFILLER_1_84 vpwr vgnd scs8hd_fill_2
XFILLER_20_49 vgnd vpwr scs8hd_fill_1
XFILLER_29_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_14 vgnd vpwr scs8hd_decap_12
XFILLER_28_145 vpwr vgnd scs8hd_fill_2
XFILLER_28_112 vgnd vpwr scs8hd_fill_1
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_fill_1
XFILLER_34_126 vgnd vpwr scs8hd_decap_12
XFILLER_19_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_167 vpwr vgnd scs8hd_fill_2
XFILLER_19_178 vgnd vpwr scs8hd_decap_3
XANTENNA__083__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_225 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_1 vgnd vpwr scs8hd_decap_3
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _157_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__094__B _092_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _067_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_3
XFILLER_32_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_133 vgnd vpwr scs8hd_decap_4
XFILLER_8_144 vpwr vgnd scs8hd_fill_2
XFILLER_12_173 vgnd vpwr scs8hd_decap_12
XANTENNA__089__B _092_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_114 vgnd vpwr scs8hd_decap_6
XFILLER_4_84 vgnd vpwr scs8hd_decap_8
XFILLER_4_73 vgnd vpwr scs8hd_fill_1
XFILLER_4_51 vgnd vpwr scs8hd_decap_3
XFILLER_23_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _060_/A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
XFILLER_13_71 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_16 vpwr vgnd scs8hd_fill_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_24_81 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_098_ _098_/A _102_/B _098_/Y vgnd vpwr scs8hd_nor2_4
X_167_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_1_52 vgnd vpwr scs8hd_decap_3
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_26 vgnd vpwr scs8hd_decap_12
XFILLER_20_17 vpwr vgnd scs8hd_fill_2
XFILLER_28_179 vgnd vpwr scs8hd_decap_6
XFILLER_28_157 vpwr vgnd scs8hd_fill_2
XANTENNA__097__B _102_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _064_/Y mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_19 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_138 vgnd vpwr scs8hd_decap_12
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_33_182 vgnd vpwr scs8hd_fill_1
XFILLER_33_160 vgnd vpwr scs8hd_decap_8
XFILLER_25_138 vpwr vgnd scs8hd_fill_2
XFILLER_18_190 vpwr vgnd scs8hd_fill_2
XFILLER_0_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_138 vpwr vgnd scs8hd_fill_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _150_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_141 vgnd vpwr scs8hd_fill_1
XFILLER_7_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _068_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_152 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vgnd vpwr scs8hd_decap_8
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _066_/A mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_141 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XFILLER_26_200 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_23_214 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_94 vgnd vpwr scs8hd_decap_3
XFILLER_1_173 vgnd vpwr scs8hd_decap_8
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _072_/Y mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _066_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_28 vgnd vpwr scs8hd_fill_1
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_217 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_097_ _097_/A _102_/B _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_232 vgnd vpwr scs8hd_fill_1
X_166_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_38 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _072_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_169 vgnd vpwr scs8hd_fill_1
XFILLER_10_73 vpwr vgnd scs8hd_fill_2
XFILLER_19_60 vgnd vpwr scs8hd_fill_1
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_4
XFILLER_27_180 vgnd vpwr scs8hd_fill_1
XFILLER_19_93 vpwr vgnd scs8hd_fill_2
X_149_ _149_/HI _149_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_194 vgnd vpwr scs8hd_decap_4
XFILLER_24_183 vgnd vpwr scs8hd_decap_4
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_94 vgnd vpwr scs8hd_fill_1
XPHY_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _141_/HI mem_bottom_track_9.LATCH_2_.latch/Q
+ mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_17 vgnd vpwr scs8hd_decap_12
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_197 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _061_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _068_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_19 vpwr vgnd scs8hd_fill_2
XFILLER_26_212 vpwr vgnd scs8hd_fill_2
XFILLER_5_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_71 vgnd vpwr scs8hd_decap_6
XFILLER_17_201 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_152 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _059_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_1_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
X_165_ _165_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
X_096_ address[5] address[6] _096_/C _102_/B vgnd vpwr scs8hd_or3_4
XFILLER_1_32 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _084_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_104 vpwr vgnd scs8hd_fill_2
XFILLER_28_126 vgnd vpwr scs8hd_decap_8
XFILLER_3_203 vpwr vgnd scs8hd_fill_2
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_41 vgnd vpwr scs8hd_decap_8
XFILLER_10_52 vgnd vpwr scs8hd_decap_6
XFILLER_10_85 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _063_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_83 vgnd vpwr scs8hd_fill_1
XFILLER_19_126 vpwr vgnd scs8hd_fill_2
XFILLER_19_148 vpwr vgnd scs8hd_fill_2
X_148_ _148_/HI _148_/LO vgnd vpwr scs8hd_conb_1
X_079_ _081_/A address[2] _083_/C _099_/A vgnd vpwr scs8hd_or3_4
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_18_170 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vpwr vgnd scs8hd_fill_2
XFILLER_24_162 vpwr vgnd scs8hd_fill_2
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
XFILLER_21_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_165 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_173 vgnd vpwr scs8hd_decap_4
XFILLER_15_195 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XFILLER_26_29 vpwr vgnd scs8hd_fill_2
XFILLER_21_110 vpwr vgnd scs8hd_fill_2
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XFILLER_29_232 vgnd vpwr scs8hd_fill_1
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_187 vgnd vpwr scs8hd_fill_1
XFILLER_16_73 vpwr vgnd scs8hd_fill_2
XFILLER_16_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__103__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _065_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_76 vgnd vpwr scs8hd_fill_1
XFILLER_4_43 vgnd vpwr scs8hd_decap_8
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_0_.latch data_in _072_/A _138_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__100__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_164_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
X_095_ _056_/Y address[3] _095_/C _096_/C vgnd vpwr scs8hd_or3_4
XFILLER_6_212 vpwr vgnd scs8hd_fill_2
XFILLER_1_11 vgnd vpwr scs8hd_decap_12
XFILLER_1_77 vpwr vgnd scs8hd_fill_2
XFILLER_1_88 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_97 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_94 vgnd vpwr scs8hd_decap_12
XFILLER_35_83 vpwr vgnd scs8hd_fill_2
X_147_ _147_/HI _147_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__106__A _099_/A vgnd vpwr scs8hd_diode_2
X_078_ _084_/A _098_/A _078_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XFILLER_31_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_141 vgnd vpwr scs8hd_fill_1
XFILLER_30_133 vpwr vgnd scs8hd_fill_2
XFILLER_30_122 vgnd vpwr scs8hd_decap_8
XFILLER_7_32 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _062_/Y mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_148 vgnd vpwr scs8hd_decap_4
XFILLER_32_84 vgnd vpwr scs8hd_decap_4
XANTENNA__103__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_203 vpwr vgnd scs8hd_fill_2
XFILLER_32_206 vgnd vpwr scs8hd_decap_8
XFILLER_17_214 vpwr vgnd scs8hd_fill_2
XFILLER_17_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_195 vgnd vpwr scs8hd_fill_1
XANTENNA__114__A _099_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_31 vgnd vpwr scs8hd_fill_1
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_198 vpwr vgnd scs8hd_fill_2
XFILLER_1_187 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_85 vgnd vpwr scs8hd_fill_1
X_163_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_224 vgnd vpwr scs8hd_decap_8
X_094_ _102_/A _092_/B _094_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__111__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _151_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_45 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _092_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _067_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _068_/Y mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_172 vpwr vgnd scs8hd_fill_2
XFILLER_27_150 vpwr vgnd scs8hd_fill_2
XFILLER_19_52 vpwr vgnd scs8hd_fill_2
XANTENNA__122__A _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA__106__B _106_/B vgnd vpwr scs8hd_diode_2
X_077_ address[1] _077_/B address[0] _098_/A vgnd vpwr scs8hd_or3_4
X_146_ _146_/HI _146_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_6 vgnd vpwr scs8hd_decap_12
XFILLER_18_194 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_208 vgnd vpwr scs8hd_decap_8
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_86 vpwr vgnd scs8hd_fill_2
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_145 vgnd vpwr scs8hd_decap_8
XFILLER_7_88 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _102_/A vgnd vpwr scs8hd_diode_2
X_129_ _130_/A address[6] _130_/C _083_/C _129_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_156 vpwr vgnd scs8hd_fill_2
XFILLER_32_74 vgnd vpwr scs8hd_fill_1
XFILLER_32_30 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__103__C _096_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_215 vpwr vgnd scs8hd_fill_2
XFILLER_7_160 vpwr vgnd scs8hd_fill_2
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _142_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_204 vgnd vpwr scs8hd_fill_1
XFILLER_32_218 vgnd vpwr scs8hd_decap_12
XANTENNA__114__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_185 vpwr vgnd scs8hd_fill_2
XFILLER_4_174 vgnd vpwr scs8hd_decap_3
XFILLER_4_56 vpwr vgnd scs8hd_fill_2
XANTENNA__130__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _071_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_133 vpwr vgnd scs8hd_fill_2
XFILLER_9_211 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_9_ mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _064_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
X_162_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_10_232 vgnd vpwr scs8hd_fill_1
X_093_ _084_/B _092_/B _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_9 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__111__C _111_/C vgnd vpwr scs8hd_diode_2
Xmem_right_track_10.LATCH_0_.latch data_in _066_/A _132_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_217 vgnd vpwr scs8hd_decap_12
XFILLER_10_77 vgnd vpwr scs8hd_decap_6
XFILLER_19_42 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_63 vgnd vpwr scs8hd_decap_12
XFILLER_27_195 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vpwr vgnd scs8hd_fill_2
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XFILLER_19_97 vpwr vgnd scs8hd_fill_2
X_145_ _145_/HI _145_/LO vgnd vpwr scs8hd_conb_1
X_076_ _097_/A _084_/A _076_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_198 vpwr vgnd scs8hd_fill_2
XFILLER_33_176 vgnd vpwr scs8hd_decap_6
XFILLER_33_132 vgnd vpwr scs8hd_decap_8
XFILLER_33_110 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_121 vpwr vgnd scs8hd_fill_2
XFILLER_24_110 vpwr vgnd scs8hd_fill_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_4
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_65 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_7_12 vpwr vgnd scs8hd_fill_2
XFILLER_7_23 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A address[5] vgnd vpwr scs8hd_diode_2
X_128_ _130_/A address[6] _075_/C address[0] _128_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__117__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
X_059_ _059_/A _059_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _062_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_29_224 vgnd vpwr scs8hd_decap_8
XFILLER_16_21 vgnd vpwr scs8hd_decap_8
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XANTENNA__128__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_150 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _070_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_11 vpwr vgnd scs8hd_fill_2
XFILLER_14_219 vgnd vpwr scs8hd_decap_12
XFILLER_13_44 vgnd vpwr scs8hd_decap_3
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
XFILLER_13_99 vpwr vgnd scs8hd_fill_2
XFILLER_1_156 vpwr vgnd scs8hd_fill_2
XFILLER_1_101 vpwr vgnd scs8hd_fill_2
XFILLER_1_123 vgnd vpwr scs8hd_fill_1
Xmem_right_track_6.LATCH_0_.latch data_in _064_/A _130_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_223 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__051__A address[1] vgnd vpwr scs8hd_diode_2
X_161_ _161_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_24_54 vgnd vpwr scs8hd_decap_3
XFILLER_24_32 vpwr vgnd scs8hd_fill_2
XFILLER_24_10 vpwr vgnd scs8hd_fill_2
X_092_ _100_/A _092_/B _092_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__136__A _130_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _064_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_108 vgnd vpwr scs8hd_decap_4
XFILLER_3_229 vgnd vpwr scs8hd_decap_4
XFILLER_3_207 vgnd vpwr scs8hd_decap_8
XFILLER_10_89 vgnd vpwr scs8hd_fill_1
XFILLER_35_75 vgnd vpwr scs8hd_decap_4
XFILLER_27_130 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _151_/HI mem_top_track_8.LATCH_2_.latch/Q
+ mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_144_ _144_/HI _144_/LO vgnd vpwr scs8hd_conb_1
X_075_ address[5] address[6] _075_/C _084_/A vgnd vpwr scs8hd_or3_4
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _159_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_174 vgnd vpwr scs8hd_decap_4
XFILLER_33_188 vgnd vpwr scs8hd_decap_6
XFILLER_33_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_166 vpwr vgnd scs8hd_fill_2
XFILLER_24_133 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_1_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_44 vpwr vgnd scs8hd_fill_2
XFILLER_21_55 vpwr vgnd scs8hd_fill_2
XFILLER_30_169 vgnd vpwr scs8hd_decap_4
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_111 vgnd vpwr scs8hd_decap_4
XFILLER_15_144 vpwr vgnd scs8hd_fill_2
XFILLER_15_199 vgnd vpwr scs8hd_decap_6
X_058_ enable _095_/C vgnd vpwr scs8hd_inv_8
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_127_ _130_/A address[6] _075_/C _083_/C _127_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_16_3 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _169_/A vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vgnd vpwr scs8hd_decap_6
XFILLER_21_136 vgnd vpwr scs8hd_decap_3
XFILLER_8_107 vgnd vpwr scs8hd_decap_12
XFILLER_12_125 vgnd vpwr scs8hd_fill_1
XFILLER_12_158 vpwr vgnd scs8hd_fill_2
XFILLER_16_88 vgnd vpwr scs8hd_decap_4
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_8_129 vpwr vgnd scs8hd_fill_2
XANTENNA__128__B address[6] vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _060_/Y mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__054__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_98 vpwr vgnd scs8hd_fill_2
XFILLER_27_21 vgnd vpwr scs8hd_decap_4
XFILLER_4_154 vgnd vpwr scs8hd_decap_3
XFILLER_4_143 vgnd vpwr scs8hd_decap_8
XFILLER_4_110 vgnd vpwr scs8hd_decap_6
XFILLER_4_69 vgnd vpwr scs8hd_decap_4
XANTENNA__130__C _130_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vpwr vgnd scs8hd_fill_2
XFILLER_14_209 vgnd vpwr scs8hd_decap_4
XFILLER_13_34 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_113 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_220 vpwr vgnd scs8hd_fill_2
XANTENNA__125__C _111_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_88 vgnd vpwr scs8hd_decap_4
XFILLER_24_77 vpwr vgnd scs8hd_fill_2
XFILLER_24_66 vgnd vpwr scs8hd_decap_8
X_091_ _099_/A _092_/B _091_/Y vgnd vpwr scs8hd_nor2_4
X_160_ right_top_grid_pin_10_ chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_10_212 vpwr vgnd scs8hd_fill_2
XANTENNA__136__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__062__A _062_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_87 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
X_074_ address[4] address[3] _095_/C _075_/C vgnd vpwr scs8hd_or3_4
X_143_ _143_/HI _143_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_131 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_145 vpwr vgnd scs8hd_fill_2
XANTENNA__057__A address[3] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_23 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _066_/Y mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_3
XFILLER_30_137 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_057_ address[3] _057_/Y vgnd vpwr scs8hd_inv_8
X_126_ address[5] address[6] _111_/C address[0] _126_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__133__C _075_/C vgnd vpwr scs8hd_diode_2
XFILLER_30_6 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_10.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_119 vgnd vpwr scs8hd_fill_1
XFILLER_12_104 vgnd vpwr scs8hd_decap_6
XFILLER_12_115 vgnd vpwr scs8hd_decap_8
XFILLER_12_137 vpwr vgnd scs8hd_fill_2
XFILLER_16_67 vgnd vpwr scs8hd_decap_4
XFILLER_32_88 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_218 vgnd vpwr scs8hd_decap_12
XFILLER_35_207 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _072_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__128__C _075_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__160__A right_top_grid_pin_10_ vgnd vpwr scs8hd_diode_2
X_109_ _102_/A _106_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__070__A _070_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_88 vgnd vpwr scs8hd_decap_8
XFILLER_17_218 vpwr vgnd scs8hd_fill_2
XFILLER_17_229 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__130__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_fill_1
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__065__A _065_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_169 vpwr vgnd scs8hd_fill_2
XFILLER_9_203 vgnd vpwr scs8hd_fill_1
XFILLER_13_232 vgnd vpwr scs8hd_fill_1
XANTENNA__125__D _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_8
X_090_ _098_/A _092_/B _090_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_206 vgnd vpwr scs8hd_decap_4
XFILLER_10_224 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _068_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_49 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__136__C _096_/C vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_0_.latch data_in _060_/A _126_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_69 vpwr vgnd scs8hd_fill_2
XFILLER_27_176 vgnd vpwr scs8hd_decap_4
XFILLER_27_165 vgnd vpwr scs8hd_decap_4
XFILLER_27_143 vgnd vpwr scs8hd_decap_4
XFILLER_27_121 vgnd vpwr scs8hd_fill_1
XFILLER_19_23 vgnd vpwr scs8hd_decap_4
XFILLER_19_56 vpwr vgnd scs8hd_fill_2
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
X_142_ _142_/HI _142_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
X_073_ address[1] _077_/B _083_/C _097_/A vgnd vpwr scs8hd_or3_4
XFILLER_33_168 vgnd vpwr scs8hd_fill_1
XFILLER_18_154 vgnd vpwr scs8hd_fill_1
XANTENNA__163__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vpwr vgnd scs8hd_fill_2
XFILLER_24_179 vpwr vgnd scs8hd_fill_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_135 vgnd vpwr scs8hd_decap_6
XFILLER_30_105 vgnd vpwr scs8hd_decap_8
X_125_ address[5] address[6] _111_/C _083_/C _125_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_056_ address[4] _056_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__133__D _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA__158__A _158_/A vgnd vpwr scs8hd_diode_2
XANTENNA__068__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_13 vpwr vgnd scs8hd_fill_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_149 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _082_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__128__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_164 vpwr vgnd scs8hd_fill_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vgnd vpwr scs8hd_decap_6
X_108_ _084_/B _106_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_3 vgnd vpwr scs8hd_decap_3
XFILLER_26_219 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _063_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _174_/A vgnd vpwr scs8hd_inv_1
XFILLER_8_80 vgnd vpwr scs8hd_fill_1
XFILLER_27_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _143_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_189 vgnd vpwr scs8hd_decap_6
XFILLER_4_16 vgnd vpwr scs8hd_decap_8
XANTENNA__171__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_137 vpwr vgnd scs8hd_fill_2
XFILLER_8_7 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A _081_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_181 vgnd vpwr scs8hd_decap_4
XANTENNA__166__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__076__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_46 vgnd vpwr scs8hd_decap_8
XFILLER_1_28 vpwr vgnd scs8hd_fill_2
XANTENNA__136__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _105_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_46 vgnd vpwr scs8hd_decap_3
XFILLER_35_56 vgnd vpwr scs8hd_decap_6
XFILLER_27_199 vpwr vgnd scs8hd_fill_2
XFILLER_19_79 vpwr vgnd scs8hd_fill_2
X_141_ _141_/HI _141_/LO vgnd vpwr scs8hd_conb_1
X_072_ _072_/A _072_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XFILLER_18_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _069_/A vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _071_/A _137_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_125 vgnd vpwr scs8hd_decap_8
XFILLER_24_158 vgnd vpwr scs8hd_fill_1
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _077_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_69 vgnd vpwr scs8hd_decap_4
XFILLER_15_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_7_16 vpwr vgnd scs8hd_fill_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_3
X_055_ address[6] _134_/B vgnd vpwr scs8hd_inv_8
X_124_ _102_/A _121_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_36 vgnd vpwr scs8hd_decap_3
XFILLER_32_68 vgnd vpwr scs8hd_decap_6
XANTENNA__084__A _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_161 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_110 vpwr vgnd scs8hd_fill_2
X_107_ _100_/A _106_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_194 vpwr vgnd scs8hd_fill_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_3
XANTENNA__169__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _081_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_4_135 vpwr vgnd scs8hd_fill_2
XFILLER_4_179 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_3
XANTENNA__081__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_1_105 vpwr vgnd scs8hd_fill_2
XFILLER_13_201 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__076__B _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_36 vgnd vpwr scs8hd_fill_1
XFILLER_10_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _100_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
XFILLER_30_90 vpwr vgnd scs8hd_fill_2
XANTENNA__177__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_79 vgnd vpwr scs8hd_fill_1
XANTENNA__087__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_071_ _071_/A _071_/Y vgnd vpwr scs8hd_inv_8
X_140_ _140_/HI _140_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_101 vgnd vpwr scs8hd_decap_4
XFILLER_18_123 vpwr vgnd scs8hd_fill_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XFILLER_33_148 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_178 vgnd vpwr scs8hd_fill_1
XFILLER_2_83 vgnd vpwr scs8hd_decap_6
XANTENNA__073__C _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_115 vgnd vpwr scs8hd_fill_1
XFILLER_15_148 vpwr vgnd scs8hd_fill_2
X_054_ address[5] _130_/A vgnd vpwr scs8hd_inv_8
X_123_ _084_/B _121_/B _123_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _091_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_48 vgnd vpwr scs8hd_decap_8
XANTENNA__084__B _084_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_151 vpwr vgnd scs8hd_fill_2
XFILLER_11_151 vgnd vpwr scs8hd_fill_1
XFILLER_11_173 vpwr vgnd scs8hd_fill_2
XFILLER_7_133 vpwr vgnd scs8hd_fill_2
XFILLER_11_184 vgnd vpwr scs8hd_fill_1
X_106_ _099_/A _106_/B _106_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_93 vgnd vpwr scs8hd_decap_4
XFILLER_27_25 vgnd vpwr scs8hd_fill_1
XANTENNA__079__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _056_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_224 vgnd vpwr scs8hd_decap_8
XFILLER_31_213 vpwr vgnd scs8hd_fill_2
XFILLER_16_210 vpwr vgnd scs8hd_fill_2
XFILLER_16_232 vgnd vpwr scs8hd_fill_1
XFILLER_22_213 vgnd vpwr scs8hd_fill_1
XFILLER_13_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_49 vpwr vgnd scs8hd_fill_2
XANTENNA__081__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_224 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_94 vgnd vpwr scs8hd_fill_1
XANTENNA__092__B _092_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_231 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_113 vpwr vgnd scs8hd_fill_2
XFILLER_27_102 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vpwr vgnd scs8hd_fill_2
XANTENNA__087__B _057_/Y vgnd vpwr scs8hd_diode_2
X_070_ _070_/A _070_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _071_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_113 vgnd vpwr scs8hd_fill_1
XFILLER_18_135 vgnd vpwr scs8hd_fill_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _144_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_62 vpwr vgnd scs8hd_fill_2
XFILLER_24_149 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_160 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_27 vpwr vgnd scs8hd_fill_2
XANTENNA__098__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_182 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_053_ address[0] _083_/C vgnd vpwr scs8hd_inv_8
X_122_ _100_/A _121_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_208 vgnd vpwr scs8hd_decap_8
Xmem_right_track_10.LATCH_1_.latch data_in _065_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_130 vgnd vpwr scs8hd_decap_3
XFILLER_7_123 vgnd vpwr scs8hd_fill_1
XFILLER_7_156 vpwr vgnd scs8hd_fill_2
X_105_ _098_/A _106_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_81 vgnd vpwr scs8hd_decap_8
XFILLER_34_200 vgnd vpwr scs8hd_decap_3
XFILLER_19_230 vgnd vpwr scs8hd_decap_3
XFILLER_8_72 vgnd vpwr scs8hd_decap_8
XANTENNA__079__C _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_33_80 vgnd vpwr scs8hd_decap_6
XFILLER_3_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_9_207 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_0_195 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _070_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_18 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_147 vgnd vpwr scs8hd_fill_1
XANTENNA__087__C _095_/C vgnd vpwr scs8hd_diode_2
XFILLER_19_38 vpwr vgnd scs8hd_fill_2
XFILLER_35_180 vgnd vpwr scs8hd_decap_6
XFILLER_27_169 vgnd vpwr scs8hd_fill_1
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _139_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_183 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_106 vpwr vgnd scs8hd_fill_2
Xmem_right_track_6.LATCH_1_.latch data_in _063_/A _129_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_161 vpwr vgnd scs8hd_fill_2
X_121_ _099_/A _121_/B _121_/Y vgnd vpwr scs8hd_nor2_4
X_052_ address[2] _077_/B vgnd vpwr scs8hd_inv_8
XFILLER_16_17 vpwr vgnd scs8hd_fill_2
XFILLER_20_186 vgnd vpwr scs8hd_decap_3
XFILLER_28_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _064_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_168 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
X_104_ _097_/A _106_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_71 vgnd vpwr scs8hd_fill_1
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_8_84 vgnd vpwr scs8hd_decap_8
XFILLER_27_49 vgnd vpwr scs8hd_decap_6
XANTENNA__095__C _095_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_70 vpwr vgnd scs8hd_fill_2
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_9_219 vpwr vgnd scs8hd_fill_2
XFILLER_13_204 vgnd vpwr scs8hd_decap_4
XFILLER_0_185 vgnd vpwr scs8hd_fill_1
XFILLER_14_83 vpwr vgnd scs8hd_fill_2
XFILLER_30_93 vgnd vpwr scs8hd_fill_1
XFILLER_30_82 vgnd vpwr scs8hd_decap_8
XFILLER_35_27 vgnd vpwr scs8hd_decap_4
XFILLER_27_126 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _153_/A vgnd vpwr scs8hd_inv_1
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _170_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_75 vpwr vgnd scs8hd_fill_2
XFILLER_2_53 vgnd vpwr scs8hd_decap_6
XFILLER_2_42 vpwr vgnd scs8hd_fill_2
XFILLER_32_195 vpwr vgnd scs8hd_fill_2
XFILLER_32_151 vpwr vgnd scs8hd_fill_2
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vgnd vpwr scs8hd_decap_3
X_120_ _098_/A _121_/B _120_/Y vgnd vpwr scs8hd_nor2_4
X_051_ address[1] _081_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_51 vpwr vgnd scs8hd_fill_2
XFILLER_11_84 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_195 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_29 vpwr vgnd scs8hd_fill_2
XFILLER_20_143 vgnd vpwr scs8hd_decap_8
XFILLER_20_154 vgnd vpwr scs8hd_decap_4
XFILLER_20_165 vgnd vpwr scs8hd_fill_1
XFILLER_20_198 vpwr vgnd scs8hd_fill_2
X_103_ address[5] _134_/B _096_/C _106_/B vgnd vpwr scs8hd_or3_4
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_154 vpwr vgnd scs8hd_fill_2
XFILLER_11_198 vpwr vgnd scs8hd_fill_2
XFILLER_19_210 vgnd vpwr scs8hd_decap_4
XFILLER_27_28 vpwr vgnd scs8hd_fill_2
XFILLER_25_202 vpwr vgnd scs8hd_fill_2
XFILLER_4_139 vpwr vgnd scs8hd_fill_2
XFILLER_16_224 vgnd vpwr scs8hd_decap_8
XFILLER_22_227 vgnd vpwr scs8hd_decap_6
XFILLER_22_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XFILLER_5_97 vpwr vgnd scs8hd_fill_2
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vgnd vpwr scs8hd_fill_1
XFILLER_5_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _156_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_212 vpwr vgnd scs8hd_fill_2
XFILLER_14_62 vpwr vgnd scs8hd_fill_2
XFILLER_5_223 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__101__A _084_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_127 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_171 vgnd vpwr scs8hd_fill_1
XFILLER_25_83 vgnd vpwr scs8hd_fill_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_fill_1
XFILLER_21_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_174 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _139_/HI mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_14_141 vgnd vpwr scs8hd_decap_8
XFILLER_14_163 vpwr vgnd scs8hd_fill_2
XFILLER_14_174 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_18 vgnd vpwr scs8hd_decap_12
XFILLER_20_122 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_1_.latch data_in _059_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_111 vgnd vpwr scs8hd_fill_1
X_102_ _102_/A _102_/B _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_137 vpwr vgnd scs8hd_fill_2
XFILLER_11_177 vgnd vpwr scs8hd_decap_4
XFILLER_22_51 vgnd vpwr scs8hd_fill_1
XFILLER_19_222 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_97 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_51 vpwr vgnd scs8hd_fill_2
XFILLER_3_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_173 vpwr vgnd scs8hd_fill_2
XANTENNA__104__A _097_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_50 vgnd vpwr scs8hd_decap_8
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _080_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_232 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_41 vpwr vgnd scs8hd_fill_2
XFILLER_29_191 vpwr vgnd scs8hd_fill_2
XANTENNA__101__B _102_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_117 vpwr vgnd scs8hd_fill_2
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_183 vgnd vpwr scs8hd_decap_4
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_95 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XANTENNA__112__A _097_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_161 vgnd vpwr scs8hd_decap_3
XFILLER_32_164 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_153 vgnd vpwr scs8hd_decap_6
XANTENNA__107__A _100_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_112 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_178 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_101_ _084_/B _102_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_123 vgnd vpwr scs8hd_decap_3
XFILLER_22_63 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _069_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_62 vgnd vpwr scs8hd_decap_8
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_152 vgnd vpwr scs8hd_decap_4
XANTENNA__104__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _098_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_84 vgnd vpwr scs8hd_decap_8
XFILLER_28_62 vgnd vpwr scs8hd_decap_12
XFILLER_28_40 vgnd vpwr scs8hd_fill_1
XFILLER_0_199 vgnd vpwr scs8hd_fill_1
XFILLER_0_177 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _100_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_88 vgnd vpwr scs8hd_decap_6
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_14_75 vpwr vgnd scs8hd_fill_2
XFILLER_29_170 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_107 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_63 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_2_89 vgnd vpwr scs8hd_fill_1
XANTENNA__112__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_6
XFILLER_32_110 vgnd vpwr scs8hd_decap_3
XFILLER_17_184 vpwr vgnd scs8hd_fill_2
XFILLER_23_198 vpwr vgnd scs8hd_fill_2
XFILLER_23_132 vgnd vpwr scs8hd_decap_4
XFILLER_11_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_11_65 vpwr vgnd scs8hd_fill_2
X_177_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__107__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _084_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_135 vpwr vgnd scs8hd_fill_2
XFILLER_20_168 vgnd vpwr scs8hd_fill_1
XFILLER_28_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
X_100_ _100_/A _102_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_106 vpwr vgnd scs8hd_fill_2
XFILLER_22_97 vpwr vgnd scs8hd_fill_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_6
XFILLER_8_11 vpwr vgnd scs8hd_fill_2
XANTENNA__118__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_194 vgnd vpwr scs8hd_fill_1
XFILLER_8_55 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_30 vpwr vgnd scs8hd_fill_2
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XFILLER_3_120 vpwr vgnd scs8hd_fill_2
XFILLER_3_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_208 vgnd vpwr scs8hd_fill_1
XFILLER_21_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_74 vgnd vpwr scs8hd_decap_4
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _090_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_56 vpwr vgnd scs8hd_fill_2
XFILLER_5_45 vpwr vgnd scs8hd_fill_2
XFILLER_5_12 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _130_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_21 vpwr vgnd scs8hd_fill_2
XFILLER_14_87 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_182 vgnd vpwr scs8hd_fill_1
XANTENNA__126__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_163 vgnd vpwr scs8hd_decap_8
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_79 vpwr vgnd scs8hd_fill_2
XFILLER_2_46 vgnd vpwr scs8hd_decap_4
XFILLER_32_122 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_111 vgnd vpwr scs8hd_fill_1
XFILLER_11_33 vpwr vgnd scs8hd_fill_2
XFILLER_11_55 vgnd vpwr scs8hd_decap_4
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_176_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__123__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_103 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_214 vgnd vpwr scs8hd_fill_1
XFILLER_8_45 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__134__A address[5] vgnd vpwr scs8hd_diode_2
X_159_ _159_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_8
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
XFILLER_17_43 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_fill_1
XFILLER_31_209 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _130_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_146 vgnd vpwr scs8hd_decap_3
XFILLER_28_97 vgnd vpwr scs8hd_decap_3
XFILLER_8_202 vgnd vpwr scs8hd_fill_1
XFILLER_8_224 vgnd vpwr scs8hd_decap_8
XFILLER_5_24 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_216 vpwr vgnd scs8hd_fill_2
XFILLER_5_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__126__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__052__A address[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_3_ mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_43 vgnd vpwr scs8hd_decap_4
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_175 vgnd vpwr scs8hd_decap_4
XFILLER_17_197 vgnd vpwr scs8hd_decap_4
XFILLER_23_189 vgnd vpwr scs8hd_decap_6
XFILLER_23_178 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_101 vgnd vpwr scs8hd_fill_1
XFILLER_14_167 vgnd vpwr scs8hd_decap_4
X_175_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_9_160 vpwr vgnd scs8hd_fill_2
XFILLER_20_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ _064_/A mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_226 vpwr vgnd scs8hd_fill_2
XFILLER_8_24 vgnd vpwr scs8hd_fill_1
XFILLER_8_68 vpwr vgnd scs8hd_fill_2
XANTENNA__118__C _075_/C vgnd vpwr scs8hd_diode_2
X_089_ _097_/A _092_/B _089_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_163 vgnd vpwr scs8hd_decap_3
X_158_ _158_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__134__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA__060__A _060_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_22 vpwr vgnd scs8hd_fill_2
XFILLER_17_55 vgnd vpwr scs8hd_decap_4
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XFILLER_33_76 vpwr vgnd scs8hd_fill_2
XFILLER_3_177 vpwr vgnd scs8hd_fill_2
XFILLER_3_188 vgnd vpwr scs8hd_decap_4
XANTENNA__129__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__055__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_103 vgnd vpwr scs8hd_decap_6
XFILLER_28_32 vgnd vpwr scs8hd_decap_8
XFILLER_0_169 vgnd vpwr scs8hd_decap_4
XFILLER_12_232 vgnd vpwr scs8hd_fill_1
XANTENNA__131__C _111_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_45 vpwr vgnd scs8hd_fill_2
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_195 vpwr vgnd scs8hd_fill_2
XFILLER_29_184 vpwr vgnd scs8hd_fill_2
XFILLER_29_162 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__126__C _111_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_187 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _149_/HI mem_top_track_0.LATCH_2_.latch/Q
+ mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_132 vpwr vgnd scs8hd_fill_2
XFILLER_25_99 vgnd vpwr scs8hd_decap_4
XFILLER_25_11 vpwr vgnd scs8hd_fill_2
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_2_59 vgnd vpwr scs8hd_fill_1
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_102 vgnd vpwr scs8hd_decap_8
XFILLER_17_132 vgnd vpwr scs8hd_decap_4
XFILLER_32_168 vgnd vpwr scs8hd_decap_6
XANTENNA__137__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _153_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__063__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_13 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_174_ _174_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_91 vpwr vgnd scs8hd_fill_2
XANTENNA__058__A enable vgnd vpwr scs8hd_diode_2
XFILLER_22_67 vgnd vpwr scs8hd_decap_4
XFILLER_22_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _157_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__134__C _075_/C vgnd vpwr scs8hd_diode_2
XFILLER_10_171 vgnd vpwr scs8hd_decap_12
XFILLER_10_193 vpwr vgnd scs8hd_fill_2
X_088_ address[5] address[6] _130_/C _092_/B vgnd vpwr scs8hd_or3_4
XFILLER_25_219 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_156 vgnd vpwr scs8hd_fill_1
XFILLER_3_112 vpwr vgnd scs8hd_fill_2
XFILLER_30_200 vpwr vgnd scs8hd_fill_2
XANTENNA__129__C _130_/C vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_211 vgnd vpwr scs8hd_decap_4
XFILLER_21_222 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_115 vpwr vgnd scs8hd_fill_2
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_11 vgnd vpwr scs8hd_fill_1
XANTENNA__131__D _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _155_/A vgnd vpwr scs8hd_inv_1
XANTENNA__156__A _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA__066__A _066_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_35 vgnd vpwr scs8hd_decap_4
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_79 vpwr vgnd scs8hd_fill_2
XFILLER_29_174 vpwr vgnd scs8hd_fill_2
XFILLER_29_130 vpwr vgnd scs8hd_fill_2
XANTENNA__126__D address[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_199 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_232 vgnd vpwr scs8hd_fill_1
XFILLER_17_100 vpwr vgnd scs8hd_fill_2
XFILLER_17_188 vgnd vpwr scs8hd_decap_6
XANTENNA__137__C _130_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _060_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_25 vgnd vpwr scs8hd_fill_1
XFILLER_11_47 vpwr vgnd scs8hd_fill_2
XFILLER_11_69 vgnd vpwr scs8hd_decap_4
XFILLER_14_125 vgnd vpwr scs8hd_fill_1
X_173_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_20_139 vpwr vgnd scs8hd_fill_2
XANTENNA__164__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_9_184 vpwr vgnd scs8hd_fill_2
XFILLER_9_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_70 vpwr vgnd scs8hd_fill_2
XFILLER_28_206 vgnd vpwr scs8hd_decap_8
XANTENNA__074__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_11_128 vpwr vgnd scs8hd_fill_2
XFILLER_11_139 vgnd vpwr scs8hd_decap_12
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_217 vgnd vpwr scs8hd_fill_1
X_087_ address[4] _057_/Y _095_/C _130_/C vgnd vpwr scs8hd_or3_4
X_156_ _156_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_6_154 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_11_ mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__134__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_10_183 vgnd vpwr scs8hd_fill_1
XANTENNA__159__A _159_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_231 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_79 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_212 vpwr vgnd scs8hd_fill_2
XANTENNA__129__D _083_/C vgnd vpwr scs8hd_diode_2
X_139_ _139_/HI _139_/LO vgnd vpwr scs8hd_conb_1
XFILLER_31_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _158_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_78 vgnd vpwr scs8hd_fill_1
XFILLER_5_49 vgnd vpwr scs8hd_decap_4
XFILLER_5_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_25 vpwr vgnd scs8hd_fill_2
XFILLER_14_58 vpwr vgnd scs8hd_fill_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A _084_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_26_189 vpwr vgnd scs8hd_fill_2
XFILLER_26_145 vgnd vpwr scs8hd_decap_8
XFILLER_25_24 vpwr vgnd scs8hd_fill_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_79 vgnd vpwr scs8hd_decap_4
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_222 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_126 vgnd vpwr scs8hd_decap_4
XANTENNA__137__D _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_192 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _078_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_37 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _069_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_172_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _145_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_152 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__074__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_11_107 vgnd vpwr scs8hd_decap_4
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XFILLER_22_47 vgnd vpwr scs8hd_decap_4
XANTENNA__090__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
XFILLER_8_49 vgnd vpwr scs8hd_decap_4
X_155_ _155_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_122 vpwr vgnd scs8hd_fill_2
XFILLER_6_188 vgnd vpwr scs8hd_decap_6
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
X_086_ _084_/A _102_/A _086_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__175__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_14 vpwr vgnd scs8hd_fill_2
XFILLER_33_35 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_3_169 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_232 vgnd vpwr scs8hd_fill_1
X_138_ address[5] _134_/B _130_/C address[0] _138_/Y vgnd vpwr scs8hd_nor4_4
X_069_ _069_/A _069_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ _062_/A mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_9_92 vgnd vpwr scs8hd_decap_3
XFILLER_8_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XFILLER_12_224 vgnd vpwr scs8hd_decap_8
Xmem_right_track_12.LATCH_0_.latch data_in _068_/A _134_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__082__B _100_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_6_71 vgnd vpwr scs8hd_decap_4
XFILLER_6_93 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _178_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_124 vgnd vpwr scs8hd_decap_8
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _077_/B vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _084_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_157 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_138 vpwr vgnd scs8hd_fill_2
XFILLER_23_149 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_149 vpwr vgnd scs8hd_fill_2
X_171_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_22_182 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_164 vgnd vpwr scs8hd_decap_8
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_20_108 vgnd vpwr scs8hd_decap_4
XFILLER_28_219 vgnd vpwr scs8hd_decap_12
XANTENNA__074__C _095_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__090__B _092_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ _068_/A mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_154_ _154_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_145 vgnd vpwr scs8hd_decap_8
X_085_ address[1] address[2] address[0] _102_/A vgnd vpwr scs8hd_or3_4
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_26 vpwr vgnd scs8hd_fill_2
XFILLER_33_14 vpwr vgnd scs8hd_fill_2
XANTENNA__085__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_159 vgnd vpwr scs8hd_fill_1
XFILLER_3_126 vgnd vpwr scs8hd_decap_3
Xmem_right_track_8.LATCH_0_.latch data_in _070_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_137_ address[5] _134_/B _130_/C _083_/C _137_/Y vgnd vpwr scs8hd_nor4_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_068_ _068_/A _068_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_14 vgnd vpwr scs8hd_decap_12
XFILLER_28_58 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _066_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_80 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_29_166 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_232 vgnd vpwr scs8hd_fill_1
XFILLER_35_125 vgnd vpwr scs8hd_decap_12
XFILLER_29_90 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA__077__C address[0] vgnd vpwr scs8hd_diode_2
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__B _092_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_32_139 vgnd vpwr scs8hd_decap_12
XFILLER_31_91 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _089_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__088__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_22_194 vpwr vgnd scs8hd_fill_2
XFILLER_22_172 vgnd vpwr scs8hd_fill_1
XFILLER_22_150 vgnd vpwr scs8hd_decap_3
X_170_ _170_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_14_128 vpwr vgnd scs8hd_fill_2
XFILLER_9_110 vpwr vgnd scs8hd_fill_2
XFILLER_3_95 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_18 vgnd vpwr scs8hd_decap_6
X_153_ _153_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
X_084_ _084_/A _084_/B _084_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_197 vgnd vpwr scs8hd_decap_4
XFILLER_12_82 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_223 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_24_201 vgnd vpwr scs8hd_decap_4
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__085__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_116 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_92 vpwr vgnd scs8hd_fill_2
X_136_ _130_/A address[6] _096_/C address[0] _136_/Y vgnd vpwr scs8hd_nor4_4
X_067_ _067_/A _067_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_63 vpwr vgnd scs8hd_fill_2
XFILLER_0_74 vgnd vpwr scs8hd_decap_6
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_28_26 vgnd vpwr scs8hd_decap_4
XFILLER_0_119 vgnd vpwr scs8hd_decap_3
XANTENNA__096__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _149_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _059_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
X_119_ _097_/A _121_/B _119_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_2.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_178 vpwr vgnd scs8hd_fill_2
XFILLER_29_134 vgnd vpwr scs8hd_decap_3
XFILLER_20_71 vgnd vpwr scs8hd_fill_1
XFILLER_35_137 vgnd vpwr scs8hd_decap_12
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XFILLER_25_49 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_1_214 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_104 vgnd vpwr scs8hd_decap_4
XFILLER_15_93 vgnd vpwr scs8hd_decap_3
XFILLER_31_151 vpwr vgnd scs8hd_fill_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_107 vgnd vpwr scs8hd_decap_4
XFILLER_16_181 vgnd vpwr scs8hd_decap_3
XFILLER_31_184 vgnd vpwr scs8hd_decap_3
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
XANTENNA__088__C _130_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_199 vpwr vgnd scs8hd_fill_2
XFILLER_13_173 vgnd vpwr scs8hd_decap_4
XFILLER_3_52 vpwr vgnd scs8hd_fill_2
XFILLER_3_41 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__099__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_232 vgnd vpwr scs8hd_fill_1
X_152_ _152_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_12_61 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_083_ address[1] address[2] _083_/C _084_/B vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_6_169 vgnd vpwr scs8hd_decap_6
XFILLER_33_202 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _063_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_210 vgnd vpwr scs8hd_decap_4
XFILLER_18_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_39 vpwr vgnd scs8hd_fill_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_6
XFILLER_15_224 vgnd vpwr scs8hd_decap_8
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
X_135_ _130_/A address[6] _096_/C _083_/C _135_/Y vgnd vpwr scs8hd_nor4_4
X_066_ _066_/A _066_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_7 vgnd vpwr scs8hd_decap_12
XFILLER_24_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_194 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__096__C _096_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
X_118_ _130_/A _134_/B _075_/C _121_/B vgnd vpwr scs8hd_or3_4
Xmem_right_track_4.LATCH_0_.latch data_in _062_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_3
XFILLER_14_29 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _060_/A mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_70 vgnd vpwr scs8hd_fill_1
XFILLER_35_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_30 vgnd vpwr scs8hd_fill_1
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_25_28 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_1_226 vgnd vpwr scs8hd_decap_6
XFILLER_25_160 vpwr vgnd scs8hd_fill_2
XFILLER_17_138 vpwr vgnd scs8hd_fill_2
XFILLER_17_149 vgnd vpwr scs8hd_decap_6
XFILLER_15_72 vpwr vgnd scs8hd_fill_2
XFILLER_31_163 vgnd vpwr scs8hd_decap_3
XFILLER_31_130 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _071_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_108 vpwr vgnd scs8hd_fill_2
XFILLER_14_119 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _147_/HI _064_/Y mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_3
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _146_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_222 vpwr vgnd scs8hd_fill_2
X_151_ _151_/HI _151_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_126 vgnd vpwr scs8hd_decap_12
XFILLER_6_159 vpwr vgnd scs8hd_fill_2
XFILLER_10_133 vpwr vgnd scs8hd_fill_2
XFILLER_12_40 vpwr vgnd scs8hd_fill_2
X_082_ _084_/A _100_/A _082_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _150_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_214 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_50 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_065_ _065_/A _065_/Y vgnd vpwr scs8hd_inv_8
X_134_ address[5] _134_/B _075_/C address[0] _134_/Y vgnd vpwr scs8hd_nor4_4
Xmux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ _066_/A mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
X_117_ _102_/A _116_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_18 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _070_/A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_103 vpwr vgnd scs8hd_fill_2
XFILLER_29_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_224 vgnd vpwr scs8hd_decap_8
XFILLER_4_213 vgnd vpwr scs8hd_fill_1
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
XFILLER_34_150 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_15_51 vgnd vpwr scs8hd_fill_1
XFILLER_15_62 vgnd vpwr scs8hd_decap_3
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_142 vpwr vgnd scs8hd_fill_2
XFILLER_26_72 vgnd vpwr scs8hd_fill_1
XFILLER_13_197 vgnd vpwr scs8hd_decap_4
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_190 vpwr vgnd scs8hd_fill_2
XFILLER_22_19 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _065_/A vgnd
+ vpwr scs8hd_diode_2
X_150_ _150_/HI _150_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_138 vgnd vpwr scs8hd_decap_4
XFILLER_12_74 vgnd vpwr scs8hd_decap_8
X_081_ _081_/A address[2] address[0] _100_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_18 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XFILLER_3_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _060_/Y vgnd vpwr
+ scs8hd_diode_2
X_133_ address[5] _134_/B _075_/C _083_/C _133_/Y vgnd vpwr scs8hd_nor4_4
X_064_ _064_/A _064_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_163 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A _056_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_207 vpwr vgnd scs8hd_fill_2
XFILLER_21_218 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XFILLER_9_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_83 vgnd vpwr scs8hd_decap_8
X_116_ _084_/B _116_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_126 vpwr vgnd scs8hd_fill_2
XFILLER_20_41 vgnd vpwr scs8hd_decap_8
XFILLER_20_63 vpwr vgnd scs8hd_fill_2
XFILLER_20_74 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vgnd vpwr scs8hd_decap_6
XFILLER_29_50 vgnd vpwr scs8hd_decap_8
XFILLER_28_192 vgnd vpwr scs8hd_fill_1
XFILLER_26_107 vgnd vpwr scs8hd_decap_8
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _094_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_25_184 vgnd vpwr scs8hd_decap_3
XFILLER_25_151 vgnd vpwr scs8hd_decap_3
XFILLER_15_30 vpwr vgnd scs8hd_fill_2
XFILLER_31_95 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XANTENNA__102__B _102_/B vgnd vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_143 vgnd vpwr scs8hd_decap_8
XFILLER_22_165 vgnd vpwr scs8hd_decap_4
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _062_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vgnd vpwr scs8hd_decap_12
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XFILLER_13_143 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_080_ _084_/A _099_/A _080_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_15_ mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_64 vgnd vpwr scs8hd_fill_1
XFILLER_18_224 vgnd vpwr scs8hd_decap_8
XANTENNA__108__A _084_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_6
XFILLER_24_205 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_216 vpwr vgnd scs8hd_fill_2
X_063_ _063_/A _063_/Y vgnd vpwr scs8hd_inv_8
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _076_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_30 vgnd vpwr scs8hd_fill_1
X_132_ _130_/A address[6] _111_/C address[0] _132_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_186 vgnd vpwr scs8hd_decap_8
XFILLER_2_175 vgnd vpwr scs8hd_decap_8
XFILLER_2_131 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__110__B _057_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_23 vgnd vpwr scs8hd_decap_8
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_9_21 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _061_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _060_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_41 vgnd vpwr scs8hd_decap_8
XFILLER_18_85 vpwr vgnd scs8hd_fill_2
XFILLER_11_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
X_115_ _100_/A _116_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_223 vpwr vgnd scs8hd_fill_2
XANTENNA__105__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__121__A _099_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_8
XFILLER_29_73 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _084_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_55 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vpwr scs8hd_fill_1
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_218 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _148_/HI _069_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_108 vgnd vpwr scs8hd_fill_1
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _141_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

