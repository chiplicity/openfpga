magic
tech EFS8A
magscale 1 2
timestamp 1602873619
<< locali >>
rect 11655 24225 11690 24259
rect 8493 23171 8527 23205
rect 7331 23137 7366 23171
rect 8493 23137 8654 23171
rect 11287 23137 11322 23171
rect 15427 23137 15554 23171
rect 6227 22049 6262 22083
rect 11563 22049 11598 22083
rect 6831 21097 6837 21131
rect 6831 21029 6865 21097
rect 13271 20009 13277 20043
rect 13271 19941 13305 20009
rect 1443 19873 1478 19907
rect 8119 19159 8153 19227
rect 12903 19159 12937 19227
rect 15295 19159 15329 19227
rect 8119 19125 8125 19159
rect 12903 19125 12909 19159
rect 15295 19125 15301 19159
rect 13179 18921 13185 18955
rect 8493 18819 8527 18921
rect 13179 18853 13213 18921
rect 1903 18785 2030 18819
rect 8493 18785 8654 18819
rect 11747 18785 11782 18819
rect 8493 18751 8527 18785
rect 12081 18207 12115 18377
rect 6371 17833 6377 17867
rect 6371 17765 6405 17833
rect 16899 17765 16944 17799
rect 7849 17051 7883 17221
rect 3755 17017 3893 17051
rect 21051 16745 21097 16779
rect 22971 16609 23006 16643
rect 15669 16031 15703 16201
rect 16129 15963 16163 16201
rect 4531 15895 4565 15963
rect 4531 15861 4537 15895
rect 13363 15657 13369 15691
rect 13363 15589 13397 15657
rect 8619 15521 8654 15555
rect 6469 14875 6503 15113
rect 19435 14569 19441 14603
rect 19435 14501 19469 14569
rect 14841 13923 14875 14025
rect 4439 13481 4445 13515
rect 6647 13481 6653 13515
rect 12995 13481 13001 13515
rect 4439 13413 4473 13481
rect 6647 13413 6681 13481
rect 12995 13413 13029 13481
rect 5457 12835 5491 12937
rect 13277 12631 13311 12937
rect 15209 12631 15243 12937
rect 21275 12393 21281 12427
rect 21275 12325 21309 12393
rect 10609 11747 10643 11849
rect 7935 11305 7941 11339
rect 13731 11305 13737 11339
rect 7935 11237 7969 11305
rect 13731 11237 13765 11305
rect 25375 10761 25513 10795
rect 3433 10523 3467 10761
rect 22287 10217 22293 10251
rect 22287 10149 22321 10217
rect 949 9707 983 10149
rect 12023 10081 12058 10115
rect 20855 10081 20982 10115
rect 17233 9503 17267 9673
rect 7935 9129 7941 9163
rect 12443 9129 12449 9163
rect 7935 9061 7969 9129
rect 12443 9061 12477 9129
rect 13553 8823 13587 9129
rect 20085 8415 20119 8517
rect 7935 8279 7969 8347
rect 15847 8279 15881 8347
rect 7935 8245 7941 8279
rect 15847 8245 15853 8279
rect 11799 8041 11805 8075
rect 11799 7973 11833 8041
rect 5359 7191 5393 7259
rect 5359 7157 5365 7191
rect 12587 7157 12725 7191
rect 18239 6953 18245 6987
rect 6043 6885 6088 6919
rect 18239 6885 18273 6953
rect 15243 6817 15370 6851
rect 22937 6647 22971 6953
rect 17233 6239 17267 6409
rect 22937 6307 22971 6409
rect 3249 5559 3283 5865
rect 4715 5865 4721 5899
rect 7383 5865 7389 5899
rect 15663 5865 15669 5899
rect 4715 5797 4749 5865
rect 7383 5797 7417 5865
rect 15663 5797 15697 5865
rect 7199 5015 7233 5083
rect 7199 4981 7205 5015
rect 3617 3451 3651 3689
rect 9229 3587 9263 3689
rect 10517 3587 10551 3689
rect 22707 3145 22845 3179
rect 7291 2839 7325 2907
rect 7291 2805 7297 2839
rect 8493 2295 8527 2601
rect 10885 2295 10919 2601
rect 24869 2499 24903 2601
<< viali >>
rect 18245 24361 18279 24395
rect 10676 24225 10710 24259
rect 11621 24225 11655 24259
rect 16957 24225 16991 24259
rect 18061 24225 18095 24259
rect 17141 24089 17175 24123
rect 10747 24021 10781 24055
rect 11759 24021 11793 24055
rect 1593 23817 1627 23851
rect 10701 23817 10735 23851
rect 14565 23817 14599 23851
rect 16221 23817 16255 23851
rect 18613 23817 18647 23851
rect 20361 23817 20395 23851
rect 22569 23817 22603 23851
rect 24777 23817 24811 23851
rect 21465 23749 21499 23783
rect 1409 23613 1443 23647
rect 1961 23613 1995 23647
rect 8953 23613 8987 23647
rect 9413 23613 9447 23647
rect 11136 23613 11170 23647
rect 12484 23613 12518 23647
rect 12909 23613 12943 23647
rect 14381 23613 14415 23647
rect 14933 23613 14967 23647
rect 16037 23613 16071 23647
rect 16589 23613 16623 23647
rect 17877 23613 17911 23647
rect 18061 23613 18095 23647
rect 20177 23613 20211 23647
rect 21281 23613 21315 23647
rect 21833 23613 21867 23647
rect 22385 23613 22419 23647
rect 22937 23613 22971 23647
rect 24593 23613 24627 23647
rect 25145 23613 25179 23647
rect 16957 23545 16991 23579
rect 9137 23477 9171 23511
rect 9965 23477 9999 23511
rect 11207 23477 11241 23511
rect 11713 23477 11747 23511
rect 12587 23477 12621 23511
rect 18245 23477 18279 23511
rect 20821 23477 20855 23511
rect 1593 23273 1627 23307
rect 11161 23273 11195 23307
rect 13691 23273 13725 23307
rect 18245 23273 18279 23307
rect 24777 23273 24811 23307
rect 8493 23205 8527 23239
rect 9873 23205 9907 23239
rect 1409 23137 1443 23171
rect 7297 23137 7331 23171
rect 11253 23137 11287 23171
rect 12300 23137 12334 23171
rect 13620 23137 13654 23171
rect 15393 23137 15427 23171
rect 16808 23137 16842 23171
rect 18061 23137 18095 23171
rect 24593 23137 24627 23171
rect 9781 23069 9815 23103
rect 10057 23069 10091 23103
rect 7435 22933 7469 22967
rect 7757 22933 7791 22967
rect 8723 22933 8757 22967
rect 11391 22933 11425 22967
rect 12403 22933 12437 22967
rect 15623 22933 15657 22967
rect 16911 22933 16945 22967
rect 1593 22729 1627 22763
rect 7205 22729 7239 22763
rect 8585 22729 8619 22763
rect 10241 22729 10275 22763
rect 14933 22729 14967 22763
rect 16773 22729 16807 22763
rect 10609 22661 10643 22695
rect 11345 22661 11379 22695
rect 17095 22661 17129 22695
rect 18245 22661 18279 22695
rect 7389 22593 7423 22627
rect 7665 22593 7699 22627
rect 9597 22593 9631 22627
rect 14289 22593 14323 22627
rect 1409 22525 1443 22559
rect 1961 22525 1995 22559
rect 5768 22525 5802 22559
rect 10860 22525 10894 22559
rect 11621 22525 11655 22559
rect 12449 22525 12483 22559
rect 13277 22525 13311 22559
rect 13528 22525 13562 22559
rect 14013 22525 14047 22559
rect 14508 22525 14542 22559
rect 17024 22525 17058 22559
rect 17417 22525 17451 22559
rect 5871 22457 5905 22491
rect 6653 22457 6687 22491
rect 7481 22457 7515 22491
rect 9321 22457 9355 22491
rect 9413 22457 9447 22491
rect 12909 22457 12943 22491
rect 14611 22457 14645 22491
rect 15577 22457 15611 22491
rect 6285 22389 6319 22423
rect 9045 22389 9079 22423
rect 10931 22389 10965 22423
rect 12633 22389 12667 22423
rect 13599 22389 13633 22423
rect 15669 22389 15703 22423
rect 24593 22389 24627 22423
rect 1685 22185 1719 22219
rect 6331 22185 6365 22219
rect 8861 22185 8895 22219
rect 11069 22185 11103 22219
rect 12449 22185 12483 22219
rect 7389 22117 7423 22151
rect 10149 22117 10183 22151
rect 13185 22117 13219 22151
rect 13277 22117 13311 22151
rect 16129 22117 16163 22151
rect 6193 22049 6227 22083
rect 11529 22049 11563 22083
rect 5181 21981 5215 22015
rect 7297 21981 7331 22015
rect 7573 21981 7607 22015
rect 10057 21981 10091 22015
rect 16037 21981 16071 22015
rect 10609 21913 10643 21947
rect 13737 21913 13771 21947
rect 14289 21913 14323 21947
rect 16589 21913 16623 21947
rect 9321 21845 9355 21879
rect 11667 21845 11701 21879
rect 12817 21845 12851 21879
rect 1593 21641 1627 21675
rect 11529 21641 11563 21675
rect 13737 21641 13771 21675
rect 24777 21641 24811 21675
rect 10977 21573 11011 21607
rect 12265 21573 12299 21607
rect 14933 21573 14967 21607
rect 5641 21505 5675 21539
rect 7573 21505 7607 21539
rect 8217 21505 8251 21539
rect 8861 21505 8895 21539
rect 9137 21505 9171 21539
rect 10425 21505 10459 21539
rect 12817 21505 12851 21539
rect 13461 21505 13495 21539
rect 14381 21505 14415 21539
rect 15669 21505 15703 21539
rect 15945 21505 15979 21539
rect 17233 21505 17267 21539
rect 1409 21437 1443 21471
rect 1961 21437 1995 21471
rect 4572 21437 4606 21471
rect 4675 21437 4709 21471
rect 5784 21437 5818 21471
rect 6285 21437 6319 21471
rect 18128 21437 18162 21471
rect 18521 21437 18555 21471
rect 24593 21437 24627 21471
rect 25145 21437 25179 21471
rect 5871 21369 5905 21403
rect 7297 21369 7331 21403
rect 7389 21369 7423 21403
rect 8953 21369 8987 21403
rect 10517 21369 10551 21403
rect 12909 21369 12943 21403
rect 14473 21369 14507 21403
rect 16037 21369 16071 21403
rect 16589 21369 16623 21403
rect 5089 21301 5123 21335
rect 6653 21301 6687 21335
rect 7113 21301 7147 21335
rect 8585 21301 8619 21335
rect 9873 21301 9907 21335
rect 10149 21301 10183 21335
rect 14197 21301 14231 21335
rect 15301 21301 15335 21335
rect 16957 21301 16991 21335
rect 18199 21301 18233 21335
rect 5273 21097 5307 21131
rect 6837 21097 6871 21131
rect 7389 21097 7423 21131
rect 8033 21097 8067 21131
rect 8723 21097 8757 21131
rect 9505 21097 9539 21131
rect 10609 21029 10643 21063
rect 13737 21029 13771 21063
rect 13829 21029 13863 21063
rect 14381 21029 14415 21063
rect 15945 21029 15979 21063
rect 16037 21029 16071 21063
rect 17509 21029 17543 21063
rect 17601 21029 17635 21063
rect 4445 20961 4479 20995
rect 5524 20961 5558 20995
rect 8652 20961 8686 20995
rect 12081 20961 12115 20995
rect 12541 20961 12575 20995
rect 6469 20893 6503 20927
rect 10517 20893 10551 20927
rect 12817 20893 12851 20927
rect 13277 20893 13311 20927
rect 16405 20893 16439 20927
rect 17785 20893 17819 20927
rect 11069 20825 11103 20859
rect 15761 20825 15795 20859
rect 4629 20757 4663 20791
rect 5595 20757 5629 20791
rect 6285 20757 6319 20791
rect 7665 20757 7699 20791
rect 9045 20757 9079 20791
rect 10149 20757 10183 20791
rect 16865 20757 16899 20791
rect 3341 20553 3375 20587
rect 7757 20553 7791 20587
rect 8493 20553 8527 20587
rect 9689 20553 9723 20587
rect 9965 20553 9999 20587
rect 11161 20553 11195 20587
rect 12081 20553 12115 20587
rect 12633 20553 12667 20587
rect 14197 20553 14231 20587
rect 15853 20553 15887 20587
rect 17417 20553 17451 20587
rect 17785 20553 17819 20587
rect 4629 20485 4663 20519
rect 18199 20485 18233 20519
rect 8677 20417 8711 20451
rect 9137 20417 9171 20451
rect 10241 20417 10275 20451
rect 10609 20417 10643 20451
rect 13277 20417 13311 20451
rect 16221 20417 16255 20451
rect 16865 20417 16899 20451
rect 18613 20417 18647 20451
rect 1752 20349 1786 20383
rect 2856 20349 2890 20383
rect 3836 20349 3870 20383
rect 4261 20349 4295 20383
rect 5089 20349 5123 20383
rect 5181 20349 5215 20383
rect 5641 20349 5675 20383
rect 6837 20349 6871 20383
rect 15092 20349 15126 20383
rect 18128 20349 18162 20383
rect 19124 20349 19158 20383
rect 19533 20349 19567 20383
rect 5917 20281 5951 20315
rect 7199 20281 7233 20315
rect 8769 20281 8803 20315
rect 10333 20281 10367 20315
rect 13598 20281 13632 20315
rect 16313 20281 16347 20315
rect 19211 20281 19245 20315
rect 1823 20213 1857 20247
rect 2237 20213 2271 20247
rect 2927 20213 2961 20247
rect 3939 20213 3973 20247
rect 6193 20213 6227 20247
rect 6561 20213 6595 20247
rect 8033 20213 8067 20247
rect 13185 20213 13219 20247
rect 14473 20213 14507 20247
rect 15163 20213 15197 20247
rect 15577 20213 15611 20247
rect 7297 20009 7331 20043
rect 8723 20009 8757 20043
rect 9137 20009 9171 20043
rect 10609 20009 10643 20043
rect 11575 20009 11609 20043
rect 13277 20009 13311 20043
rect 14105 20009 14139 20043
rect 15853 20009 15887 20043
rect 5549 19941 5583 19975
rect 6698 19941 6732 19975
rect 10010 19941 10044 19975
rect 16221 19941 16255 19975
rect 16773 19941 16807 19975
rect 17785 19941 17819 19975
rect 1409 19873 1443 19907
rect 2973 19873 3007 19907
rect 5089 19873 5123 19907
rect 5273 19873 5307 19907
rect 5825 19873 5859 19907
rect 8652 19873 8686 19907
rect 11504 19873 11538 19907
rect 13829 19873 13863 19907
rect 19200 19873 19234 19907
rect 6377 19805 6411 19839
rect 9689 19805 9723 19839
rect 12909 19805 12943 19839
rect 16129 19805 16163 19839
rect 17693 19805 17727 19839
rect 17969 19805 18003 19839
rect 1547 19669 1581 19703
rect 3157 19669 3191 19703
rect 7757 19669 7791 19703
rect 12541 19669 12575 19703
rect 19303 19669 19337 19703
rect 1593 19465 1627 19499
rect 4721 19465 4755 19499
rect 10425 19465 10459 19499
rect 10701 19465 10735 19499
rect 15853 19465 15887 19499
rect 16221 19465 16255 19499
rect 16589 19465 16623 19499
rect 24777 19465 24811 19499
rect 8677 19397 8711 19431
rect 11529 19397 11563 19431
rect 17693 19397 17727 19431
rect 5917 19329 5951 19363
rect 7021 19329 7055 19363
rect 12173 19329 12207 19363
rect 20085 19329 20119 19363
rect 1409 19261 1443 19295
rect 2672 19261 2706 19295
rect 3617 19261 3651 19295
rect 4077 19261 4111 19295
rect 5089 19261 5123 19295
rect 5273 19261 5307 19295
rect 5641 19261 5675 19295
rect 7757 19261 7791 19295
rect 9505 19261 9539 19295
rect 11345 19261 11379 19295
rect 12541 19261 12575 19295
rect 13461 19261 13495 19295
rect 14933 19261 14967 19295
rect 16732 19261 16766 19295
rect 17141 19261 17175 19295
rect 18096 19261 18130 19295
rect 18521 19261 18555 19295
rect 19099 19261 19133 19295
rect 24593 19261 24627 19295
rect 25145 19261 25179 19295
rect 2053 19193 2087 19227
rect 3157 19193 3191 19227
rect 4353 19193 4387 19227
rect 8953 19193 8987 19227
rect 9826 19193 9860 19227
rect 13829 19193 13863 19227
rect 16819 19193 16853 19227
rect 19533 19193 19567 19227
rect 2513 19125 2547 19159
rect 2743 19125 2777 19159
rect 3433 19125 3467 19159
rect 6377 19125 6411 19159
rect 7573 19125 7607 19159
rect 8125 19125 8159 19159
rect 9413 19125 9447 19159
rect 11161 19125 11195 19159
rect 11897 19125 11931 19159
rect 12909 19125 12943 19159
rect 14105 19125 14139 19159
rect 14841 19125 14875 19159
rect 15301 19125 15335 19159
rect 18199 19125 18233 19159
rect 19257 19125 19291 19159
rect 19901 19125 19935 19159
rect 8493 18921 8527 18955
rect 9413 18921 9447 18955
rect 12449 18921 12483 18955
rect 13185 18921 13219 18955
rect 13737 18921 13771 18955
rect 16221 18921 16255 18955
rect 16589 18921 16623 18955
rect 17141 18921 17175 18955
rect 18061 18921 18095 18955
rect 24777 18921 24811 18955
rect 4905 18853 4939 18887
rect 6101 18853 6135 18887
rect 10333 18853 10367 18887
rect 10885 18853 10919 18887
rect 15622 18853 15656 18887
rect 1869 18785 1903 18819
rect 3008 18785 3042 18819
rect 5365 18785 5399 18819
rect 5825 18785 5859 18819
rect 7021 18785 7055 18819
rect 7389 18785 7423 18819
rect 11713 18785 11747 18819
rect 17049 18785 17083 18819
rect 17509 18785 17543 18819
rect 18680 18785 18714 18819
rect 19660 18785 19694 18819
rect 24593 18785 24627 18819
rect 4077 18717 4111 18751
rect 7665 18717 7699 18751
rect 8493 18717 8527 18751
rect 10241 18717 10275 18751
rect 12817 18717 12851 18751
rect 15301 18717 15335 18751
rect 20913 18717 20947 18751
rect 2099 18649 2133 18683
rect 11253 18649 11287 18683
rect 19763 18649 19797 18683
rect 1593 18581 1627 18615
rect 3111 18581 3145 18615
rect 3709 18581 3743 18615
rect 5273 18581 5307 18615
rect 8033 18581 8067 18615
rect 8723 18581 8757 18615
rect 9873 18581 9907 18615
rect 11851 18581 11885 18615
rect 14105 18581 14139 18615
rect 14933 18581 14967 18615
rect 18751 18581 18785 18615
rect 2053 18377 2087 18411
rect 2513 18377 2547 18411
rect 5089 18377 5123 18411
rect 7021 18377 7055 18411
rect 9045 18377 9079 18411
rect 12081 18377 12115 18411
rect 12173 18377 12207 18411
rect 13461 18377 13495 18411
rect 15761 18377 15795 18411
rect 17049 18377 17083 18411
rect 19073 18377 19107 18411
rect 20085 18377 20119 18411
rect 3065 18309 3099 18343
rect 6561 18309 6595 18343
rect 4353 18241 4387 18275
rect 8033 18241 8067 18275
rect 10333 18241 10367 18275
rect 11529 18241 11563 18275
rect 14749 18241 14783 18275
rect 16037 18241 16071 18275
rect 16497 18241 16531 18275
rect 1660 18173 1694 18207
rect 3525 18173 3559 18207
rect 3617 18173 3651 18207
rect 4077 18173 4111 18207
rect 5181 18173 5215 18207
rect 5733 18173 5767 18207
rect 9229 18173 9263 18207
rect 9689 18173 9723 18207
rect 10793 18173 10827 18207
rect 11345 18173 11379 18207
rect 12081 18173 12115 18207
rect 12449 18173 12483 18207
rect 12909 18173 12943 18207
rect 13921 18173 13955 18207
rect 14013 18173 14047 18207
rect 14473 18173 14507 18207
rect 18680 18173 18714 18207
rect 19441 18173 19475 18207
rect 19660 18173 19694 18207
rect 20453 18173 20487 18207
rect 5917 18105 5951 18139
rect 7389 18105 7423 18139
rect 7481 18105 7515 18139
rect 9965 18105 9999 18139
rect 13185 18105 13219 18139
rect 16129 18105 16163 18139
rect 19763 18105 19797 18139
rect 1731 18037 1765 18071
rect 2605 18037 2639 18071
rect 6285 18037 6319 18071
rect 8677 18037 8711 18071
rect 10701 18037 10735 18071
rect 11805 18037 11839 18071
rect 15393 18037 15427 18071
rect 17417 18037 17451 18071
rect 18751 18037 18785 18071
rect 20637 18037 20671 18071
rect 21649 18037 21683 18071
rect 24593 18037 24627 18071
rect 3709 17833 3743 17867
rect 5457 17833 5491 17867
rect 6377 17833 6411 17867
rect 6929 17833 6963 17867
rect 7389 17833 7423 17867
rect 10149 17833 10183 17867
rect 13093 17833 13127 17867
rect 16497 17833 16531 17867
rect 18429 17833 18463 17867
rect 7941 17765 7975 17799
rect 8493 17765 8527 17799
rect 10609 17765 10643 17799
rect 14289 17765 14323 17799
rect 16037 17765 16071 17799
rect 16865 17765 16899 17799
rect 1961 17697 1995 17731
rect 4721 17697 4755 17731
rect 4997 17697 5031 17731
rect 11989 17697 12023 17731
rect 12449 17697 12483 17731
rect 13829 17697 13863 17731
rect 14105 17697 14139 17731
rect 15644 17697 15678 17731
rect 16589 17697 16623 17731
rect 18613 17697 18647 17731
rect 18797 17697 18831 17731
rect 20948 17697 20982 17731
rect 22268 17697 22302 17731
rect 23280 17697 23314 17731
rect 2973 17629 3007 17663
rect 5181 17629 5215 17663
rect 6009 17629 6043 17663
rect 7849 17629 7883 17663
rect 10517 17629 10551 17663
rect 10793 17629 10827 17663
rect 12541 17629 12575 17663
rect 15715 17561 15749 17595
rect 2145 17493 2179 17527
rect 4353 17493 4387 17527
rect 9321 17493 9355 17527
rect 14565 17493 14599 17527
rect 17509 17493 17543 17527
rect 18153 17493 18187 17527
rect 21051 17493 21085 17527
rect 22339 17493 22373 17527
rect 23351 17493 23385 17527
rect 1593 17289 1627 17323
rect 4537 17289 4571 17323
rect 7757 17289 7791 17323
rect 8033 17289 8067 17323
rect 11713 17289 11747 17323
rect 13921 17289 13955 17323
rect 17785 17289 17819 17323
rect 24777 17289 24811 17323
rect 2053 17221 2087 17255
rect 7849 17221 7883 17255
rect 17049 17221 17083 17255
rect 5733 17153 5767 17187
rect 6837 17153 6871 17187
rect 1409 17085 1443 17119
rect 2605 17085 2639 17119
rect 3684 17085 3718 17119
rect 4169 17085 4203 17119
rect 8585 17153 8619 17187
rect 10425 17153 10459 17187
rect 13553 17153 13587 17187
rect 14381 17153 14415 17187
rect 16129 17153 16163 17187
rect 20775 17153 20809 17187
rect 21097 17153 21131 17187
rect 22109 17153 22143 17187
rect 12817 17085 12851 17119
rect 13277 17085 13311 17119
rect 15669 17085 15703 17119
rect 19660 17085 19694 17119
rect 20085 17085 20119 17119
rect 20672 17085 20706 17119
rect 21465 17085 21499 17119
rect 21700 17085 21734 17119
rect 22569 17085 22603 17119
rect 24593 17085 24627 17119
rect 25145 17085 25179 17119
rect 3893 17017 3927 17051
rect 4721 17017 4755 17051
rect 4813 17017 4847 17051
rect 5365 17017 5399 17051
rect 7158 17017 7192 17051
rect 7849 17017 7883 17051
rect 8906 17017 8940 17051
rect 10517 17017 10551 17051
rect 11069 17017 11103 17051
rect 14702 17017 14736 17051
rect 16037 17017 16071 17051
rect 16450 17017 16484 17051
rect 17325 17017 17359 17051
rect 18153 17017 18187 17051
rect 18245 17017 18279 17051
rect 18797 17017 18831 17051
rect 21787 17017 21821 17051
rect 2329 16949 2363 16983
rect 2789 16949 2823 16983
rect 3065 16949 3099 16983
rect 6009 16949 6043 16983
rect 6561 16949 6595 16983
rect 8401 16949 8435 16983
rect 9505 16949 9539 16983
rect 9873 16949 9907 16983
rect 10241 16949 10275 16983
rect 11989 16949 12023 16983
rect 12725 16949 12759 16983
rect 14197 16949 14231 16983
rect 15301 16949 15335 16983
rect 19073 16949 19107 16983
rect 19763 16949 19797 16983
rect 23305 16949 23339 16983
rect 4997 16745 5031 16779
rect 6837 16745 6871 16779
rect 7573 16745 7607 16779
rect 8677 16745 8711 16779
rect 10701 16745 10735 16779
rect 14381 16745 14415 16779
rect 16681 16745 16715 16779
rect 18613 16745 18647 16779
rect 21097 16745 21131 16779
rect 4439 16677 4473 16711
rect 5273 16677 5307 16711
rect 6009 16677 6043 16711
rect 7849 16677 7883 16711
rect 9781 16677 9815 16711
rect 9873 16677 9907 16711
rect 11437 16677 11471 16711
rect 13547 16677 13581 16711
rect 15761 16677 15795 16711
rect 17785 16677 17819 16711
rect 19349 16677 19383 16711
rect 19901 16677 19935 16711
rect 1961 16609 1995 16643
rect 3040 16609 3074 16643
rect 20980 16609 21014 16643
rect 21992 16609 22026 16643
rect 22937 16609 22971 16643
rect 25028 16609 25062 16643
rect 4077 16541 4111 16575
rect 5917 16541 5951 16575
rect 7757 16541 7791 16575
rect 10057 16541 10091 16575
rect 11345 16541 11379 16575
rect 11713 16541 11747 16575
rect 13185 16541 13219 16575
rect 15117 16541 15151 16575
rect 15669 16541 15703 16575
rect 17509 16541 17543 16575
rect 17693 16541 17727 16575
rect 17969 16541 18003 16575
rect 19257 16541 19291 16575
rect 23949 16541 23983 16575
rect 6469 16473 6503 16507
rect 8309 16473 8343 16507
rect 16221 16473 16255 16507
rect 22063 16473 22097 16507
rect 2145 16405 2179 16439
rect 3111 16405 3145 16439
rect 11161 16405 11195 16439
rect 12817 16405 12851 16439
rect 14105 16405 14139 16439
rect 23075 16405 23109 16439
rect 25099 16405 25133 16439
rect 1593 16201 1627 16235
rect 5089 16201 5123 16235
rect 5917 16201 5951 16235
rect 6193 16201 6227 16235
rect 6653 16201 6687 16235
rect 7205 16201 7239 16235
rect 7573 16201 7607 16235
rect 9045 16201 9079 16235
rect 9689 16201 9723 16235
rect 10793 16201 10827 16235
rect 14013 16201 14047 16235
rect 15669 16201 15703 16235
rect 15853 16201 15887 16235
rect 16129 16201 16163 16235
rect 17509 16201 17543 16235
rect 20637 16201 20671 16235
rect 21097 16201 21131 16235
rect 22017 16201 22051 16235
rect 24777 16201 24811 16235
rect 11253 16133 11287 16167
rect 15485 16133 15519 16167
rect 7757 16065 7791 16099
rect 8401 16065 8435 16099
rect 14749 16065 14783 16099
rect 14933 16065 14967 16099
rect 1409 15997 1443 16031
rect 2053 15997 2087 16031
rect 2513 15997 2547 16031
rect 2605 15997 2639 16031
rect 3065 15997 3099 16031
rect 4169 15997 4203 16031
rect 9873 15997 9907 16031
rect 13093 15997 13127 16031
rect 14289 15997 14323 16031
rect 15669 15997 15703 16031
rect 17785 16133 17819 16167
rect 21327 16133 21361 16167
rect 16497 16065 16531 16099
rect 16773 16065 16807 16099
rect 18153 16065 18187 16099
rect 19717 16065 19751 16099
rect 19993 16065 20027 16099
rect 22339 16065 22373 16099
rect 16221 15997 16255 16031
rect 21256 15997 21290 16031
rect 22236 15997 22270 16031
rect 24593 15997 24627 16031
rect 25145 15997 25179 16031
rect 3341 15929 3375 15963
rect 7849 15929 7883 15963
rect 9321 15929 9355 15963
rect 10194 15929 10228 15963
rect 12173 15929 12207 15963
rect 12909 15929 12943 15963
rect 13414 15929 13448 15963
rect 15025 15929 15059 15963
rect 16129 15929 16163 15963
rect 16589 15929 16623 15963
rect 18245 15929 18279 15963
rect 18797 15929 18831 15963
rect 19441 15929 19475 15963
rect 19809 15929 19843 15963
rect 3617 15861 3651 15895
rect 4077 15861 4111 15895
rect 4537 15861 4571 15895
rect 5365 15861 5399 15895
rect 11621 15861 11655 15895
rect 19073 15861 19107 15895
rect 21741 15861 21775 15895
rect 22937 15861 22971 15895
rect 25513 15861 25547 15895
rect 1593 15657 1627 15691
rect 3157 15657 3191 15691
rect 4629 15657 4663 15691
rect 7481 15657 7515 15691
rect 9413 15657 9447 15691
rect 12541 15657 12575 15691
rect 13369 15657 13403 15691
rect 14933 15657 14967 15691
rect 16497 15657 16531 15691
rect 18245 15657 18279 15691
rect 18613 15657 18647 15691
rect 19717 15657 19751 15691
rect 24823 15657 24857 15691
rect 4261 15589 4295 15623
rect 6923 15589 6957 15623
rect 8125 15589 8159 15623
rect 8723 15589 8757 15623
rect 12173 15589 12207 15623
rect 15485 15589 15519 15623
rect 17325 15589 17359 15623
rect 17877 15589 17911 15623
rect 18889 15589 18923 15623
rect 19441 15589 19475 15623
rect 21281 15589 21315 15623
rect 1409 15521 1443 15555
rect 2973 15521 3007 15555
rect 5089 15521 5123 15555
rect 5549 15521 5583 15555
rect 5733 15521 5767 15555
rect 8585 15521 8619 15555
rect 9873 15521 9907 15555
rect 10333 15521 10367 15555
rect 11437 15521 11471 15555
rect 11897 15521 11931 15555
rect 22728 15521 22762 15555
rect 23740 15521 23774 15555
rect 24752 15521 24786 15555
rect 2053 15453 2087 15487
rect 6561 15453 6595 15487
rect 10609 15453 10643 15487
rect 13001 15453 13035 15487
rect 15393 15453 15427 15487
rect 15669 15453 15703 15487
rect 17222 15453 17256 15487
rect 18797 15453 18831 15487
rect 21189 15453 21223 15487
rect 21465 15453 21499 15487
rect 22109 15453 22143 15487
rect 22799 15385 22833 15419
rect 2605 15317 2639 15351
rect 3709 15317 3743 15351
rect 6377 15317 6411 15351
rect 7849 15317 7883 15351
rect 12817 15317 12851 15351
rect 13921 15317 13955 15351
rect 23811 15317 23845 15351
rect 2145 15113 2179 15147
rect 3065 15113 3099 15147
rect 3433 15113 3467 15147
rect 4721 15113 4755 15147
rect 6193 15113 6227 15147
rect 6469 15113 6503 15147
rect 6561 15113 6595 15147
rect 8033 15113 8067 15147
rect 9873 15113 9907 15147
rect 10609 15113 10643 15147
rect 12587 15113 12621 15147
rect 13277 15113 13311 15147
rect 14749 15113 14783 15147
rect 16773 15113 16807 15147
rect 19073 15113 19107 15147
rect 21465 15113 21499 15147
rect 22109 15113 22143 15147
rect 22845 15113 22879 15147
rect 23121 15113 23155 15147
rect 25145 15113 25179 15147
rect 2421 15045 2455 15079
rect 2743 15045 2777 15079
rect 4353 14977 4387 15011
rect 5917 14977 5951 15011
rect 1593 14909 1627 14943
rect 2672 14909 2706 14943
rect 3617 14909 3651 14943
rect 4077 14909 4111 14943
rect 5181 14909 5215 14943
rect 5641 14909 5675 14943
rect 10241 15045 10275 15079
rect 11805 15045 11839 15079
rect 19441 15045 19475 15079
rect 21741 15045 21775 15079
rect 6837 14977 6871 15011
rect 8953 14977 8987 15011
rect 11529 14977 11563 15011
rect 13829 14977 13863 15011
rect 14105 14977 14139 15011
rect 15853 14977 15887 15011
rect 17785 14977 17819 15011
rect 18153 14977 18187 15011
rect 18797 14977 18831 15011
rect 10793 14909 10827 14943
rect 11253 14909 11287 14943
rect 12173 14909 12207 14943
rect 12516 14909 12550 14943
rect 17024 14909 17058 14943
rect 20361 14909 20395 14943
rect 20545 14909 20579 14943
rect 22360 14909 22394 14943
rect 23740 14909 23774 14943
rect 24133 14909 24167 14943
rect 6469 14841 6503 14875
rect 7158 14841 7192 14875
rect 8677 14841 8711 14875
rect 8769 14841 8803 14875
rect 13921 14841 13955 14875
rect 15393 14841 15427 14875
rect 15485 14841 15519 14875
rect 18245 14841 18279 14875
rect 20866 14841 20900 14875
rect 24685 14841 24719 14875
rect 1777 14773 1811 14807
rect 5089 14773 5123 14807
rect 7757 14773 7791 14807
rect 8493 14773 8527 14807
rect 13001 14773 13035 14807
rect 15209 14773 15243 14807
rect 16405 14773 16439 14807
rect 17095 14773 17129 14807
rect 17509 14773 17543 14807
rect 22431 14773 22465 14807
rect 23811 14773 23845 14807
rect 24501 14773 24535 14807
rect 1593 14569 1627 14603
rect 3617 14569 3651 14603
rect 4169 14569 4203 14603
rect 8953 14569 8987 14603
rect 10793 14569 10827 14603
rect 13829 14569 13863 14603
rect 14197 14569 14231 14603
rect 15117 14569 15151 14603
rect 17233 14569 17267 14603
rect 19441 14569 19475 14603
rect 20637 14569 20671 14603
rect 22569 14569 22603 14603
rect 24777 14569 24811 14603
rect 3111 14501 3145 14535
rect 7757 14501 7791 14535
rect 8585 14501 8619 14535
rect 11989 14501 12023 14535
rect 13001 14501 13035 14535
rect 13553 14501 13587 14535
rect 15485 14501 15519 14535
rect 17601 14501 17635 14535
rect 17693 14501 17727 14535
rect 21097 14501 21131 14535
rect 1409 14433 1443 14467
rect 3008 14433 3042 14467
rect 4077 14433 4111 14467
rect 4537 14433 4571 14467
rect 5181 14433 5215 14467
rect 5549 14433 5583 14467
rect 6101 14433 6135 14467
rect 6285 14433 6319 14467
rect 9873 14433 9907 14467
rect 10149 14433 10183 14467
rect 11253 14433 11287 14467
rect 11713 14433 11747 14467
rect 22477 14433 22511 14467
rect 23029 14433 23063 14467
rect 24593 14433 24627 14467
rect 6377 14365 6411 14399
rect 7665 14365 7699 14399
rect 8309 14365 8343 14399
rect 10425 14365 10459 14399
rect 12909 14365 12943 14399
rect 15393 14365 15427 14399
rect 15669 14365 15703 14399
rect 19073 14365 19107 14399
rect 21005 14365 21039 14399
rect 21465 14365 21499 14399
rect 18153 14297 18187 14331
rect 22293 14297 22327 14331
rect 7205 14229 7239 14263
rect 9505 14229 9539 14263
rect 19993 14229 20027 14263
rect 21925 14229 21959 14263
rect 23673 14229 23707 14263
rect 1777 14025 1811 14059
rect 5641 14025 5675 14059
rect 6377 14025 6411 14059
rect 8125 14025 8159 14059
rect 9781 14025 9815 14059
rect 13369 14025 13403 14059
rect 13645 14025 13679 14059
rect 14013 14025 14047 14059
rect 14841 14025 14875 14059
rect 14933 14025 14967 14059
rect 16865 14025 16899 14059
rect 20913 14025 20947 14059
rect 22477 14025 22511 14059
rect 24777 14025 24811 14059
rect 8815 13957 8849 13991
rect 11713 13957 11747 13991
rect 15761 13957 15795 13991
rect 2697 13889 2731 13923
rect 4169 13889 4203 13923
rect 5365 13889 5399 13923
rect 7481 13889 7515 13923
rect 12449 13889 12483 13923
rect 14841 13889 14875 13923
rect 16129 13889 16163 13923
rect 19901 13889 19935 13923
rect 20177 13889 20211 13923
rect 21465 13889 21499 13923
rect 21741 13889 21775 13923
rect 1869 13821 1903 13855
rect 2881 13821 2915 13855
rect 4537 13821 4571 13855
rect 4905 13821 4939 13855
rect 5181 13821 5215 13855
rect 8712 13821 8746 13855
rect 16992 13821 17026 13855
rect 17417 13821 17451 13855
rect 19073 13821 19107 13855
rect 23673 13821 23707 13855
rect 24087 13821 24121 13855
rect 25304 13821 25338 13855
rect 25697 13821 25731 13855
rect 2421 13753 2455 13787
rect 3243 13753 3277 13787
rect 6101 13753 6135 13787
rect 7205 13753 7239 13787
rect 7297 13753 7331 13787
rect 10057 13753 10091 13787
rect 10149 13753 10183 13787
rect 10701 13753 10735 13787
rect 11253 13753 11287 13787
rect 12770 13753 12804 13787
rect 14657 13753 14691 13787
rect 15209 13753 15243 13787
rect 15301 13753 15335 13787
rect 17095 13753 17129 13787
rect 18153 13753 18187 13787
rect 18245 13753 18279 13787
rect 18797 13753 18831 13787
rect 19717 13753 19751 13787
rect 19993 13753 20027 13787
rect 21557 13753 21591 13787
rect 2053 13685 2087 13719
rect 3801 13685 3835 13719
rect 9229 13685 9263 13719
rect 12173 13685 12207 13719
rect 17877 13685 17911 13719
rect 22937 13685 22971 13719
rect 23489 13685 23523 13719
rect 23765 13685 23799 13719
rect 25375 13685 25409 13719
rect 3893 13481 3927 13515
rect 4445 13481 4479 13515
rect 6193 13481 6227 13515
rect 6653 13481 6687 13515
rect 7205 13481 7239 13515
rect 11621 13481 11655 13515
rect 12449 13481 12483 13515
rect 13001 13481 13035 13515
rect 13553 13481 13587 13515
rect 17877 13481 17911 13515
rect 18245 13481 18279 13515
rect 19901 13481 19935 13515
rect 20729 13481 20763 13515
rect 2421 13413 2455 13447
rect 8217 13413 8251 13447
rect 8769 13413 8803 13447
rect 10010 13413 10044 13447
rect 15485 13413 15519 13447
rect 17049 13413 17083 13447
rect 18613 13413 18647 13447
rect 19165 13413 19199 13447
rect 19533 13413 19567 13447
rect 21557 13413 21591 13447
rect 23121 13413 23155 13447
rect 6285 13345 6319 13379
rect 10609 13345 10643 13379
rect 11437 13345 11471 13379
rect 24552 13345 24586 13379
rect 2329 13277 2363 13311
rect 2605 13277 2639 13311
rect 4077 13277 4111 13311
rect 8125 13277 8159 13311
rect 9045 13277 9079 13311
rect 9689 13277 9723 13311
rect 12633 13277 12667 13311
rect 15393 13277 15427 13311
rect 16957 13277 16991 13311
rect 17233 13277 17267 13311
rect 18521 13277 18555 13311
rect 21465 13277 21499 13311
rect 21741 13277 21775 13311
rect 23029 13277 23063 13311
rect 24639 13277 24673 13311
rect 9505 13209 9539 13243
rect 15117 13209 15151 13243
rect 15945 13209 15979 13243
rect 23581 13209 23615 13243
rect 1593 13141 1627 13175
rect 3249 13141 3283 13175
rect 4997 13141 5031 13175
rect 7573 13141 7607 13175
rect 7941 13141 7975 13175
rect 13829 13141 13863 13175
rect 21097 13141 21131 13175
rect 1685 12937 1719 12971
rect 1961 12937 1995 12971
rect 2697 12937 2731 12971
rect 3709 12937 3743 12971
rect 4813 12937 4847 12971
rect 5457 12937 5491 12971
rect 7757 12937 7791 12971
rect 8125 12937 8159 12971
rect 11483 12937 11517 12971
rect 13277 12937 13311 12971
rect 13369 12937 13403 12971
rect 14933 12937 14967 12971
rect 15209 12937 15243 12971
rect 15393 12937 15427 12971
rect 22017 12937 22051 12971
rect 22477 12937 22511 12971
rect 24961 12937 24995 12971
rect 2973 12869 3007 12903
rect 4445 12869 4479 12903
rect 8769 12869 8803 12903
rect 12679 12869 12713 12903
rect 3893 12801 3927 12835
rect 5181 12801 5215 12835
rect 5457 12801 5491 12835
rect 6285 12801 6319 12835
rect 9873 12801 9907 12835
rect 11161 12801 11195 12835
rect 1777 12733 1811 12767
rect 2329 12733 2363 12767
rect 2789 12733 2823 12767
rect 5733 12733 5767 12767
rect 6837 12733 6871 12767
rect 8585 12733 8619 12767
rect 9045 12733 9079 12767
rect 11412 12733 11446 12767
rect 12608 12733 12642 12767
rect 3985 12665 4019 12699
rect 5641 12665 5675 12699
rect 7158 12665 7192 12699
rect 9965 12665 9999 12699
rect 10517 12665 10551 12699
rect 13645 12801 13679 12835
rect 14105 12801 14139 12835
rect 13737 12665 13771 12699
rect 25191 12869 25225 12903
rect 25605 12869 25639 12903
rect 15853 12801 15887 12835
rect 16129 12801 16163 12835
rect 18337 12801 18371 12835
rect 18981 12801 19015 12835
rect 20361 12801 20395 12835
rect 23121 12801 23155 12835
rect 19876 12733 19910 12767
rect 20821 12733 20855 12767
rect 22636 12733 22670 12767
rect 24108 12733 24142 12767
rect 25120 12733 25154 12767
rect 15945 12665 15979 12699
rect 18429 12665 18463 12699
rect 21183 12665 21217 12699
rect 23397 12665 23431 12699
rect 3341 12597 3375 12631
rect 5917 12597 5951 12631
rect 8493 12597 8527 12631
rect 9597 12597 9631 12631
rect 10793 12597 10827 12631
rect 11897 12597 11931 12631
rect 12173 12597 12207 12631
rect 13001 12597 13035 12631
rect 13277 12597 13311 12631
rect 14565 12597 14599 12631
rect 15209 12597 15243 12631
rect 16865 12597 16899 12631
rect 17233 12597 17267 12631
rect 17877 12597 17911 12631
rect 19257 12597 19291 12631
rect 19947 12597 19981 12631
rect 20729 12597 20763 12631
rect 21741 12597 21775 12631
rect 22707 12597 22741 12631
rect 24179 12597 24213 12631
rect 24593 12597 24627 12631
rect 4169 12393 4203 12427
rect 6929 12393 6963 12427
rect 9873 12393 9907 12427
rect 10241 12393 10275 12427
rect 12449 12393 12483 12427
rect 13461 12393 13495 12427
rect 13737 12393 13771 12427
rect 16405 12393 16439 12427
rect 18153 12393 18187 12427
rect 18521 12393 18555 12427
rect 21281 12393 21315 12427
rect 21833 12393 21867 12427
rect 22109 12393 22143 12427
rect 6377 12325 6411 12359
rect 7205 12325 7239 12359
rect 8769 12325 8803 12359
rect 10701 12325 10735 12359
rect 12862 12325 12896 12359
rect 15485 12325 15519 12359
rect 16037 12325 16071 12359
rect 17554 12325 17588 12359
rect 18797 12325 18831 12359
rect 19441 12325 19475 12359
rect 22753 12325 22787 12359
rect 22845 12325 22879 12359
rect 1409 12257 1443 12291
rect 2697 12257 2731 12291
rect 2881 12257 2915 12291
rect 4077 12257 4111 12291
rect 4629 12257 4663 12291
rect 5641 12257 5675 12291
rect 6101 12257 6135 12291
rect 8309 12257 8343 12291
rect 8585 12257 8619 12291
rect 19993 12257 20027 12291
rect 24501 12257 24535 12291
rect 24685 12257 24719 12291
rect 3157 12189 3191 12223
rect 3893 12189 3927 12223
rect 10609 12189 10643 12223
rect 10977 12189 11011 12223
rect 12541 12189 12575 12223
rect 15393 12189 15427 12223
rect 17233 12189 17267 12223
rect 19349 12189 19383 12223
rect 20913 12189 20947 12223
rect 23029 12189 23063 12223
rect 24777 12189 24811 12223
rect 1593 12121 1627 12155
rect 1961 12053 1995 12087
rect 2237 12053 2271 12087
rect 5089 12053 5123 12087
rect 7941 12053 7975 12087
rect 14197 12053 14231 12087
rect 20729 12053 20763 12087
rect 23673 12053 23707 12087
rect 2237 11849 2271 11883
rect 3249 11849 3283 11883
rect 5641 11849 5675 11883
rect 7021 11849 7055 11883
rect 8953 11849 8987 11883
rect 10609 11849 10643 11883
rect 11161 11849 11195 11883
rect 16957 11849 16991 11883
rect 21649 11849 21683 11883
rect 22293 11849 22327 11883
rect 24685 11849 24719 11883
rect 8493 11781 8527 11815
rect 11529 11781 11563 11815
rect 18429 11781 18463 11815
rect 19809 11781 19843 11815
rect 22615 11781 22649 11815
rect 25421 11781 25455 11815
rect 2881 11713 2915 11747
rect 4813 11713 4847 11747
rect 9597 11713 9631 11747
rect 10609 11713 10643 11747
rect 13553 11713 13587 11747
rect 14105 11713 14139 11747
rect 15945 11713 15979 11747
rect 16221 11713 16255 11747
rect 20729 11713 20763 11747
rect 22937 11713 22971 11747
rect 2329 11645 2363 11679
rect 3341 11645 3375 11679
rect 4353 11645 4387 11679
rect 4445 11645 4479 11679
rect 4629 11645 4663 11679
rect 6837 11645 6871 11679
rect 7297 11645 7331 11679
rect 11345 11645 11379 11679
rect 11805 11645 11839 11679
rect 12817 11645 12851 11679
rect 13001 11645 13035 11679
rect 15025 11645 15059 11679
rect 15669 11645 15703 11679
rect 18889 11645 18923 11679
rect 21925 11645 21959 11679
rect 22544 11645 22578 11679
rect 23673 11645 23707 11679
rect 24133 11645 24167 11679
rect 25237 11645 25271 11679
rect 25789 11645 25823 11679
rect 3801 11577 3835 11611
rect 6101 11577 6135 11611
rect 7941 11577 7975 11611
rect 8033 11577 8067 11611
rect 9918 11577 9952 11611
rect 12173 11577 12207 11611
rect 13277 11577 13311 11611
rect 14426 11577 14460 11611
rect 16037 11577 16071 11611
rect 18705 11577 18739 11611
rect 19210 11577 19244 11611
rect 20177 11577 20211 11611
rect 20545 11577 20579 11611
rect 21050 11577 21084 11611
rect 23397 11577 23431 11611
rect 23489 11577 23523 11611
rect 1593 11509 1627 11543
rect 2513 11509 2547 11543
rect 3525 11509 3559 11543
rect 4261 11509 4295 11543
rect 7665 11509 7699 11543
rect 9413 11509 9447 11543
rect 10517 11509 10551 11543
rect 10885 11509 10919 11543
rect 14013 11509 14047 11543
rect 15301 11509 15335 11543
rect 17233 11509 17267 11543
rect 17693 11509 17727 11543
rect 23765 11509 23799 11543
rect 25145 11509 25179 11543
rect 1593 11305 1627 11339
rect 4905 11305 4939 11339
rect 7941 11305 7975 11339
rect 8493 11305 8527 11339
rect 12817 11305 12851 11339
rect 13093 11305 13127 11339
rect 13737 11305 13771 11339
rect 14289 11305 14323 11339
rect 18245 11305 18279 11339
rect 18613 11305 18647 11339
rect 20453 11305 20487 11339
rect 21005 11305 21039 11339
rect 22661 11305 22695 11339
rect 24961 11305 24995 11339
rect 3801 11237 3835 11271
rect 7389 11237 7423 11271
rect 10885 11237 10919 11271
rect 15025 11237 15059 11271
rect 15669 11237 15703 11271
rect 17646 11237 17680 11271
rect 19993 11237 20027 11271
rect 23489 11237 23523 11271
rect 1409 11169 1443 11203
rect 2421 11169 2455 11203
rect 2697 11169 2731 11203
rect 4261 11169 4295 11203
rect 4445 11169 4479 11203
rect 4721 11169 4755 11203
rect 6009 11169 6043 11203
rect 6469 11169 6503 11203
rect 9689 11169 9723 11203
rect 12265 11169 12299 11203
rect 13369 11169 13403 11203
rect 19441 11169 19475 11203
rect 19717 11169 19751 11203
rect 20913 11169 20947 11203
rect 21373 11169 21407 11203
rect 25145 11169 25179 11203
rect 25329 11169 25363 11203
rect 2881 11101 2915 11135
rect 6745 11101 6779 11135
rect 7573 11101 7607 11135
rect 10793 11101 10827 11135
rect 15577 11101 15611 11135
rect 17325 11101 17359 11135
rect 23397 11101 23431 11135
rect 2513 11033 2547 11067
rect 3525 11033 3559 11067
rect 4537 11033 4571 11067
rect 11345 11033 11379 11067
rect 12173 11033 12207 11067
rect 16129 11033 16163 11067
rect 23949 11033 23983 11067
rect 1869 10965 1903 10999
rect 2329 10965 2363 10999
rect 9873 10965 9907 10999
rect 12449 10965 12483 10999
rect 18981 10965 19015 10999
rect 22109 10965 22143 10999
rect 24317 10965 24351 10999
rect 1685 10761 1719 10795
rect 3249 10761 3283 10795
rect 3433 10761 3467 10795
rect 5549 10761 5583 10795
rect 6561 10761 6595 10795
rect 7205 10761 7239 10795
rect 7665 10761 7699 10795
rect 9137 10761 9171 10795
rect 10517 10761 10551 10795
rect 10885 10761 10919 10795
rect 11253 10761 11287 10795
rect 12173 10761 12207 10795
rect 15945 10761 15979 10795
rect 21557 10761 21591 10795
rect 21833 10761 21867 10795
rect 25513 10761 25547 10795
rect 2329 10693 2363 10727
rect 2973 10625 3007 10659
rect 2237 10557 2271 10591
rect 2513 10557 2547 10591
rect 6285 10693 6319 10727
rect 8401 10693 8435 10727
rect 15485 10693 15519 10727
rect 20269 10693 20303 10727
rect 7849 10625 7883 10659
rect 8769 10625 8803 10659
rect 13185 10625 13219 10659
rect 24041 10625 24075 10659
rect 25697 10625 25731 10659
rect 3709 10557 3743 10591
rect 4353 10557 4387 10591
rect 5733 10557 5767 10591
rect 9321 10557 9355 10591
rect 11069 10557 11103 10591
rect 11529 10557 11563 10591
rect 14289 10557 14323 10591
rect 16313 10557 16347 10591
rect 16497 10557 16531 10591
rect 17877 10557 17911 10591
rect 18337 10557 18371 10591
rect 18521 10557 18555 10591
rect 20453 10557 20487 10591
rect 20913 10557 20947 10591
rect 22201 10557 22235 10591
rect 22477 10557 22511 10591
rect 25304 10557 25338 10591
rect 26065 10557 26099 10591
rect 2145 10489 2179 10523
rect 3433 10489 3467 10523
rect 7941 10489 7975 10523
rect 9642 10489 9676 10523
rect 12541 10489 12575 10523
rect 12633 10489 12667 10523
rect 13553 10489 13587 10523
rect 14610 10489 14644 10523
rect 21189 10489 21223 10523
rect 23765 10489 23799 10523
rect 23857 10489 23891 10523
rect 4077 10421 4111 10455
rect 4813 10421 4847 10455
rect 5181 10421 5215 10455
rect 5917 10421 5951 10455
rect 10241 10421 10275 10455
rect 14197 10421 14231 10455
rect 15209 10421 15243 10455
rect 16129 10421 16163 10455
rect 17325 10421 17359 10455
rect 18153 10421 18187 10455
rect 19257 10421 19291 10455
rect 19717 10421 19751 10455
rect 22109 10421 22143 10455
rect 23029 10421 23063 10455
rect 23397 10421 23431 10455
rect 24961 10421 24995 10455
rect 4353 10217 4387 10251
rect 7849 10217 7883 10251
rect 11253 10217 11287 10251
rect 12541 10217 12575 10251
rect 12909 10217 12943 10251
rect 14381 10217 14415 10251
rect 16313 10217 16347 10251
rect 17233 10217 17267 10251
rect 18429 10217 18463 10251
rect 18981 10217 19015 10251
rect 21741 10217 21775 10251
rect 22293 10217 22327 10251
rect 22845 10217 22879 10251
rect 949 10149 983 10183
rect 5549 10149 5583 10183
rect 8769 10149 8803 10183
rect 9321 10149 9355 10183
rect 10425 10149 10459 10183
rect 10977 10149 11011 10183
rect 13185 10149 13219 10183
rect 15117 10149 15151 10183
rect 17509 10149 17543 10183
rect 21051 10149 21085 10183
rect 23397 10149 23431 10183
rect 23857 10149 23891 10183
rect 24409 10149 24443 10183
rect 1409 10081 1443 10115
rect 2421 10081 2455 10115
rect 2697 10081 2731 10115
rect 3433 10081 3467 10115
rect 4813 10081 4847 10115
rect 5089 10081 5123 10115
rect 6377 10081 6411 10115
rect 6653 10081 6687 10115
rect 8033 10081 8067 10115
rect 8493 10081 8527 10115
rect 11989 10081 12023 10115
rect 15301 10081 15335 10115
rect 15761 10081 15795 10115
rect 19165 10081 19199 10115
rect 19441 10081 19475 10115
rect 20821 10081 20855 10115
rect 25237 10081 25271 10115
rect 2881 10013 2915 10047
rect 7113 10013 7147 10047
rect 10333 10013 10367 10047
rect 13093 10013 13127 10047
rect 13553 10013 13587 10047
rect 15853 10013 15887 10047
rect 17417 10013 17451 10047
rect 21925 10013 21959 10047
rect 23765 10013 23799 10047
rect 2513 9945 2547 9979
rect 4721 9945 4755 9979
rect 4905 9945 4939 9979
rect 6285 9945 6319 9979
rect 6469 9945 6503 9979
rect 12127 9945 12161 9979
rect 17969 9945 18003 9979
rect 1593 9877 1627 9911
rect 1869 9877 1903 9911
rect 2329 9877 2363 9911
rect 3801 9877 3835 9911
rect 16681 9877 16715 9911
rect 19901 9877 19935 9911
rect 20545 9877 20579 9911
rect 25421 9877 25455 9911
rect 949 9673 983 9707
rect 1869 9673 1903 9707
rect 2237 9673 2271 9707
rect 2697 9673 2731 9707
rect 4721 9673 4755 9707
rect 6377 9673 6411 9707
rect 8033 9673 8067 9707
rect 8401 9673 8435 9707
rect 9689 9673 9723 9707
rect 10057 9673 10091 9707
rect 12909 9673 12943 9707
rect 15209 9673 15243 9707
rect 17233 9673 17267 9707
rect 17417 9673 17451 9707
rect 18245 9673 18279 9707
rect 18981 9673 19015 9707
rect 21189 9673 21223 9707
rect 22753 9673 22787 9707
rect 24685 9673 24719 9707
rect 26065 9673 26099 9707
rect 10793 9605 10827 9639
rect 11989 9605 12023 9639
rect 14105 9605 14139 9639
rect 1961 9537 1995 9571
rect 4905 9537 4939 9571
rect 5549 9537 5583 9571
rect 8677 9537 8711 9571
rect 10241 9537 10275 9571
rect 11161 9537 11195 9571
rect 13369 9537 13403 9571
rect 14933 9537 14967 9571
rect 19257 9537 19291 9571
rect 21833 9537 21867 9571
rect 24225 9537 24259 9571
rect 1740 9469 1774 9503
rect 3157 9469 3191 9503
rect 3617 9469 3651 9503
rect 4813 9469 4847 9503
rect 5089 9469 5123 9503
rect 6929 9469 6963 9503
rect 7481 9469 7515 9503
rect 15025 9469 15059 9503
rect 15485 9469 15519 9503
rect 17233 9469 17267 9503
rect 18061 9469 18095 9503
rect 18521 9469 18555 9503
rect 20177 9469 20211 9503
rect 20796 9469 20830 9503
rect 21557 9469 21591 9503
rect 25304 9469 25338 9503
rect 25697 9469 25731 9503
rect 1593 9401 1627 9435
rect 2973 9401 3007 9435
rect 6009 9401 6043 9435
rect 8769 9401 8803 9435
rect 9321 9401 9355 9435
rect 10333 9401 10367 9435
rect 13093 9401 13127 9435
rect 13185 9401 13219 9435
rect 16129 9401 16163 9435
rect 16221 9401 16255 9435
rect 16773 9401 16807 9435
rect 19349 9401 19383 9435
rect 19901 9401 19935 9435
rect 22154 9401 22188 9435
rect 23765 9401 23799 9435
rect 23857 9401 23891 9435
rect 25053 9401 25087 9435
rect 3249 9333 3283 9367
rect 4353 9333 4387 9367
rect 7021 9333 7055 9367
rect 15945 9333 15979 9367
rect 17693 9333 17727 9367
rect 20867 9333 20901 9367
rect 23029 9333 23063 9367
rect 23397 9333 23431 9367
rect 25375 9333 25409 9367
rect 1593 9129 1627 9163
rect 1961 9129 1995 9163
rect 2237 9129 2271 9163
rect 3525 9129 3559 9163
rect 3801 9129 3835 9163
rect 5825 9129 5859 9163
rect 7941 9129 7975 9163
rect 10701 9129 10735 9163
rect 12449 9129 12483 9163
rect 13553 9129 13587 9163
rect 13645 9129 13679 9163
rect 21557 9129 21591 9163
rect 22569 9129 22603 9163
rect 23673 9129 23707 9163
rect 24409 9129 24443 9163
rect 4077 9061 4111 9095
rect 9873 9061 9907 9095
rect 1409 8993 1443 9027
rect 2697 8993 2731 9027
rect 4445 8993 4479 9027
rect 5089 8993 5123 9027
rect 6101 8993 6135 9027
rect 6561 8993 6595 9027
rect 2421 8925 2455 8959
rect 6745 8925 6779 8959
rect 7573 8925 7607 8959
rect 9781 8925 9815 8959
rect 10057 8925 10091 8959
rect 12081 8925 12115 8959
rect 8493 8857 8527 8891
rect 13001 8857 13035 8891
rect 13369 8857 13403 8891
rect 15577 9061 15611 9095
rect 17141 9061 17175 9095
rect 18934 9061 18968 9095
rect 21970 9061 22004 9095
rect 14232 8993 14266 9027
rect 16129 8993 16163 9027
rect 18613 8993 18647 9027
rect 23213 8993 23247 9027
rect 23397 8993 23431 9027
rect 23857 8993 23891 9027
rect 25028 8993 25062 9027
rect 15485 8925 15519 8959
rect 17049 8925 17083 8959
rect 17325 8925 17359 8959
rect 21649 8925 21683 8959
rect 22845 8925 22879 8959
rect 14335 8857 14369 8891
rect 15025 8857 15059 8891
rect 25099 8857 25133 8891
rect 5457 8789 5491 8823
rect 7021 8789 7055 8823
rect 7481 8789 7515 8823
rect 8769 8789 8803 8823
rect 9229 8789 9263 8823
rect 13553 8789 13587 8823
rect 16405 8789 16439 8823
rect 19533 8789 19567 8823
rect 19809 8789 19843 8823
rect 21189 8789 21223 8823
rect 4813 8585 4847 8619
rect 6101 8585 6135 8619
rect 6469 8585 6503 8619
rect 7021 8585 7055 8619
rect 8493 8585 8527 8619
rect 8861 8585 8895 8619
rect 9137 8585 9171 8619
rect 11483 8585 11517 8619
rect 13369 8585 13403 8619
rect 14611 8585 14645 8619
rect 17049 8585 17083 8619
rect 18291 8585 18325 8619
rect 20269 8585 20303 8619
rect 23029 8585 23063 8619
rect 9965 8517 9999 8551
rect 11805 8517 11839 8551
rect 14289 8517 14323 8551
rect 17877 8517 17911 8551
rect 20085 8517 20119 8551
rect 25375 8517 25409 8551
rect 3157 8449 3191 8483
rect 5549 8449 5583 8483
rect 7573 8449 7607 8483
rect 10701 8449 10735 8483
rect 15485 8449 15519 8483
rect 19257 8449 19291 8483
rect 21833 8449 21867 8483
rect 24225 8449 24259 8483
rect 1685 8381 1719 8415
rect 4997 8381 5031 8415
rect 5457 8381 5491 8415
rect 11412 8381 11446 8415
rect 12449 8381 12483 8415
rect 14508 8381 14542 8415
rect 14933 8381 14967 8415
rect 18188 8381 18222 8415
rect 18613 8381 18647 8415
rect 20085 8381 20119 8415
rect 20780 8381 20814 8415
rect 21281 8381 21315 8415
rect 25304 8381 25338 8415
rect 3065 8313 3099 8347
rect 3478 8313 3512 8347
rect 9413 8313 9447 8347
rect 9505 8313 9539 8347
rect 12811 8313 12845 8347
rect 19349 8313 19383 8347
rect 19901 8313 19935 8347
rect 20867 8313 20901 8347
rect 22154 8313 22188 8347
rect 23397 8313 23431 8347
rect 23765 8313 23799 8347
rect 23857 8313 23891 8347
rect 2053 8245 2087 8279
rect 2697 8245 2731 8279
rect 4077 8245 4111 8279
rect 4445 8245 4479 8279
rect 7481 8245 7515 8279
rect 7941 8245 7975 8279
rect 10333 8245 10367 8279
rect 11253 8245 11287 8279
rect 12265 8245 12299 8279
rect 13737 8245 13771 8279
rect 15393 8245 15427 8279
rect 15853 8245 15887 8279
rect 16405 8245 16439 8279
rect 17325 8245 17359 8279
rect 18981 8245 19015 8279
rect 21649 8245 21683 8279
rect 22753 8245 22787 8279
rect 25053 8245 25087 8279
rect 25789 8245 25823 8279
rect 2053 8041 2087 8075
rect 3157 8041 3191 8075
rect 5825 8041 5859 8075
rect 11805 8041 11839 8075
rect 12357 8041 12391 8075
rect 15117 8041 15151 8075
rect 16129 8041 16163 8075
rect 17509 8041 17543 8075
rect 18429 8041 18463 8075
rect 19349 8041 19383 8075
rect 23489 8041 23523 8075
rect 2329 7973 2363 8007
rect 4261 7973 4295 8007
rect 6653 7973 6687 8007
rect 7665 7973 7699 8007
rect 10051 7973 10085 8007
rect 13829 7973 13863 8007
rect 15715 7973 15749 8007
rect 16951 7973 16985 8007
rect 22154 7973 22188 8007
rect 23765 7973 23799 8007
rect 8309 7905 8343 7939
rect 8493 7905 8527 7939
rect 8769 7905 8803 7939
rect 13001 7905 13035 7939
rect 15612 7905 15646 7939
rect 16589 7905 16623 7939
rect 18337 7905 18371 7939
rect 18797 7905 18831 7939
rect 25196 7905 25230 7939
rect 2237 7837 2271 7871
rect 2513 7837 2547 7871
rect 4169 7837 4203 7871
rect 4445 7837 4479 7871
rect 5181 7837 5215 7871
rect 6377 7837 6411 7871
rect 6561 7837 6595 7871
rect 9689 7837 9723 7871
rect 11437 7837 11471 7871
rect 13553 7837 13587 7871
rect 13737 7837 13771 7871
rect 21833 7837 21867 7871
rect 23673 7837 23707 7871
rect 25283 7837 25317 7871
rect 7113 7769 7147 7803
rect 9413 7769 9447 7803
rect 14289 7769 14323 7803
rect 21373 7769 21407 7803
rect 22753 7769 22787 7803
rect 24225 7769 24259 7803
rect 1685 7701 1719 7735
rect 3617 7701 3651 7735
rect 5457 7701 5491 7735
rect 10609 7701 10643 7735
rect 12633 7701 12667 7735
rect 21649 7701 21683 7735
rect 1731 7497 1765 7531
rect 3985 7497 4019 7531
rect 4353 7497 4387 7531
rect 5917 7497 5951 7531
rect 6285 7497 6319 7531
rect 8539 7497 8573 7531
rect 8953 7497 8987 7531
rect 13461 7497 13495 7531
rect 15025 7497 15059 7531
rect 16221 7497 16255 7531
rect 17095 7497 17129 7531
rect 19993 7497 20027 7531
rect 22845 7497 22879 7531
rect 25053 7497 25087 7531
rect 25697 7497 25731 7531
rect 2237 7429 2271 7463
rect 3709 7429 3743 7463
rect 8125 7429 8159 7463
rect 10149 7429 10183 7463
rect 11345 7429 11379 7463
rect 13001 7429 13035 7463
rect 14289 7429 14323 7463
rect 2697 7361 2731 7395
rect 4997 7361 5031 7395
rect 10885 7361 10919 7395
rect 17877 7361 17911 7395
rect 18705 7361 18739 7395
rect 19625 7361 19659 7395
rect 20729 7361 20763 7395
rect 1660 7293 1694 7327
rect 2789 7293 2823 7327
rect 6653 7293 6687 7327
rect 7021 7293 7055 7327
rect 7297 7293 7331 7327
rect 8468 7293 8502 7327
rect 11161 7293 11195 7327
rect 11989 7293 12023 7327
rect 12516 7293 12550 7327
rect 15209 7293 15243 7327
rect 15761 7293 15795 7327
rect 16992 7293 17026 7327
rect 17417 7293 17451 7327
rect 20453 7293 20487 7327
rect 20637 7293 20671 7327
rect 21741 7293 21775 7327
rect 22293 7293 22327 7327
rect 23673 7293 23707 7327
rect 24225 7293 24259 7327
rect 24685 7293 24719 7327
rect 25272 7293 25306 7327
rect 26065 7293 26099 7327
rect 3110 7225 3144 7259
rect 9597 7225 9631 7259
rect 9689 7225 9723 7259
rect 13737 7225 13771 7259
rect 13829 7225 13863 7259
rect 14749 7225 14783 7259
rect 16681 7225 16715 7259
rect 18797 7225 18831 7259
rect 19349 7225 19383 7259
rect 4905 7157 4939 7191
rect 5365 7157 5399 7191
rect 6929 7157 6963 7191
rect 9413 7157 9447 7191
rect 10517 7157 10551 7191
rect 11621 7157 11655 7191
rect 12725 7157 12759 7191
rect 15485 7157 15519 7191
rect 18429 7157 18463 7191
rect 21189 7157 21223 7191
rect 21557 7157 21591 7191
rect 21833 7157 21867 7191
rect 23397 7157 23431 7191
rect 23765 7157 23799 7191
rect 25375 7157 25409 7191
rect 1961 6953 1995 6987
rect 3433 6953 3467 6987
rect 5549 6953 5583 6987
rect 7021 6953 7055 6987
rect 9781 6953 9815 6987
rect 13737 6953 13771 6987
rect 15439 6953 15473 6987
rect 17417 6953 17451 6987
rect 18245 6953 18279 6987
rect 18797 6953 18831 6987
rect 19073 6953 19107 6987
rect 19763 6953 19797 6987
rect 20269 6953 20303 6987
rect 22753 6953 22787 6987
rect 22937 6953 22971 6987
rect 24317 6953 24351 6987
rect 24961 6953 24995 6987
rect 3157 6885 3191 6919
rect 4905 6885 4939 6919
rect 6009 6885 6043 6919
rect 7665 6885 7699 6919
rect 9505 6885 9539 6919
rect 11391 6885 11425 6919
rect 12725 6885 12759 6919
rect 13277 6885 13311 6919
rect 21878 6885 21912 6919
rect 1476 6817 1510 6851
rect 2421 6817 2455 6851
rect 3801 6817 3835 6851
rect 4169 6817 4203 6851
rect 4721 6817 4755 6851
rect 5733 6817 5767 6851
rect 6653 6817 6687 6851
rect 9873 6817 9907 6851
rect 10149 6817 10183 6851
rect 10701 6817 10735 6851
rect 11288 6817 11322 6851
rect 14264 6817 14298 6851
rect 15209 6817 15243 6851
rect 16313 6817 16347 6851
rect 16773 6817 16807 6851
rect 19660 6817 19694 6851
rect 2789 6749 2823 6783
rect 7573 6749 7607 6783
rect 8861 6749 8895 6783
rect 12633 6749 12667 6783
rect 17049 6749 17083 6783
rect 17877 6749 17911 6783
rect 21557 6749 21591 6783
rect 1547 6681 1581 6715
rect 8125 6681 8159 6715
rect 8585 6681 8619 6715
rect 22477 6681 22511 6715
rect 23489 6885 23523 6919
rect 24041 6885 24075 6919
rect 25145 6817 25179 6851
rect 25421 6817 25455 6851
rect 23397 6749 23431 6783
rect 24685 6749 24719 6783
rect 23121 6681 23155 6715
rect 2329 6613 2363 6647
rect 2559 6613 2593 6647
rect 2697 6613 2731 6647
rect 5181 6613 5215 6647
rect 7297 6613 7331 6647
rect 11713 6613 11747 6647
rect 14105 6613 14139 6647
rect 14335 6613 14369 6647
rect 15761 6613 15795 6647
rect 16221 6613 16255 6647
rect 17785 6613 17819 6647
rect 21465 6613 21499 6647
rect 22937 6613 22971 6647
rect 3065 6409 3099 6443
rect 4261 6409 4295 6443
rect 6193 6409 6227 6443
rect 7297 6409 7331 6443
rect 8493 6409 8527 6443
rect 8953 6409 8987 6443
rect 11529 6409 11563 6443
rect 12265 6409 12299 6443
rect 16313 6409 16347 6443
rect 17003 6409 17037 6443
rect 17233 6409 17267 6443
rect 17417 6409 17451 6443
rect 22937 6409 22971 6443
rect 23121 6409 23155 6443
rect 23397 6409 23431 6443
rect 4721 6341 4755 6375
rect 5917 6341 5951 6375
rect 9413 6341 9447 6375
rect 14381 6341 14415 6375
rect 3801 6273 3835 6307
rect 4905 6273 4939 6307
rect 7573 6273 7607 6307
rect 10333 6273 10367 6307
rect 11253 6273 11287 6307
rect 13829 6273 13863 6307
rect 15209 6273 15243 6307
rect 15393 6273 15427 6307
rect 24961 6341 24995 6375
rect 25421 6341 25455 6375
rect 18153 6273 18187 6307
rect 20453 6273 20487 6307
rect 22937 6273 22971 6307
rect 25789 6273 25823 6307
rect 2053 6205 2087 6239
rect 3525 6205 3559 6239
rect 3709 6205 3743 6239
rect 5549 6205 5583 6239
rect 9505 6205 9539 6239
rect 9965 6205 9999 6239
rect 10517 6205 10551 6239
rect 10977 6205 11011 6239
rect 12792 6205 12826 6239
rect 13185 6205 13219 6239
rect 14749 6205 14783 6239
rect 16932 6205 16966 6239
rect 17233 6205 17267 6239
rect 19625 6205 19659 6239
rect 19993 6205 20027 6239
rect 20361 6205 20395 6239
rect 21557 6205 21591 6239
rect 23673 6205 23707 6239
rect 24133 6205 24167 6239
rect 25237 6205 25271 6239
rect 2421 6137 2455 6171
rect 4997 6137 5031 6171
rect 6653 6137 6687 6171
rect 7665 6137 7699 6171
rect 8217 6137 8251 6171
rect 13921 6137 13955 6171
rect 15485 6137 15519 6171
rect 16037 6137 16071 6171
rect 16773 6137 16807 6171
rect 18474 6137 18508 6171
rect 21878 6137 21912 6171
rect 2789 6069 2823 6103
rect 9689 6069 9723 6103
rect 12863 6069 12897 6103
rect 13645 6069 13679 6103
rect 17877 6069 17911 6103
rect 19073 6069 19107 6103
rect 21005 6069 21039 6103
rect 21373 6069 21407 6103
rect 22477 6069 22511 6103
rect 23765 6069 23799 6103
rect 3065 5865 3099 5899
rect 3249 5865 3283 5899
rect 1547 5797 1581 5831
rect 1444 5729 1478 5763
rect 2421 5729 2455 5763
rect 2789 5661 2823 5695
rect 2329 5593 2363 5627
rect 4721 5865 4755 5899
rect 5273 5865 5307 5899
rect 6929 5865 6963 5899
rect 7389 5865 7423 5899
rect 7941 5865 7975 5899
rect 8217 5865 8251 5899
rect 13461 5865 13495 5899
rect 15669 5865 15703 5899
rect 16221 5865 16255 5899
rect 18429 5865 18463 5899
rect 21005 5865 21039 5899
rect 24225 5865 24259 5899
rect 6285 5797 6319 5831
rect 11069 5797 11103 5831
rect 13737 5797 13771 5831
rect 13829 5797 13863 5831
rect 14381 5797 14415 5831
rect 17233 5797 17267 5831
rect 19073 5797 19107 5831
rect 19993 5797 20027 5831
rect 20361 5797 20395 5831
rect 22293 5797 22327 5831
rect 22753 5797 22787 5831
rect 23305 5797 23339 5831
rect 10149 5729 10183 5763
rect 10333 5729 10367 5763
rect 12357 5729 12391 5763
rect 12541 5729 12575 5763
rect 13093 5729 13127 5763
rect 20913 5729 20947 5763
rect 21373 5729 21407 5763
rect 24133 5729 24167 5763
rect 24593 5729 24627 5763
rect 4353 5661 4387 5695
rect 5549 5661 5583 5695
rect 7021 5661 7055 5695
rect 10701 5661 10735 5695
rect 12817 5661 12851 5695
rect 15301 5661 15335 5695
rect 17141 5661 17175 5695
rect 18981 5661 19015 5695
rect 19257 5661 19291 5695
rect 22661 5661 22695 5695
rect 10609 5593 10643 5627
rect 14749 5593 14783 5627
rect 17693 5593 17727 5627
rect 22017 5593 22051 5627
rect 1961 5525 1995 5559
rect 2559 5525 2593 5559
rect 2697 5525 2731 5559
rect 3249 5525 3283 5559
rect 3433 5525 3467 5559
rect 3893 5525 3927 5559
rect 5917 5525 5951 5559
rect 10498 5525 10532 5559
rect 11345 5525 11379 5559
rect 18061 5525 18095 5559
rect 23765 5525 23799 5559
rect 25145 5525 25179 5559
rect 6285 5321 6319 5355
rect 9689 5321 9723 5355
rect 9965 5321 9999 5355
rect 10333 5321 10367 5355
rect 10655 5321 10689 5355
rect 11161 5321 11195 5355
rect 12173 5321 12207 5355
rect 12633 5321 12667 5355
rect 13093 5321 13127 5355
rect 14841 5321 14875 5355
rect 17233 5321 17267 5355
rect 19257 5321 19291 5355
rect 19625 5321 19659 5355
rect 21097 5321 21131 5355
rect 22477 5321 22511 5355
rect 22753 5321 22787 5355
rect 23397 5321 23431 5355
rect 24685 5321 24719 5355
rect 1961 5253 1995 5287
rect 3065 5253 3099 5287
rect 4445 5253 4479 5287
rect 10793 5253 10827 5287
rect 20269 5253 20303 5287
rect 2053 5185 2087 5219
rect 3985 5185 4019 5219
rect 4905 5185 4939 5219
rect 6837 5185 6871 5219
rect 10885 5185 10919 5219
rect 13921 5185 13955 5219
rect 15669 5185 15703 5219
rect 16865 5185 16899 5219
rect 18337 5185 18371 5219
rect 20637 5185 20671 5219
rect 1832 5117 1866 5151
rect 3249 5117 3283 5151
rect 3801 5117 3835 5151
rect 8401 5117 8435 5151
rect 8585 5117 8619 5151
rect 9045 5117 9079 5151
rect 10517 5117 10551 5151
rect 12909 5117 12943 5151
rect 20085 5117 20119 5151
rect 21189 5117 21223 5151
rect 23673 5117 23707 5151
rect 24133 5117 24167 5151
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 1685 5049 1719 5083
rect 4997 5049 5031 5083
rect 5549 5049 5583 5083
rect 11529 5049 11563 5083
rect 14283 5049 14317 5083
rect 15990 5049 16024 5083
rect 18429 5049 18463 5083
rect 18981 5049 19015 5083
rect 21510 5049 21544 5083
rect 2329 4981 2363 5015
rect 2697 4981 2731 5015
rect 5825 4981 5859 5015
rect 6653 4981 6687 5015
rect 7205 4981 7239 5015
rect 7757 4981 7791 5015
rect 8033 4981 8067 5015
rect 8677 4981 8711 5015
rect 13461 4981 13495 5015
rect 13829 4981 13863 5015
rect 15301 4981 15335 5015
rect 16589 4981 16623 5015
rect 17785 4981 17819 5015
rect 22109 4981 22143 5015
rect 23765 4981 23799 5015
rect 25421 4981 25455 5015
rect 1547 4777 1581 4811
rect 2329 4777 2363 4811
rect 3525 4777 3559 4811
rect 3801 4777 3835 4811
rect 4261 4777 4295 4811
rect 4721 4777 4755 4811
rect 6469 4777 6503 4811
rect 6929 4777 6963 4811
rect 8217 4777 8251 4811
rect 8677 4777 8711 4811
rect 10333 4777 10367 4811
rect 10701 4777 10735 4811
rect 11345 4777 11379 4811
rect 14473 4777 14507 4811
rect 15025 4777 15059 4811
rect 17049 4777 17083 4811
rect 18153 4777 18187 4811
rect 19257 4777 19291 4811
rect 20637 4777 20671 4811
rect 22569 4777 22603 4811
rect 24501 4777 24535 4811
rect 1869 4709 1903 4743
rect 3157 4709 3191 4743
rect 5089 4709 5123 4743
rect 5641 4709 5675 4743
rect 7297 4709 7331 4743
rect 7389 4709 7423 4743
rect 9045 4709 9079 4743
rect 9689 4709 9723 4743
rect 13645 4709 13679 4743
rect 14197 4709 14231 4743
rect 16221 4709 16255 4743
rect 16773 4709 16807 4743
rect 18429 4709 18463 4743
rect 21418 4709 21452 4743
rect 23029 4709 23063 4743
rect 23581 4709 23615 4743
rect 24133 4709 24167 4743
rect 1476 4641 1510 4675
rect 2421 4641 2455 4675
rect 11529 4641 11563 4675
rect 11805 4641 11839 4675
rect 19876 4641 19910 4675
rect 24409 4641 24443 4675
rect 24869 4641 24903 4675
rect 2789 4573 2823 4607
rect 4997 4573 5031 4607
rect 5917 4573 5951 4607
rect 7573 4573 7607 4607
rect 10057 4573 10091 4607
rect 13553 4573 13587 4607
rect 16129 4573 16163 4607
rect 18337 4573 18371 4607
rect 18981 4573 19015 4607
rect 21097 4573 21131 4607
rect 22937 4573 22971 4607
rect 2697 4505 2731 4539
rect 9965 4505 9999 4539
rect 19947 4505 19981 4539
rect 2559 4437 2593 4471
rect 9413 4437 9447 4471
rect 9854 4437 9888 4471
rect 11069 4437 11103 4471
rect 12265 4437 12299 4471
rect 13277 4437 13311 4471
rect 15669 4437 15703 4471
rect 17509 4437 17543 4471
rect 22017 4437 22051 4471
rect 7849 4233 7883 4267
rect 9597 4233 9631 4267
rect 10057 4233 10091 4267
rect 11253 4233 11287 4267
rect 12173 4233 12207 4267
rect 12633 4233 12667 4267
rect 16129 4233 16163 4267
rect 17509 4233 17543 4267
rect 18981 4233 19015 4267
rect 19349 4233 19383 4267
rect 21833 4233 21867 4267
rect 24685 4233 24719 4267
rect 2973 4165 3007 4199
rect 5641 4165 5675 4199
rect 9919 4165 9953 4199
rect 11529 4165 11563 4199
rect 14565 4165 14599 4199
rect 15761 4165 15795 4199
rect 17049 4165 17083 4199
rect 19717 4165 19751 4199
rect 22569 4165 22603 4199
rect 25421 4165 25455 4199
rect 1777 4097 1811 4131
rect 5089 4097 5123 4131
rect 6929 4097 6963 4131
rect 10149 4097 10183 4131
rect 14013 4097 14047 4131
rect 16497 4097 16531 4131
rect 20545 4097 20579 4131
rect 25789 4097 25823 4131
rect 1869 4029 1903 4063
rect 2237 4029 2271 4063
rect 2421 4029 2455 4063
rect 3709 4029 3743 4063
rect 3985 4029 4019 4063
rect 8585 4029 8619 4063
rect 9229 4029 9263 4063
rect 10517 4029 10551 4063
rect 11345 4029 11379 4063
rect 11805 4029 11839 4063
rect 12449 4029 12483 4063
rect 18061 4029 18095 4063
rect 23489 4029 23523 4063
rect 23673 4029 23707 4063
rect 24225 4029 24259 4063
rect 25237 4029 25271 4063
rect 3341 3961 3375 3995
rect 4169 3961 4203 3995
rect 4905 3961 4939 3995
rect 5181 3961 5215 3995
rect 6653 3961 6687 3995
rect 7021 3961 7055 3995
rect 7573 3961 7607 3995
rect 8401 3961 8435 3995
rect 8953 3961 8987 3995
rect 9781 3961 9815 3995
rect 14105 3961 14139 3995
rect 14933 3961 14967 3995
rect 16589 3961 16623 3995
rect 18382 3961 18416 3995
rect 19901 3961 19935 3995
rect 19993 3961 20027 3995
rect 22017 3961 22051 3995
rect 22109 3961 22143 3995
rect 4537 3893 4571 3927
rect 6009 3893 6043 3927
rect 8309 3893 8343 3927
rect 10793 3893 10827 3927
rect 13001 3893 13035 3927
rect 13553 3893 13587 3927
rect 15393 3893 15427 3927
rect 17877 3893 17911 3927
rect 21097 3893 21131 3927
rect 23029 3893 23063 3927
rect 23765 3893 23799 3927
rect 25145 3893 25179 3927
rect 2697 3689 2731 3723
rect 3433 3689 3467 3723
rect 3617 3689 3651 3723
rect 3801 3689 3835 3723
rect 5365 3689 5399 3723
rect 5641 3689 5675 3723
rect 9045 3689 9079 3723
rect 9229 3689 9263 3723
rect 9873 3689 9907 3723
rect 10241 3689 10275 3723
rect 10517 3689 10551 3723
rect 11621 3689 11655 3723
rect 16865 3689 16899 3723
rect 19349 3689 19383 3723
rect 21189 3689 21223 3723
rect 22661 3689 22695 3723
rect 24869 3689 24903 3723
rect 1547 3621 1581 3655
rect 1460 3553 1494 3587
rect 3065 3553 3099 3587
rect 1961 3485 1995 3519
rect 4261 3621 4295 3655
rect 4766 3621 4800 3655
rect 7389 3621 7423 3655
rect 7941 3621 7975 3655
rect 4445 3553 4479 3587
rect 6009 3553 6043 3587
rect 6193 3553 6227 3587
rect 9229 3553 9263 3587
rect 12173 3621 12207 3655
rect 13001 3621 13035 3655
rect 13829 3621 13863 3655
rect 14381 3621 14415 3655
rect 15485 3621 15519 3655
rect 16037 3621 16071 3655
rect 16497 3621 16531 3655
rect 18429 3621 18463 3655
rect 18981 3621 19015 3655
rect 20269 3621 20303 3655
rect 21833 3621 21867 3655
rect 10517 3553 10551 3587
rect 10609 3553 10643 3587
rect 12357 3553 12391 3587
rect 17141 3553 17175 3587
rect 19809 3553 19843 3587
rect 21465 3553 21499 3587
rect 22385 3553 22419 3587
rect 23305 3553 23339 3587
rect 23673 3553 23707 3587
rect 25053 3553 25087 3587
rect 25329 3553 25363 3587
rect 7297 3485 7331 3519
rect 8217 3485 8251 3519
rect 10977 3485 11011 3519
rect 13737 3485 13771 3519
rect 14657 3485 14691 3519
rect 15117 3485 15151 3519
rect 15393 3485 15427 3519
rect 17785 3485 17819 3519
rect 18337 3485 18371 3519
rect 21741 3485 21775 3519
rect 23121 3485 23155 3519
rect 23765 3485 23799 3519
rect 3617 3417 3651 3451
rect 6377 3417 6411 3451
rect 8677 3417 8711 3451
rect 11989 3417 12023 3451
rect 17325 3417 17359 3451
rect 19993 3417 20027 3451
rect 24593 3417 24627 3451
rect 2237 3349 2271 3383
rect 7021 3349 7055 3383
rect 9505 3349 9539 3383
rect 10747 3349 10781 3383
rect 10885 3349 10919 3383
rect 11253 3349 11287 3383
rect 12449 3349 12483 3383
rect 13369 3349 13403 3383
rect 18153 3349 18187 3383
rect 24225 3349 24259 3383
rect 2881 3145 2915 3179
rect 6653 3145 6687 3179
rect 7849 3145 7883 3179
rect 8125 3145 8159 3179
rect 9689 3145 9723 3179
rect 10057 3145 10091 3179
rect 12265 3145 12299 3179
rect 13737 3145 13771 3179
rect 14013 3145 14047 3179
rect 15485 3145 15519 3179
rect 15761 3145 15795 3179
rect 16129 3145 16163 3179
rect 17325 3145 17359 3179
rect 19809 3145 19843 3179
rect 22385 3145 22419 3179
rect 22845 3145 22879 3179
rect 23121 3145 23155 3179
rect 24685 3145 24719 3179
rect 25053 3145 25087 3179
rect 4537 3077 4571 3111
rect 5549 3077 5583 3111
rect 8585 3077 8619 3111
rect 10379 3077 10413 3111
rect 10517 3077 10551 3111
rect 23811 3077 23845 3111
rect 23949 3077 23983 3111
rect 25421 3077 25455 3111
rect 2513 3009 2547 3043
rect 4997 3009 5031 3043
rect 10609 3009 10643 3043
rect 16405 3009 16439 3043
rect 17049 3009 17083 3043
rect 18797 3009 18831 3043
rect 19073 3009 19107 3043
rect 20361 3009 20395 3043
rect 20821 3009 20855 3043
rect 24041 3009 24075 3043
rect 24133 3009 24167 3043
rect 2237 2941 2271 2975
rect 3433 2941 3467 2975
rect 3801 2941 3835 2975
rect 6929 2941 6963 2975
rect 8953 2941 8987 2975
rect 9137 2941 9171 2975
rect 10241 2941 10275 2975
rect 11253 2941 11287 2975
rect 12817 2941 12851 2975
rect 14565 2941 14599 2975
rect 22636 2941 22670 2975
rect 23397 2941 23431 2975
rect 23673 2941 23707 2975
rect 25237 2941 25271 2975
rect 4077 2873 4111 2907
rect 5089 2873 5123 2907
rect 10977 2873 11011 2907
rect 13138 2873 13172 2907
rect 14381 2873 14415 2907
rect 14886 2873 14920 2907
rect 16497 2873 16531 2907
rect 18889 2873 18923 2907
rect 20729 2873 20763 2907
rect 21142 2873 21176 2907
rect 26157 2873 26191 2907
rect 1685 2805 1719 2839
rect 3249 2805 3283 2839
rect 6193 2805 6227 2839
rect 7297 2805 7331 2839
rect 8769 2805 8803 2839
rect 11713 2805 11747 2839
rect 12633 2805 12667 2839
rect 17785 2805 17819 2839
rect 18337 2805 18371 2839
rect 21741 2805 21775 2839
rect 22017 2805 22051 2839
rect 25789 2805 25823 2839
rect 3433 2601 3467 2635
rect 3801 2601 3835 2635
rect 4905 2601 4939 2635
rect 6009 2601 6043 2635
rect 6653 2601 6687 2635
rect 7941 2601 7975 2635
rect 8309 2601 8343 2635
rect 8493 2601 8527 2635
rect 9597 2601 9631 2635
rect 10885 2601 10919 2635
rect 11989 2601 12023 2635
rect 13645 2601 13679 2635
rect 16313 2601 16347 2635
rect 17417 2601 17451 2635
rect 19257 2601 19291 2635
rect 20223 2601 20257 2635
rect 22293 2601 22327 2635
rect 23857 2601 23891 2635
rect 24133 2601 24167 2635
rect 24869 2601 24903 2635
rect 25513 2601 25547 2635
rect 2329 2533 2363 2567
rect 5410 2533 5444 2567
rect 7021 2533 7055 2567
rect 7113 2533 7147 2567
rect 7665 2533 7699 2567
rect 1444 2465 1478 2499
rect 1869 2465 1903 2499
rect 2697 2465 2731 2499
rect 2973 2465 3007 2499
rect 4144 2465 4178 2499
rect 5089 2465 5123 2499
rect 6285 2465 6319 2499
rect 3157 2397 3191 2431
rect 4215 2329 4249 2363
rect 8677 2465 8711 2499
rect 9137 2465 9171 2499
rect 9781 2465 9815 2499
rect 11713 2533 11747 2567
rect 13046 2533 13080 2567
rect 16818 2533 16852 2567
rect 18061 2533 18095 2567
rect 18658 2533 18692 2567
rect 21005 2533 21039 2567
rect 21465 2533 21499 2567
rect 22017 2533 22051 2567
rect 25053 2533 25087 2567
rect 11253 2465 11287 2499
rect 11437 2465 11471 2499
rect 15485 2465 15519 2499
rect 15945 2465 15979 2499
rect 17785 2465 17819 2499
rect 18337 2465 18371 2499
rect 20120 2465 20154 2499
rect 20545 2465 20579 2499
rect 22845 2465 22879 2499
rect 23489 2465 23523 2499
rect 24225 2465 24259 2499
rect 24593 2465 24627 2499
rect 24869 2465 24903 2499
rect 25672 2465 25706 2499
rect 12725 2397 12759 2431
rect 13921 2397 13955 2431
rect 15301 2397 15335 2431
rect 16497 2397 16531 2431
rect 21373 2397 21407 2431
rect 12357 2329 12391 2363
rect 15669 2329 15703 2363
rect 23029 2329 23063 2363
rect 25743 2329 25777 2363
rect 1547 2261 1581 2295
rect 4629 2261 4663 2295
rect 8493 2261 8527 2295
rect 8861 2261 8895 2295
rect 9965 2261 9999 2295
rect 10333 2261 10367 2295
rect 10701 2261 10735 2295
rect 10885 2261 10919 2295
rect 14657 2261 14691 2295
rect 22661 2261 22695 2295
rect 26157 2261 26191 2295
<< metal1 >>
rect 5534 27480 5540 27532
rect 5592 27520 5598 27532
rect 6178 27520 6184 27532
rect 5592 27492 6184 27520
rect 5592 27480 5598 27492
rect 6178 27480 6184 27492
rect 6236 27480 6242 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 18322 24828 18328 24880
rect 18380 24868 18386 24880
rect 27614 24868 27620 24880
rect 18380 24840 27620 24868
rect 18380 24828 18386 24840
rect 27614 24828 27620 24840
rect 27672 24828 27678 24880
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 18233 24395 18291 24401
rect 18233 24361 18245 24395
rect 18279 24392 18291 24395
rect 20162 24392 20168 24404
rect 18279 24364 20168 24392
rect 18279 24361 18291 24364
rect 18233 24355 18291 24361
rect 20162 24352 20168 24364
rect 20220 24352 20226 24404
rect 10686 24265 10692 24268
rect 10664 24259 10692 24265
rect 10664 24256 10676 24259
rect 10599 24228 10676 24256
rect 10664 24225 10676 24228
rect 10744 24256 10750 24268
rect 11514 24256 11520 24268
rect 10744 24228 11520 24256
rect 10664 24219 10692 24225
rect 10686 24216 10692 24219
rect 10744 24216 10750 24228
rect 11514 24216 11520 24228
rect 11572 24216 11578 24268
rect 11609 24259 11667 24265
rect 11609 24225 11621 24259
rect 11655 24256 11667 24259
rect 11698 24256 11704 24268
rect 11655 24228 11704 24256
rect 11655 24225 11667 24228
rect 11609 24219 11667 24225
rect 11698 24216 11704 24228
rect 11756 24216 11762 24268
rect 16942 24256 16948 24268
rect 16903 24228 16948 24256
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 18046 24256 18052 24268
rect 18007 24228 18052 24256
rect 18046 24216 18052 24228
rect 18104 24216 18110 24268
rect 17129 24123 17187 24129
rect 17129 24089 17141 24123
rect 17175 24120 17187 24123
rect 18782 24120 18788 24132
rect 17175 24092 18788 24120
rect 17175 24089 17187 24092
rect 17129 24083 17187 24089
rect 18782 24080 18788 24092
rect 18840 24080 18846 24132
rect 9766 24012 9772 24064
rect 9824 24052 9830 24064
rect 10735 24055 10793 24061
rect 10735 24052 10747 24055
rect 9824 24024 10747 24052
rect 9824 24012 9830 24024
rect 10735 24021 10747 24024
rect 10781 24021 10793 24055
rect 10735 24015 10793 24021
rect 11330 24012 11336 24064
rect 11388 24052 11394 24064
rect 11747 24055 11805 24061
rect 11747 24052 11759 24055
rect 11388 24024 11759 24052
rect 11388 24012 11394 24024
rect 11747 24021 11759 24024
rect 11793 24021 11805 24055
rect 11747 24015 11805 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 10686 23848 10692 23860
rect 10647 23820 10692 23848
rect 10686 23808 10692 23820
rect 10744 23808 10750 23860
rect 14553 23851 14611 23857
rect 14553 23817 14565 23851
rect 14599 23848 14611 23851
rect 16022 23848 16028 23860
rect 14599 23820 16028 23848
rect 14599 23817 14611 23820
rect 14553 23811 14611 23817
rect 16022 23808 16028 23820
rect 16080 23808 16086 23860
rect 16209 23851 16267 23857
rect 16209 23817 16221 23851
rect 16255 23848 16267 23851
rect 17402 23848 17408 23860
rect 16255 23820 17408 23848
rect 16255 23817 16267 23820
rect 16209 23811 16267 23817
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 18046 23808 18052 23860
rect 18104 23848 18110 23860
rect 18506 23848 18512 23860
rect 18104 23820 18512 23848
rect 18104 23808 18110 23820
rect 18506 23808 18512 23820
rect 18564 23848 18570 23860
rect 18601 23851 18659 23857
rect 18601 23848 18613 23851
rect 18564 23820 18613 23848
rect 18564 23808 18570 23820
rect 18601 23817 18613 23820
rect 18647 23817 18659 23851
rect 18601 23811 18659 23817
rect 20349 23851 20407 23857
rect 20349 23817 20361 23851
rect 20395 23848 20407 23851
rect 21634 23848 21640 23860
rect 20395 23820 21640 23848
rect 20395 23817 20407 23820
rect 20349 23811 20407 23817
rect 21634 23808 21640 23820
rect 21692 23808 21698 23860
rect 22557 23851 22615 23857
rect 22557 23817 22569 23851
rect 22603 23848 22615 23851
rect 24210 23848 24216 23860
rect 22603 23820 24216 23848
rect 22603 23817 22615 23820
rect 22557 23811 22615 23817
rect 24210 23808 24216 23820
rect 24268 23808 24274 23860
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 21453 23783 21511 23789
rect 21453 23749 21465 23783
rect 21499 23780 21511 23783
rect 22646 23780 22652 23792
rect 21499 23752 22652 23780
rect 21499 23749 21511 23752
rect 21453 23743 21511 23749
rect 22646 23740 22652 23752
rect 22704 23740 22710 23792
rect 24210 23672 24216 23724
rect 24268 23712 24274 23724
rect 27154 23712 27160 23724
rect 24268 23684 27160 23712
rect 24268 23672 24274 23684
rect 27154 23672 27160 23684
rect 27212 23672 27218 23724
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 1946 23644 1952 23656
rect 1443 23616 1952 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 1946 23604 1952 23616
rect 2004 23604 2010 23656
rect 7190 23604 7196 23656
rect 7248 23644 7254 23656
rect 8941 23647 8999 23653
rect 8941 23644 8953 23647
rect 7248 23616 8953 23644
rect 7248 23604 7254 23616
rect 8941 23613 8953 23616
rect 8987 23644 8999 23647
rect 9401 23647 9459 23653
rect 9401 23644 9413 23647
rect 8987 23616 9413 23644
rect 8987 23613 8999 23616
rect 8941 23607 8999 23613
rect 9401 23613 9413 23616
rect 9447 23613 9459 23647
rect 9401 23607 9459 23613
rect 11124 23647 11182 23653
rect 11124 23613 11136 23647
rect 11170 23644 11182 23647
rect 11238 23644 11244 23656
rect 11170 23616 11244 23644
rect 11170 23613 11182 23616
rect 11124 23607 11182 23613
rect 11238 23604 11244 23616
rect 11296 23604 11302 23656
rect 11514 23604 11520 23656
rect 11572 23644 11578 23656
rect 12472 23647 12530 23653
rect 12472 23644 12484 23647
rect 11572 23616 12484 23644
rect 11572 23604 11578 23616
rect 12472 23613 12484 23616
rect 12518 23644 12530 23647
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12518 23616 12909 23644
rect 12518 23613 12530 23616
rect 12472 23607 12530 23613
rect 12897 23613 12909 23616
rect 12943 23613 12955 23647
rect 14366 23644 14372 23656
rect 14279 23616 14372 23644
rect 12897 23607 12955 23613
rect 14366 23604 14372 23616
rect 14424 23644 14430 23656
rect 14921 23647 14979 23653
rect 14921 23644 14933 23647
rect 14424 23616 14933 23644
rect 14424 23604 14430 23616
rect 14921 23613 14933 23616
rect 14967 23613 14979 23647
rect 16025 23647 16083 23653
rect 16025 23644 16037 23647
rect 14921 23607 14979 23613
rect 15212 23616 16037 23644
rect 12986 23536 12992 23588
rect 13044 23576 13050 23588
rect 15212 23576 15240 23616
rect 16025 23613 16037 23616
rect 16071 23644 16083 23647
rect 16577 23647 16635 23653
rect 16577 23644 16589 23647
rect 16071 23616 16589 23644
rect 16071 23613 16083 23616
rect 16025 23607 16083 23613
rect 16577 23613 16589 23616
rect 16623 23613 16635 23647
rect 16577 23607 16635 23613
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17911 23616 18061 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18049 23613 18061 23616
rect 18095 23644 18107 23647
rect 18138 23644 18144 23656
rect 18095 23616 18144 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 18138 23604 18144 23616
rect 18196 23604 18202 23656
rect 20165 23647 20223 23653
rect 20165 23613 20177 23647
rect 20211 23644 20223 23647
rect 21266 23644 21272 23656
rect 20211 23616 20852 23644
rect 21179 23616 21272 23644
rect 20211 23613 20223 23616
rect 20165 23607 20223 23613
rect 13044 23548 15240 23576
rect 13044 23536 13050 23548
rect 15286 23536 15292 23588
rect 15344 23576 15350 23588
rect 16942 23576 16948 23588
rect 15344 23548 16948 23576
rect 15344 23536 15350 23548
rect 16942 23536 16948 23548
rect 17000 23536 17006 23588
rect 5258 23468 5264 23520
rect 5316 23508 5322 23520
rect 9125 23511 9183 23517
rect 9125 23508 9137 23511
rect 5316 23480 9137 23508
rect 5316 23468 5322 23480
rect 9125 23477 9137 23480
rect 9171 23477 9183 23511
rect 9950 23508 9956 23520
rect 9911 23480 9956 23508
rect 9125 23471 9183 23477
rect 9950 23468 9956 23480
rect 10008 23468 10014 23520
rect 10686 23468 10692 23520
rect 10744 23508 10750 23520
rect 11195 23511 11253 23517
rect 11195 23508 11207 23511
rect 10744 23480 11207 23508
rect 10744 23468 10750 23480
rect 11195 23477 11207 23480
rect 11241 23477 11253 23511
rect 11698 23508 11704 23520
rect 11611 23480 11704 23508
rect 11195 23471 11253 23477
rect 11698 23468 11704 23480
rect 11756 23508 11762 23520
rect 12250 23508 12256 23520
rect 11756 23480 12256 23508
rect 11756 23468 11762 23480
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 12575 23511 12633 23517
rect 12575 23477 12587 23511
rect 12621 23508 12633 23511
rect 12710 23508 12716 23520
rect 12621 23480 12716 23508
rect 12621 23477 12633 23480
rect 12575 23471 12633 23477
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 18230 23508 18236 23520
rect 18191 23480 18236 23508
rect 18230 23468 18236 23480
rect 18288 23468 18294 23520
rect 20824 23517 20852 23616
rect 21266 23604 21272 23616
rect 21324 23644 21330 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21324 23616 21833 23644
rect 21324 23604 21330 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 21910 23604 21916 23656
rect 21968 23644 21974 23656
rect 22373 23647 22431 23653
rect 22373 23644 22385 23647
rect 21968 23616 22385 23644
rect 21968 23604 21974 23616
rect 22373 23613 22385 23616
rect 22419 23644 22431 23647
rect 22925 23647 22983 23653
rect 22925 23644 22937 23647
rect 22419 23616 22937 23644
rect 22419 23613 22431 23616
rect 22373 23607 22431 23613
rect 22925 23613 22937 23616
rect 22971 23613 22983 23647
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 22925 23607 22983 23613
rect 23446 23616 24593 23644
rect 23446 23576 23474 23616
rect 24581 23613 24593 23616
rect 24627 23644 24639 23647
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 24627 23616 25145 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 22388 23548 23474 23576
rect 22388 23520 22416 23548
rect 20809 23511 20867 23517
rect 20809 23477 20821 23511
rect 20855 23508 20867 23511
rect 21082 23508 21088 23520
rect 20855 23480 21088 23508
rect 20855 23477 20867 23480
rect 20809 23471 20867 23477
rect 21082 23468 21088 23480
rect 21140 23468 21146 23520
rect 22370 23468 22376 23520
rect 22428 23468 22434 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1118 23264 1124 23316
rect 1176 23304 1182 23316
rect 1581 23307 1639 23313
rect 1581 23304 1593 23307
rect 1176 23276 1593 23304
rect 1176 23264 1182 23276
rect 1581 23273 1593 23276
rect 1627 23273 1639 23307
rect 11146 23304 11152 23316
rect 11059 23276 11152 23304
rect 1581 23267 1639 23273
rect 11146 23264 11152 23276
rect 11204 23304 11210 23316
rect 13170 23304 13176 23316
rect 11204 23276 13176 23304
rect 11204 23264 11210 23276
rect 13170 23264 13176 23276
rect 13228 23264 13234 23316
rect 13679 23307 13737 23313
rect 13679 23273 13691 23307
rect 13725 23304 13737 23307
rect 14366 23304 14372 23316
rect 13725 23276 14372 23304
rect 13725 23273 13737 23276
rect 13679 23267 13737 23273
rect 14366 23264 14372 23276
rect 14424 23264 14430 23316
rect 18233 23307 18291 23313
rect 18233 23273 18245 23307
rect 18279 23304 18291 23307
rect 18322 23304 18328 23316
rect 18279 23276 18328 23304
rect 18279 23273 18291 23276
rect 18233 23267 18291 23273
rect 18322 23264 18328 23276
rect 18380 23264 18386 23316
rect 24765 23307 24823 23313
rect 24765 23273 24777 23307
rect 24811 23304 24823 23307
rect 24854 23304 24860 23316
rect 24811 23276 24860 23304
rect 24811 23273 24823 23276
rect 24765 23267 24823 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 1946 23196 1952 23248
rect 2004 23236 2010 23248
rect 8481 23239 8539 23245
rect 8481 23236 8493 23239
rect 2004 23208 8493 23236
rect 2004 23196 2010 23208
rect 8481 23205 8493 23208
rect 8527 23236 8539 23239
rect 8570 23236 8576 23248
rect 8527 23208 8576 23236
rect 8527 23205 8539 23208
rect 8481 23199 8539 23205
rect 8570 23196 8576 23208
rect 8628 23196 8634 23248
rect 9858 23236 9864 23248
rect 9819 23208 9864 23236
rect 9858 23196 9864 23208
rect 9916 23196 9922 23248
rect 14642 23196 14648 23248
rect 14700 23236 14706 23248
rect 14700 23208 16481 23236
rect 14700 23196 14706 23208
rect 1394 23168 1400 23180
rect 1355 23140 1400 23168
rect 1394 23128 1400 23140
rect 1452 23128 1458 23180
rect 7190 23128 7196 23180
rect 7248 23168 7254 23180
rect 7285 23171 7343 23177
rect 7285 23168 7297 23171
rect 7248 23140 7297 23168
rect 7248 23128 7254 23140
rect 7285 23137 7297 23140
rect 7331 23137 7343 23171
rect 7285 23131 7343 23137
rect 11241 23171 11299 23177
rect 11241 23137 11253 23171
rect 11287 23168 11299 23171
rect 11330 23168 11336 23180
rect 11287 23140 11336 23168
rect 11287 23137 11299 23140
rect 11241 23131 11299 23137
rect 11330 23128 11336 23140
rect 11388 23128 11394 23180
rect 12158 23128 12164 23180
rect 12216 23168 12222 23180
rect 12288 23171 12346 23177
rect 12288 23168 12300 23171
rect 12216 23140 12300 23168
rect 12216 23128 12222 23140
rect 12288 23137 12300 23140
rect 12334 23137 12346 23171
rect 12288 23131 12346 23137
rect 13608 23171 13666 23177
rect 13608 23137 13620 23171
rect 13654 23168 13666 23171
rect 13814 23168 13820 23180
rect 13654 23140 13820 23168
rect 13654 23137 13666 23140
rect 13608 23131 13666 23137
rect 13814 23128 13820 23140
rect 13872 23128 13878 23180
rect 15378 23168 15384 23180
rect 15339 23140 15384 23168
rect 15378 23128 15384 23140
rect 15436 23128 15442 23180
rect 16453 23168 16481 23208
rect 16758 23168 16764 23180
rect 16816 23177 16822 23180
rect 16816 23171 16854 23177
rect 16453 23140 16764 23168
rect 16758 23128 16764 23140
rect 16842 23137 16854 23171
rect 18046 23168 18052 23180
rect 18007 23140 18052 23168
rect 16816 23131 16854 23137
rect 16816 23128 16822 23131
rect 18046 23128 18052 23140
rect 18104 23128 18110 23180
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 9214 23060 9220 23112
rect 9272 23100 9278 23112
rect 9769 23103 9827 23109
rect 9769 23100 9781 23103
rect 9272 23072 9781 23100
rect 9272 23060 9278 23072
rect 9769 23069 9781 23072
rect 9815 23069 9827 23103
rect 10042 23100 10048 23112
rect 10003 23072 10048 23100
rect 9769 23063 9827 23069
rect 10042 23060 10048 23072
rect 10100 23060 10106 23112
rect 6270 22992 6276 23044
rect 6328 23032 6334 23044
rect 12986 23032 12992 23044
rect 6328 23004 12992 23032
rect 6328 22992 6334 23004
rect 12986 22992 12992 23004
rect 13044 22992 13050 23044
rect 7282 22924 7288 22976
rect 7340 22964 7346 22976
rect 7423 22967 7481 22973
rect 7423 22964 7435 22967
rect 7340 22936 7435 22964
rect 7340 22924 7346 22936
rect 7423 22933 7435 22936
rect 7469 22933 7481 22967
rect 7742 22964 7748 22976
rect 7703 22936 7748 22964
rect 7423 22927 7481 22933
rect 7742 22924 7748 22936
rect 7800 22924 7806 22976
rect 8711 22967 8769 22973
rect 8711 22933 8723 22967
rect 8757 22964 8769 22967
rect 8846 22964 8852 22976
rect 8757 22936 8852 22964
rect 8757 22933 8769 22936
rect 8711 22927 8769 22933
rect 8846 22924 8852 22936
rect 8904 22924 8910 22976
rect 11054 22924 11060 22976
rect 11112 22964 11118 22976
rect 11379 22967 11437 22973
rect 11379 22964 11391 22967
rect 11112 22936 11391 22964
rect 11112 22924 11118 22936
rect 11379 22933 11391 22936
rect 11425 22933 11437 22967
rect 11379 22927 11437 22933
rect 12391 22967 12449 22973
rect 12391 22933 12403 22967
rect 12437 22964 12449 22967
rect 12526 22964 12532 22976
rect 12437 22936 12532 22964
rect 12437 22933 12449 22936
rect 12391 22927 12449 22933
rect 12526 22924 12532 22936
rect 12584 22924 12590 22976
rect 15611 22967 15669 22973
rect 15611 22933 15623 22967
rect 15657 22964 15669 22967
rect 15930 22964 15936 22976
rect 15657 22936 15936 22964
rect 15657 22933 15669 22936
rect 15611 22927 15669 22933
rect 15930 22924 15936 22936
rect 15988 22924 15994 22976
rect 16899 22967 16957 22973
rect 16899 22933 16911 22967
rect 16945 22964 16957 22967
rect 17586 22964 17592 22976
rect 16945 22936 17592 22964
rect 16945 22933 16957 22936
rect 16899 22927 16957 22933
rect 17586 22924 17592 22936
rect 17644 22924 17650 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1210 22720 1216 22772
rect 1268 22760 1274 22772
rect 1581 22763 1639 22769
rect 1581 22760 1593 22763
rect 1268 22732 1593 22760
rect 1268 22720 1274 22732
rect 1581 22729 1593 22732
rect 1627 22729 1639 22763
rect 7190 22760 7196 22772
rect 7103 22732 7196 22760
rect 1581 22723 1639 22729
rect 7190 22720 7196 22732
rect 7248 22760 7254 22772
rect 8202 22760 8208 22772
rect 7248 22732 8208 22760
rect 7248 22720 7254 22732
rect 8202 22720 8208 22732
rect 8260 22720 8266 22772
rect 8570 22760 8576 22772
rect 8531 22732 8576 22760
rect 8570 22720 8576 22732
rect 8628 22720 8634 22772
rect 9858 22720 9864 22772
rect 9916 22760 9922 22772
rect 10229 22763 10287 22769
rect 10229 22760 10241 22763
rect 9916 22732 10241 22760
rect 9916 22720 9922 22732
rect 10229 22729 10241 22732
rect 10275 22729 10287 22763
rect 10229 22723 10287 22729
rect 11514 22720 11520 22772
rect 11572 22760 11578 22772
rect 13078 22760 13084 22772
rect 11572 22732 13084 22760
rect 11572 22720 11578 22732
rect 13078 22720 13084 22732
rect 13136 22760 13142 22772
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 13136 22732 14933 22760
rect 13136 22720 13142 22732
rect 7742 22692 7748 22704
rect 7392 22664 7748 22692
rect 1026 22584 1032 22636
rect 1084 22624 1090 22636
rect 7392 22633 7420 22664
rect 7742 22652 7748 22664
rect 7800 22652 7806 22704
rect 9214 22652 9220 22704
rect 9272 22692 9278 22704
rect 10597 22695 10655 22701
rect 10597 22692 10609 22695
rect 9272 22664 10609 22692
rect 9272 22652 9278 22664
rect 10597 22661 10609 22664
rect 10643 22661 10655 22695
rect 11330 22692 11336 22704
rect 11243 22664 11336 22692
rect 10597 22655 10655 22661
rect 11330 22652 11336 22664
rect 11388 22692 11394 22704
rect 13446 22692 13452 22704
rect 11388 22664 13452 22692
rect 11388 22652 11394 22664
rect 13446 22652 13452 22664
rect 13504 22652 13510 22704
rect 7377 22627 7435 22633
rect 1084 22596 4154 22624
rect 1084 22584 1090 22596
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 1946 22556 1952 22568
rect 1443 22528 1952 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 1946 22516 1952 22528
rect 2004 22516 2010 22568
rect 4126 22556 4154 22596
rect 7377 22593 7389 22627
rect 7423 22593 7435 22627
rect 7377 22587 7435 22593
rect 7558 22584 7564 22636
rect 7616 22624 7622 22636
rect 7653 22627 7711 22633
rect 7653 22624 7665 22627
rect 7616 22596 7665 22624
rect 7616 22584 7622 22596
rect 7653 22593 7665 22596
rect 7699 22593 7711 22627
rect 9582 22624 9588 22636
rect 9543 22596 9588 22624
rect 7653 22587 7711 22593
rect 9582 22584 9588 22596
rect 9640 22624 9646 22636
rect 10042 22624 10048 22636
rect 9640 22596 10048 22624
rect 9640 22584 9646 22596
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 13814 22584 13820 22636
rect 13872 22624 13878 22636
rect 14277 22627 14335 22633
rect 14277 22624 14289 22627
rect 13872 22596 14289 22624
rect 13872 22584 13878 22596
rect 14277 22593 14289 22596
rect 14323 22593 14335 22627
rect 14277 22587 14335 22593
rect 10870 22565 10876 22568
rect 5756 22559 5814 22565
rect 5756 22556 5768 22559
rect 4126 22528 5768 22556
rect 5756 22525 5768 22528
rect 5802 22525 5814 22559
rect 5756 22519 5814 22525
rect 10848 22559 10876 22565
rect 10848 22525 10860 22559
rect 10928 22556 10934 22568
rect 11609 22559 11667 22565
rect 11609 22556 11621 22559
rect 10928 22528 11621 22556
rect 10848 22519 10876 22525
rect 5771 22420 5799 22519
rect 10870 22516 10876 22519
rect 10928 22516 10934 22528
rect 11609 22525 11621 22528
rect 11655 22556 11667 22559
rect 12158 22556 12164 22568
rect 11655 22528 12164 22556
rect 11655 22525 11667 22528
rect 11609 22519 11667 22525
rect 12158 22516 12164 22528
rect 12216 22556 12222 22568
rect 12434 22556 12440 22568
rect 12216 22528 12296 22556
rect 12395 22528 12440 22556
rect 12216 22516 12222 22528
rect 5859 22491 5917 22497
rect 5859 22457 5871 22491
rect 5905 22488 5917 22491
rect 6454 22488 6460 22500
rect 5905 22460 6460 22488
rect 5905 22457 5917 22460
rect 5859 22451 5917 22457
rect 6454 22448 6460 22460
rect 6512 22448 6518 22500
rect 6641 22491 6699 22497
rect 6641 22457 6653 22491
rect 6687 22488 6699 22491
rect 7469 22491 7527 22497
rect 6687 22460 7328 22488
rect 6687 22457 6699 22460
rect 6641 22451 6699 22457
rect 6273 22423 6331 22429
rect 6273 22420 6285 22423
rect 5771 22392 6285 22420
rect 6273 22389 6285 22392
rect 6319 22420 6331 22423
rect 7098 22420 7104 22432
rect 6319 22392 7104 22420
rect 6319 22389 6331 22392
rect 6273 22383 6331 22389
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 7300 22420 7328 22460
rect 7469 22457 7481 22491
rect 7515 22488 7527 22491
rect 7742 22488 7748 22500
rect 7515 22460 7748 22488
rect 7515 22457 7527 22460
rect 7469 22451 7527 22457
rect 7484 22420 7512 22451
rect 7742 22448 7748 22460
rect 7800 22448 7806 22500
rect 9306 22488 9312 22500
rect 9267 22460 9312 22488
rect 9306 22448 9312 22460
rect 9364 22448 9370 22500
rect 9401 22491 9459 22497
rect 9401 22457 9413 22491
rect 9447 22457 9459 22491
rect 12268 22488 12296 22528
rect 12434 22516 12440 22528
rect 12492 22556 12498 22568
rect 13265 22559 13323 22565
rect 13265 22556 13277 22559
rect 12492 22528 13277 22556
rect 12492 22516 12498 22528
rect 13265 22525 13277 22528
rect 13311 22525 13323 22559
rect 13265 22519 13323 22525
rect 13516 22559 13574 22565
rect 13516 22525 13528 22559
rect 13562 22556 13574 22559
rect 13998 22556 14004 22568
rect 13562 22528 14004 22556
rect 13562 22525 13574 22528
rect 13516 22519 13574 22525
rect 13998 22516 14004 22528
rect 14056 22516 14062 22568
rect 14511 22565 14539 22732
rect 14921 22729 14933 22732
rect 14967 22729 14979 22763
rect 16758 22760 16764 22772
rect 16719 22732 16764 22760
rect 14921 22723 14979 22729
rect 16758 22720 16764 22732
rect 16816 22720 16822 22772
rect 17083 22695 17141 22701
rect 17083 22661 17095 22695
rect 17129 22692 17141 22695
rect 18046 22692 18052 22704
rect 17129 22664 18052 22692
rect 17129 22661 17141 22664
rect 17083 22655 17141 22661
rect 18046 22652 18052 22664
rect 18104 22692 18110 22704
rect 18233 22695 18291 22701
rect 18233 22692 18245 22695
rect 18104 22664 18245 22692
rect 18104 22652 18110 22664
rect 18233 22661 18245 22664
rect 18279 22661 18291 22695
rect 18233 22655 18291 22661
rect 14496 22559 14554 22565
rect 14496 22525 14508 22559
rect 14542 22525 14554 22559
rect 14496 22519 14554 22525
rect 16850 22516 16856 22568
rect 16908 22556 16914 22568
rect 17012 22559 17070 22565
rect 17012 22556 17024 22559
rect 16908 22528 17024 22556
rect 16908 22516 16914 22528
rect 17012 22525 17024 22528
rect 17058 22556 17070 22559
rect 17405 22559 17463 22565
rect 17405 22556 17417 22559
rect 17058 22528 17417 22556
rect 17058 22525 17070 22528
rect 17012 22519 17070 22525
rect 17405 22525 17417 22528
rect 17451 22525 17463 22559
rect 17405 22519 17463 22525
rect 12897 22491 12955 22497
rect 12897 22488 12909 22491
rect 12268 22460 12909 22488
rect 9401 22451 9459 22457
rect 12897 22457 12909 22460
rect 12943 22457 12955 22491
rect 12897 22451 12955 22457
rect 9030 22420 9036 22432
rect 7300 22392 7512 22420
rect 8991 22392 9036 22420
rect 9030 22380 9036 22392
rect 9088 22420 9094 22432
rect 9416 22420 9444 22451
rect 13722 22448 13728 22500
rect 13780 22488 13786 22500
rect 14599 22491 14657 22497
rect 14599 22488 14611 22491
rect 13780 22460 14611 22488
rect 13780 22448 13786 22460
rect 14599 22457 14611 22460
rect 14645 22457 14657 22491
rect 14599 22451 14657 22457
rect 15378 22448 15384 22500
rect 15436 22488 15442 22500
rect 15565 22491 15623 22497
rect 15565 22488 15577 22491
rect 15436 22460 15577 22488
rect 15436 22448 15442 22460
rect 15565 22457 15577 22460
rect 15611 22488 15623 22491
rect 22370 22488 22376 22500
rect 15611 22460 22376 22488
rect 15611 22457 15623 22460
rect 15565 22451 15623 22457
rect 22370 22448 22376 22460
rect 22428 22448 22434 22500
rect 9088 22392 9444 22420
rect 9088 22380 9094 22392
rect 10778 22380 10784 22432
rect 10836 22420 10842 22432
rect 10919 22423 10977 22429
rect 10919 22420 10931 22423
rect 10836 22392 10931 22420
rect 10836 22380 10842 22392
rect 10919 22389 10931 22392
rect 10965 22389 10977 22423
rect 12618 22420 12624 22432
rect 12579 22392 12624 22420
rect 10919 22383 10977 22389
rect 12618 22380 12624 22392
rect 12676 22380 12682 22432
rect 13354 22380 13360 22432
rect 13412 22420 13418 22432
rect 13587 22423 13645 22429
rect 13587 22420 13599 22423
rect 13412 22392 13599 22420
rect 13412 22380 13418 22392
rect 13587 22389 13599 22392
rect 13633 22389 13645 22423
rect 15654 22420 15660 22432
rect 15615 22392 15660 22420
rect 13587 22383 13645 22389
rect 15654 22380 15660 22392
rect 15712 22380 15718 22432
rect 23474 22380 23480 22432
rect 23532 22420 23538 22432
rect 24581 22423 24639 22429
rect 24581 22420 24593 22423
rect 23532 22392 24593 22420
rect 23532 22380 23538 22392
rect 24581 22389 24593 22392
rect 24627 22420 24639 22423
rect 24670 22420 24676 22432
rect 24627 22392 24676 22420
rect 24627 22389 24639 22392
rect 24581 22383 24639 22389
rect 24670 22380 24676 22392
rect 24728 22380 24734 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1394 22176 1400 22228
rect 1452 22216 1458 22228
rect 1673 22219 1731 22225
rect 1673 22216 1685 22219
rect 1452 22188 1685 22216
rect 1452 22176 1458 22188
rect 1673 22185 1685 22188
rect 1719 22216 1731 22219
rect 6319 22219 6377 22225
rect 6319 22216 6331 22219
rect 1719 22188 6331 22216
rect 1719 22185 1731 22188
rect 1673 22179 1731 22185
rect 6319 22185 6331 22188
rect 6365 22185 6377 22219
rect 8846 22216 8852 22228
rect 8807 22188 8852 22216
rect 6319 22179 6377 22185
rect 8846 22176 8852 22188
rect 8904 22176 8910 22228
rect 11054 22216 11060 22228
rect 11015 22188 11060 22216
rect 11054 22176 11060 22188
rect 11112 22176 11118 22228
rect 12437 22219 12495 22225
rect 12437 22185 12449 22219
rect 12483 22216 12495 22219
rect 12526 22216 12532 22228
rect 12483 22188 12532 22216
rect 12483 22185 12495 22188
rect 12437 22179 12495 22185
rect 12526 22176 12532 22188
rect 12584 22216 12590 22228
rect 12584 22188 13216 22216
rect 12584 22176 12590 22188
rect 6822 22108 6828 22160
rect 6880 22148 6886 22160
rect 7377 22151 7435 22157
rect 7377 22148 7389 22151
rect 6880 22120 7389 22148
rect 6880 22108 6886 22120
rect 7377 22117 7389 22120
rect 7423 22117 7435 22151
rect 10134 22148 10140 22160
rect 10095 22120 10140 22148
rect 7377 22111 7435 22117
rect 10134 22108 10140 22120
rect 10192 22108 10198 22160
rect 13188 22157 13216 22188
rect 13446 22176 13452 22228
rect 13504 22216 13510 22228
rect 15286 22216 15292 22228
rect 13504 22188 15292 22216
rect 13504 22176 13510 22188
rect 15286 22176 15292 22188
rect 15344 22176 15350 22228
rect 13173 22151 13231 22157
rect 13173 22117 13185 22151
rect 13219 22117 13231 22151
rect 13173 22111 13231 22117
rect 13262 22108 13268 22160
rect 13320 22148 13326 22160
rect 13320 22120 13365 22148
rect 13320 22108 13326 22120
rect 15746 22108 15752 22160
rect 15804 22148 15810 22160
rect 16117 22151 16175 22157
rect 16117 22148 16129 22151
rect 15804 22120 16129 22148
rect 15804 22108 15810 22120
rect 16117 22117 16129 22120
rect 16163 22117 16175 22151
rect 16117 22111 16175 22117
rect 6178 22080 6184 22092
rect 6139 22052 6184 22080
rect 6178 22040 6184 22052
rect 6236 22040 6242 22092
rect 11514 22080 11520 22092
rect 11475 22052 11520 22080
rect 11514 22040 11520 22052
rect 11572 22040 11578 22092
rect 5169 22015 5227 22021
rect 5169 21981 5181 22015
rect 5215 22012 5227 22015
rect 6638 22012 6644 22024
rect 5215 21984 6644 22012
rect 5215 21981 5227 21984
rect 5169 21975 5227 21981
rect 6638 21972 6644 21984
rect 6696 21972 6702 22024
rect 7285 22015 7343 22021
rect 7285 21981 7297 22015
rect 7331 22012 7343 22015
rect 7374 22012 7380 22024
rect 7331 21984 7380 22012
rect 7331 21981 7343 21984
rect 7285 21975 7343 21981
rect 7374 21972 7380 21984
rect 7432 21972 7438 22024
rect 7558 22012 7564 22024
rect 7519 21984 7564 22012
rect 7558 21972 7564 21984
rect 7616 21972 7622 22024
rect 9490 21972 9496 22024
rect 9548 22012 9554 22024
rect 10045 22015 10103 22021
rect 10045 22012 10057 22015
rect 9548 21984 10057 22012
rect 9548 21972 9554 21984
rect 10045 21981 10057 21984
rect 10091 22012 10103 22015
rect 10778 22012 10784 22024
rect 10091 21984 10784 22012
rect 10091 21981 10103 21984
rect 10045 21975 10103 21981
rect 10778 21972 10784 21984
rect 10836 21972 10842 22024
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 22012 16083 22015
rect 16942 22012 16948 22024
rect 16071 21984 16948 22012
rect 16071 21981 16083 21984
rect 16025 21975 16083 21981
rect 16942 21972 16948 21984
rect 17000 21972 17006 22024
rect 8662 21904 8668 21956
rect 8720 21944 8726 21956
rect 9582 21944 9588 21956
rect 8720 21916 9588 21944
rect 8720 21904 8726 21916
rect 9582 21904 9588 21916
rect 9640 21944 9646 21956
rect 10597 21947 10655 21953
rect 10597 21944 10609 21947
rect 9640 21916 10609 21944
rect 9640 21904 9646 21916
rect 10597 21913 10609 21916
rect 10643 21913 10655 21947
rect 13722 21944 13728 21956
rect 13683 21916 13728 21944
rect 10597 21907 10655 21913
rect 13722 21904 13728 21916
rect 13780 21944 13786 21956
rect 14277 21947 14335 21953
rect 14277 21944 14289 21947
rect 13780 21916 14289 21944
rect 13780 21904 13786 21916
rect 14277 21913 14289 21916
rect 14323 21913 14335 21947
rect 14277 21907 14335 21913
rect 16482 21904 16488 21956
rect 16540 21944 16546 21956
rect 16577 21947 16635 21953
rect 16577 21944 16589 21947
rect 16540 21916 16589 21944
rect 16540 21904 16546 21916
rect 16577 21913 16589 21916
rect 16623 21913 16635 21947
rect 16577 21907 16635 21913
rect 9306 21876 9312 21888
rect 9219 21848 9312 21876
rect 9306 21836 9312 21848
rect 9364 21876 9370 21888
rect 11655 21879 11713 21885
rect 11655 21876 11667 21879
rect 9364 21848 11667 21876
rect 9364 21836 9370 21848
rect 11655 21845 11667 21848
rect 11701 21845 11713 21879
rect 12802 21876 12808 21888
rect 12763 21848 12808 21876
rect 11655 21839 11713 21845
rect 12802 21836 12808 21848
rect 12860 21836 12866 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 7650 21632 7656 21684
rect 7708 21672 7714 21684
rect 11514 21672 11520 21684
rect 7708 21644 11520 21672
rect 7708 21632 7714 21644
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 13262 21632 13268 21684
rect 13320 21672 13326 21684
rect 13725 21675 13783 21681
rect 13725 21672 13737 21675
rect 13320 21644 13737 21672
rect 13320 21632 13326 21644
rect 13725 21641 13737 21644
rect 13771 21641 13783 21675
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 13725 21635 13783 21641
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 7006 21564 7012 21616
rect 7064 21604 7070 21616
rect 7064 21576 7788 21604
rect 7064 21564 7070 21576
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 6178 21536 6184 21548
rect 5675 21508 6184 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 6178 21496 6184 21508
rect 6236 21536 6242 21548
rect 7558 21536 7564 21548
rect 6236 21508 7564 21536
rect 6236 21496 6242 21508
rect 7558 21496 7564 21508
rect 7616 21496 7622 21548
rect 7760 21536 7788 21576
rect 7834 21564 7840 21616
rect 7892 21604 7898 21616
rect 10965 21607 11023 21613
rect 10965 21604 10977 21607
rect 7892 21576 10977 21604
rect 7892 21564 7898 21576
rect 9140 21548 9168 21576
rect 10965 21573 10977 21576
rect 11011 21573 11023 21607
rect 10965 21567 11023 21573
rect 12253 21607 12311 21613
rect 12253 21573 12265 21607
rect 12299 21604 12311 21607
rect 13354 21604 13360 21616
rect 12299 21576 13360 21604
rect 12299 21573 12311 21576
rect 12253 21567 12311 21573
rect 8205 21539 8263 21545
rect 8205 21536 8217 21539
rect 7760 21508 8217 21536
rect 8205 21505 8217 21508
rect 8251 21536 8263 21539
rect 8662 21536 8668 21548
rect 8251 21508 8668 21536
rect 8251 21505 8263 21508
rect 8205 21499 8263 21505
rect 8662 21496 8668 21508
rect 8720 21496 8726 21548
rect 8846 21536 8852 21548
rect 8807 21508 8852 21536
rect 8846 21496 8852 21508
rect 8904 21496 8910 21548
rect 9122 21536 9128 21548
rect 9035 21508 9128 21536
rect 9122 21496 9128 21508
rect 9180 21496 9186 21548
rect 10413 21539 10471 21545
rect 10413 21505 10425 21539
rect 10459 21536 10471 21539
rect 11054 21536 11060 21548
rect 10459 21508 11060 21536
rect 10459 21505 10471 21508
rect 10413 21499 10471 21505
rect 11054 21496 11060 21508
rect 11112 21496 11118 21548
rect 12820 21545 12848 21576
rect 13354 21564 13360 21576
rect 13412 21564 13418 21616
rect 13538 21564 13544 21616
rect 13596 21604 13602 21616
rect 14921 21607 14979 21613
rect 13596 21576 14872 21604
rect 13596 21564 13602 21576
rect 12805 21539 12863 21545
rect 12805 21505 12817 21539
rect 12851 21505 12863 21539
rect 12805 21499 12863 21505
rect 13449 21539 13507 21545
rect 13449 21505 13461 21539
rect 13495 21536 13507 21539
rect 13722 21536 13728 21548
rect 13495 21508 13728 21536
rect 13495 21505 13507 21508
rect 13449 21499 13507 21505
rect 13722 21496 13728 21508
rect 13780 21536 13786 21548
rect 14366 21536 14372 21548
rect 13780 21508 14372 21536
rect 13780 21496 13786 21508
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 14844 21536 14872 21576
rect 14921 21573 14933 21607
rect 14967 21604 14979 21607
rect 16850 21604 16856 21616
rect 14967 21576 16856 21604
rect 14967 21573 14979 21576
rect 14921 21567 14979 21573
rect 16850 21564 16856 21576
rect 16908 21564 16914 21616
rect 15657 21539 15715 21545
rect 15657 21536 15669 21539
rect 14844 21508 15669 21536
rect 15657 21505 15669 21508
rect 15703 21536 15715 21539
rect 15746 21536 15752 21548
rect 15703 21508 15752 21536
rect 15703 21505 15715 21508
rect 15657 21499 15715 21505
rect 15746 21496 15752 21508
rect 15804 21496 15810 21548
rect 15930 21536 15936 21548
rect 15891 21508 15936 21536
rect 15930 21496 15936 21508
rect 15988 21536 15994 21548
rect 17221 21539 17279 21545
rect 17221 21536 17233 21539
rect 15988 21508 17233 21536
rect 15988 21496 15994 21508
rect 17221 21505 17233 21508
rect 17267 21505 17279 21539
rect 17221 21499 17279 21505
rect 658 21428 664 21480
rect 716 21468 722 21480
rect 1397 21471 1455 21477
rect 1397 21468 1409 21471
rect 716 21440 1409 21468
rect 716 21428 722 21440
rect 1397 21437 1409 21440
rect 1443 21468 1455 21471
rect 1949 21471 2007 21477
rect 1949 21468 1961 21471
rect 1443 21440 1961 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 1949 21437 1961 21440
rect 1995 21437 2007 21471
rect 1949 21431 2007 21437
rect 4560 21471 4618 21477
rect 4560 21437 4572 21471
rect 4606 21437 4618 21471
rect 4560 21431 4618 21437
rect 4663 21471 4721 21477
rect 4663 21437 4675 21471
rect 4709 21468 4721 21471
rect 4982 21468 4988 21480
rect 4709 21440 4988 21468
rect 4709 21437 4721 21440
rect 4663 21431 4721 21437
rect 4575 21332 4603 21431
rect 4982 21428 4988 21440
rect 5040 21428 5046 21480
rect 5772 21471 5830 21477
rect 5772 21437 5784 21471
rect 5818 21468 5830 21471
rect 6270 21468 6276 21480
rect 5818 21440 6276 21468
rect 5818 21437 5830 21440
rect 5772 21431 5830 21437
rect 6270 21428 6276 21440
rect 6328 21428 6334 21480
rect 18138 21477 18144 21480
rect 18116 21471 18144 21477
rect 18116 21468 18128 21471
rect 18051 21440 18128 21468
rect 18116 21437 18128 21440
rect 18196 21468 18202 21480
rect 18509 21471 18567 21477
rect 18509 21468 18521 21471
rect 18196 21440 18521 21468
rect 18116 21431 18144 21437
rect 18138 21428 18144 21431
rect 18196 21428 18202 21440
rect 18509 21437 18521 21440
rect 18555 21468 18567 21471
rect 22002 21468 22008 21480
rect 18555 21440 22008 21468
rect 18555 21437 18567 21440
rect 18509 21431 18567 21437
rect 22002 21428 22008 21440
rect 22060 21428 22066 21480
rect 24581 21471 24639 21477
rect 24581 21437 24593 21471
rect 24627 21468 24639 21471
rect 25130 21468 25136 21480
rect 24627 21440 25136 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 25130 21428 25136 21440
rect 25188 21428 25194 21480
rect 5859 21403 5917 21409
rect 5859 21369 5871 21403
rect 5905 21400 5917 21403
rect 6914 21400 6920 21412
rect 5905 21372 6920 21400
rect 5905 21369 5917 21372
rect 5859 21363 5917 21369
rect 6914 21360 6920 21372
rect 6972 21360 6978 21412
rect 7006 21360 7012 21412
rect 7064 21400 7070 21412
rect 7285 21403 7343 21409
rect 7285 21400 7297 21403
rect 7064 21372 7297 21400
rect 7064 21360 7070 21372
rect 7285 21369 7297 21372
rect 7331 21369 7343 21403
rect 7285 21363 7343 21369
rect 7374 21360 7380 21412
rect 7432 21400 7438 21412
rect 8941 21403 8999 21409
rect 7432 21372 7477 21400
rect 7432 21360 7438 21372
rect 8941 21369 8953 21403
rect 8987 21400 8999 21403
rect 9030 21400 9036 21412
rect 8987 21372 9036 21400
rect 8987 21369 8999 21372
rect 8941 21363 8999 21369
rect 5074 21332 5080 21344
rect 4575 21304 5080 21332
rect 5074 21292 5080 21304
rect 5132 21292 5138 21344
rect 6641 21335 6699 21341
rect 6641 21301 6653 21335
rect 6687 21332 6699 21335
rect 6822 21332 6828 21344
rect 6687 21304 6828 21332
rect 6687 21301 6699 21304
rect 6641 21295 6699 21301
rect 6822 21292 6828 21304
rect 6880 21292 6886 21344
rect 7101 21335 7159 21341
rect 7101 21301 7113 21335
rect 7147 21332 7159 21335
rect 7190 21332 7196 21344
rect 7147 21304 7196 21332
rect 7147 21301 7159 21304
rect 7101 21295 7159 21301
rect 7190 21292 7196 21304
rect 7248 21292 7254 21344
rect 8570 21332 8576 21344
rect 8531 21304 8576 21332
rect 8570 21292 8576 21304
rect 8628 21332 8634 21344
rect 8956 21332 8984 21363
rect 9030 21360 9036 21372
rect 9088 21360 9094 21412
rect 10505 21403 10563 21409
rect 10505 21400 10517 21403
rect 10152 21372 10517 21400
rect 10152 21344 10180 21372
rect 10505 21369 10517 21372
rect 10551 21369 10563 21403
rect 10505 21363 10563 21369
rect 12802 21360 12808 21412
rect 12860 21400 12866 21412
rect 12897 21403 12955 21409
rect 12897 21400 12909 21403
rect 12860 21372 12909 21400
rect 12860 21360 12866 21372
rect 12897 21369 12909 21372
rect 12943 21400 12955 21403
rect 13538 21400 13544 21412
rect 12943 21372 13544 21400
rect 12943 21369 12955 21372
rect 12897 21363 12955 21369
rect 13538 21360 13544 21372
rect 13596 21360 13602 21412
rect 14461 21403 14519 21409
rect 14461 21369 14473 21403
rect 14507 21369 14519 21403
rect 16022 21400 16028 21412
rect 14461 21363 14519 21369
rect 15304 21372 16028 21400
rect 8628 21304 8984 21332
rect 9861 21335 9919 21341
rect 8628 21292 8634 21304
rect 9861 21301 9873 21335
rect 9907 21332 9919 21335
rect 10134 21332 10140 21344
rect 9907 21304 10140 21332
rect 9907 21301 9919 21304
rect 9861 21295 9919 21301
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 14182 21332 14188 21344
rect 14095 21304 14188 21332
rect 14182 21292 14188 21304
rect 14240 21332 14246 21344
rect 14476 21332 14504 21363
rect 14240 21304 14504 21332
rect 14240 21292 14246 21304
rect 14550 21292 14556 21344
rect 14608 21332 14614 21344
rect 15304 21341 15332 21372
rect 16022 21360 16028 21372
rect 16080 21360 16086 21412
rect 16390 21360 16396 21412
rect 16448 21400 16454 21412
rect 16577 21403 16635 21409
rect 16577 21400 16589 21403
rect 16448 21372 16589 21400
rect 16448 21360 16454 21372
rect 16577 21369 16589 21372
rect 16623 21369 16635 21403
rect 16577 21363 16635 21369
rect 15289 21335 15347 21341
rect 15289 21332 15301 21335
rect 14608 21304 15301 21332
rect 14608 21292 14614 21304
rect 15289 21301 15301 21304
rect 15335 21301 15347 21335
rect 16942 21332 16948 21344
rect 16903 21304 16948 21332
rect 15289 21295 15347 21301
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 17494 21292 17500 21344
rect 17552 21332 17558 21344
rect 18187 21335 18245 21341
rect 18187 21332 18199 21335
rect 17552 21304 18199 21332
rect 17552 21292 17558 21304
rect 18187 21301 18199 21304
rect 18233 21301 18245 21335
rect 18187 21295 18245 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 5258 21128 5264 21140
rect 5219 21100 5264 21128
rect 5258 21088 5264 21100
rect 5316 21088 5322 21140
rect 6546 21088 6552 21140
rect 6604 21128 6610 21140
rect 6825 21131 6883 21137
rect 6825 21128 6837 21131
rect 6604 21100 6837 21128
rect 6604 21088 6610 21100
rect 6825 21097 6837 21100
rect 6871 21097 6883 21131
rect 6825 21091 6883 21097
rect 7190 21088 7196 21140
rect 7248 21128 7254 21140
rect 7374 21128 7380 21140
rect 7248 21100 7380 21128
rect 7248 21088 7254 21100
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 7466 21088 7472 21140
rect 7524 21128 7530 21140
rect 8021 21131 8079 21137
rect 8021 21128 8033 21131
rect 7524 21100 8033 21128
rect 7524 21088 7530 21100
rect 8021 21097 8033 21100
rect 8067 21097 8079 21131
rect 8021 21091 8079 21097
rect 8711 21131 8769 21137
rect 8711 21097 8723 21131
rect 8757 21128 8769 21131
rect 9214 21128 9220 21140
rect 8757 21100 9220 21128
rect 8757 21097 8769 21100
rect 8711 21091 8769 21097
rect 2038 21020 2044 21072
rect 2096 21060 2102 21072
rect 8036 21060 8064 21091
rect 9214 21088 9220 21100
rect 9272 21088 9278 21140
rect 9490 21128 9496 21140
rect 9451 21100 9496 21128
rect 9490 21088 9496 21100
rect 9548 21088 9554 21140
rect 13262 21088 13268 21140
rect 13320 21128 13326 21140
rect 13906 21128 13912 21140
rect 13320 21100 13912 21128
rect 13320 21088 13326 21100
rect 13906 21088 13912 21100
rect 13964 21128 13970 21140
rect 15838 21128 15844 21140
rect 13964 21100 15844 21128
rect 13964 21088 13970 21100
rect 15838 21088 15844 21100
rect 15896 21128 15902 21140
rect 15896 21100 16068 21128
rect 15896 21088 15902 21100
rect 2096 21032 6684 21060
rect 8036 21032 9628 21060
rect 2096 21020 2102 21032
rect 4430 20992 4436 21004
rect 4391 20964 4436 20992
rect 4430 20952 4436 20964
rect 4488 20952 4494 21004
rect 5074 20952 5080 21004
rect 5132 20992 5138 21004
rect 5512 20995 5570 21001
rect 5512 20992 5524 20995
rect 5132 20964 5524 20992
rect 5132 20952 5138 20964
rect 5512 20961 5524 20964
rect 5558 20992 5570 20995
rect 6178 20992 6184 21004
rect 5558 20964 6184 20992
rect 5558 20961 5570 20964
rect 5512 20955 5570 20961
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6656 20992 6684 21032
rect 8478 20992 8484 21004
rect 6656 20964 8484 20992
rect 8478 20952 8484 20964
rect 8536 20992 8542 21004
rect 8640 20995 8698 21001
rect 8640 20992 8652 20995
rect 8536 20964 8652 20992
rect 8536 20952 8542 20964
rect 8640 20961 8652 20964
rect 8686 20992 8698 20995
rect 8686 20964 9536 20992
rect 8686 20961 8698 20964
rect 8640 20955 8698 20961
rect 9508 20936 9536 20964
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20893 6515 20927
rect 6457 20887 6515 20893
rect 4614 20788 4620 20800
rect 4575 20760 4620 20788
rect 4614 20748 4620 20760
rect 4672 20748 4678 20800
rect 5583 20791 5641 20797
rect 5583 20757 5595 20791
rect 5629 20788 5641 20791
rect 5994 20788 6000 20800
rect 5629 20760 6000 20788
rect 5629 20757 5641 20760
rect 5583 20751 5641 20757
rect 5994 20748 6000 20760
rect 6052 20748 6058 20800
rect 6270 20788 6276 20800
rect 6231 20760 6276 20788
rect 6270 20748 6276 20760
rect 6328 20788 6334 20800
rect 6472 20788 6500 20887
rect 9490 20884 9496 20936
rect 9548 20884 9554 20936
rect 9600 20856 9628 21032
rect 9858 21020 9864 21072
rect 9916 21060 9922 21072
rect 10597 21063 10655 21069
rect 10597 21060 10609 21063
rect 9916 21032 10609 21060
rect 9916 21020 9922 21032
rect 10597 21029 10609 21032
rect 10643 21060 10655 21063
rect 11146 21060 11152 21072
rect 10643 21032 11152 21060
rect 10643 21029 10655 21032
rect 10597 21023 10655 21029
rect 11146 21020 11152 21032
rect 11204 21020 11210 21072
rect 13722 21060 13728 21072
rect 13683 21032 13728 21060
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 13814 21020 13820 21072
rect 13872 21060 13878 21072
rect 14366 21060 14372 21072
rect 13872 21032 13917 21060
rect 14327 21032 14372 21060
rect 13872 21020 13878 21032
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 15654 21020 15660 21072
rect 15712 21060 15718 21072
rect 16040 21069 16068 21100
rect 17402 21088 17408 21140
rect 17460 21128 17466 21140
rect 17460 21100 17632 21128
rect 17460 21088 17466 21100
rect 15933 21063 15991 21069
rect 15933 21060 15945 21063
rect 15712 21032 15945 21060
rect 15712 21020 15718 21032
rect 15933 21029 15945 21032
rect 15979 21029 15991 21063
rect 15933 21023 15991 21029
rect 16025 21063 16083 21069
rect 16025 21029 16037 21063
rect 16071 21029 16083 21063
rect 17494 21060 17500 21072
rect 17455 21032 17500 21060
rect 16025 21023 16083 21029
rect 17494 21020 17500 21032
rect 17552 21020 17558 21072
rect 17604 21069 17632 21100
rect 17589 21063 17647 21069
rect 17589 21029 17601 21063
rect 17635 21029 17647 21063
rect 17589 21023 17647 21029
rect 12066 20992 12072 21004
rect 12027 20964 12072 20992
rect 12066 20952 12072 20964
rect 12124 20952 12130 21004
rect 12526 20992 12532 21004
rect 12487 20964 12532 20992
rect 12526 20952 12532 20964
rect 12584 20952 12590 21004
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 10505 20927 10563 20933
rect 10505 20924 10517 20927
rect 9732 20896 10517 20924
rect 9732 20884 9738 20896
rect 10505 20893 10517 20896
rect 10551 20924 10563 20927
rect 10778 20924 10784 20936
rect 10551 20896 10784 20924
rect 10551 20893 10563 20896
rect 10505 20887 10563 20893
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 12805 20927 12863 20933
rect 12805 20893 12817 20927
rect 12851 20924 12863 20927
rect 13262 20924 13268 20936
rect 12851 20896 13268 20924
rect 12851 20893 12863 20896
rect 12805 20887 12863 20893
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 16390 20924 16396 20936
rect 16351 20896 16396 20924
rect 16390 20884 16396 20896
rect 16448 20884 16454 20936
rect 17773 20927 17831 20933
rect 17773 20893 17785 20927
rect 17819 20893 17831 20927
rect 17773 20887 17831 20893
rect 10594 20856 10600 20868
rect 9600 20828 10600 20856
rect 10594 20816 10600 20828
rect 10652 20856 10658 20868
rect 11057 20859 11115 20865
rect 11057 20856 11069 20859
rect 10652 20828 11069 20856
rect 10652 20816 10658 20828
rect 11057 20825 11069 20828
rect 11103 20825 11115 20859
rect 11057 20819 11115 20825
rect 15749 20859 15807 20865
rect 15749 20825 15761 20859
rect 15795 20856 15807 20859
rect 16482 20856 16488 20868
rect 15795 20828 16488 20856
rect 15795 20825 15807 20828
rect 15749 20819 15807 20825
rect 16482 20816 16488 20828
rect 16540 20856 16546 20868
rect 17788 20856 17816 20887
rect 16540 20828 17816 20856
rect 16540 20816 16546 20828
rect 7650 20788 7656 20800
rect 6328 20760 6500 20788
rect 7611 20760 7656 20788
rect 6328 20748 6334 20760
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 9030 20788 9036 20800
rect 8991 20760 9036 20788
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 10134 20788 10140 20800
rect 10095 20760 10140 20788
rect 10134 20748 10140 20760
rect 10192 20748 10198 20800
rect 16298 20748 16304 20800
rect 16356 20788 16362 20800
rect 16853 20791 16911 20797
rect 16853 20788 16865 20791
rect 16356 20760 16865 20788
rect 16356 20748 16362 20760
rect 16853 20757 16865 20760
rect 16899 20757 16911 20791
rect 16853 20751 16911 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 3329 20587 3387 20593
rect 3329 20553 3341 20587
rect 3375 20584 3387 20587
rect 5534 20584 5540 20596
rect 3375 20556 5540 20584
rect 3375 20553 3387 20556
rect 3329 20547 3387 20553
rect 1854 20408 1860 20460
rect 1912 20448 1918 20460
rect 1912 20420 2774 20448
rect 1912 20408 1918 20420
rect 1740 20383 1798 20389
rect 1740 20349 1752 20383
rect 1786 20380 1798 20383
rect 1786 20352 2268 20380
rect 1786 20349 1798 20352
rect 1740 20343 1798 20349
rect 1394 20204 1400 20256
rect 1452 20244 1458 20256
rect 2240 20253 2268 20352
rect 2746 20312 2774 20420
rect 2844 20383 2902 20389
rect 2844 20349 2856 20383
rect 2890 20380 2902 20383
rect 3344 20380 3372 20547
rect 5534 20544 5540 20556
rect 5592 20544 5598 20596
rect 7742 20584 7748 20596
rect 7703 20556 7748 20584
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 8478 20584 8484 20596
rect 8439 20556 8484 20584
rect 8478 20544 8484 20556
rect 8536 20544 8542 20596
rect 9674 20584 9680 20596
rect 9635 20556 9680 20584
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 9950 20584 9956 20596
rect 9911 20556 9956 20584
rect 9950 20544 9956 20556
rect 10008 20584 10014 20596
rect 11146 20584 11152 20596
rect 10008 20556 10272 20584
rect 11107 20556 11152 20584
rect 10008 20544 10014 20556
rect 3970 20476 3976 20528
rect 4028 20516 4034 20528
rect 4430 20516 4436 20528
rect 4028 20488 4436 20516
rect 4028 20476 4034 20488
rect 4430 20476 4436 20488
rect 4488 20516 4494 20528
rect 4617 20519 4675 20525
rect 4617 20516 4629 20519
rect 4488 20488 4629 20516
rect 4488 20476 4494 20488
rect 4617 20485 4629 20488
rect 4663 20485 4675 20519
rect 4617 20479 4675 20485
rect 4890 20476 4896 20528
rect 4948 20516 4954 20528
rect 8938 20516 8944 20528
rect 4948 20488 8944 20516
rect 4948 20476 4954 20488
rect 8938 20476 8944 20488
rect 8996 20476 9002 20528
rect 8665 20451 8723 20457
rect 8665 20417 8677 20451
rect 8711 20448 8723 20451
rect 9030 20448 9036 20460
rect 8711 20420 9036 20448
rect 8711 20417 8723 20420
rect 8665 20411 8723 20417
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 10244 20457 10272 20556
rect 11146 20544 11152 20556
rect 11204 20544 11210 20596
rect 12066 20584 12072 20596
rect 12027 20556 12072 20584
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 12526 20544 12532 20596
rect 12584 20584 12590 20596
rect 12621 20587 12679 20593
rect 12621 20584 12633 20587
rect 12584 20556 12633 20584
rect 12584 20544 12590 20556
rect 12621 20553 12633 20556
rect 12667 20553 12679 20587
rect 14182 20584 14188 20596
rect 14143 20556 14188 20584
rect 12621 20547 12679 20553
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 15654 20544 15660 20596
rect 15712 20584 15718 20596
rect 15841 20587 15899 20593
rect 15841 20584 15853 20587
rect 15712 20556 15853 20584
rect 15712 20544 15718 20556
rect 15841 20553 15853 20556
rect 15887 20553 15899 20587
rect 15841 20547 15899 20553
rect 16022 20544 16028 20596
rect 16080 20584 16086 20596
rect 17402 20584 17408 20596
rect 16080 20556 17408 20584
rect 16080 20544 16086 20556
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 17494 20544 17500 20596
rect 17552 20584 17558 20596
rect 17773 20587 17831 20593
rect 17773 20584 17785 20587
rect 17552 20556 17785 20584
rect 17552 20544 17558 20556
rect 17773 20553 17785 20556
rect 17819 20553 17831 20587
rect 17773 20547 17831 20553
rect 16942 20476 16948 20528
rect 17000 20516 17006 20528
rect 18187 20519 18245 20525
rect 18187 20516 18199 20519
rect 17000 20488 18199 20516
rect 17000 20476 17006 20488
rect 18187 20485 18199 20488
rect 18233 20485 18245 20519
rect 18187 20479 18245 20485
rect 10229 20451 10287 20457
rect 9180 20420 9225 20448
rect 9180 20408 9186 20420
rect 10229 20417 10241 20451
rect 10275 20417 10287 20451
rect 10594 20448 10600 20460
rect 10555 20420 10600 20448
rect 10229 20411 10287 20417
rect 10594 20408 10600 20420
rect 10652 20448 10658 20460
rect 10870 20448 10876 20460
rect 10652 20420 10876 20448
rect 10652 20408 10658 20420
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 13262 20448 13268 20460
rect 13223 20420 13268 20448
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20448 16267 20451
rect 16482 20448 16488 20460
rect 16255 20420 16488 20448
rect 16255 20417 16267 20420
rect 16209 20411 16267 20417
rect 16482 20408 16488 20420
rect 16540 20408 16546 20460
rect 16850 20448 16856 20460
rect 16811 20420 16856 20448
rect 16850 20408 16856 20420
rect 16908 20408 16914 20460
rect 18506 20448 18512 20460
rect 18131 20420 18512 20448
rect 2890 20352 3372 20380
rect 3824 20383 3882 20389
rect 2890 20349 2902 20352
rect 2844 20343 2902 20349
rect 3824 20349 3836 20383
rect 3870 20349 3882 20383
rect 4249 20383 4307 20389
rect 4249 20380 4261 20383
rect 3824 20343 3882 20349
rect 4080 20352 4261 20380
rect 3839 20312 3867 20343
rect 4080 20312 4108 20352
rect 4249 20349 4261 20352
rect 4295 20349 4307 20383
rect 5074 20380 5080 20392
rect 4987 20352 5080 20380
rect 4249 20343 4307 20349
rect 5074 20340 5080 20352
rect 5132 20380 5138 20392
rect 5169 20383 5227 20389
rect 5169 20380 5181 20383
rect 5132 20352 5181 20380
rect 5132 20340 5138 20352
rect 5169 20349 5181 20352
rect 5215 20349 5227 20383
rect 5169 20343 5227 20349
rect 5258 20340 5264 20392
rect 5316 20380 5322 20392
rect 5629 20383 5687 20389
rect 5629 20380 5641 20383
rect 5316 20352 5641 20380
rect 5316 20340 5322 20352
rect 5629 20349 5641 20352
rect 5675 20349 5687 20383
rect 5629 20343 5687 20349
rect 6086 20340 6092 20392
rect 6144 20380 6150 20392
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6144 20352 6837 20380
rect 6144 20340 6150 20352
rect 6825 20349 6837 20352
rect 6871 20380 6883 20383
rect 7650 20380 7656 20392
rect 6871 20352 7656 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 7650 20340 7656 20352
rect 7708 20340 7714 20392
rect 14550 20340 14556 20392
rect 14608 20380 14614 20392
rect 15080 20383 15138 20389
rect 15080 20380 15092 20383
rect 14608 20352 15092 20380
rect 14608 20340 14614 20352
rect 15080 20349 15092 20352
rect 15126 20380 15138 20383
rect 15562 20380 15568 20392
rect 15126 20352 15568 20380
rect 15126 20349 15138 20352
rect 15080 20343 15138 20349
rect 15562 20340 15568 20352
rect 15620 20340 15626 20392
rect 18131 20389 18159 20420
rect 18506 20408 18512 20420
rect 18564 20448 18570 20460
rect 18601 20451 18659 20457
rect 18601 20448 18613 20451
rect 18564 20420 18613 20448
rect 18564 20408 18570 20420
rect 18601 20417 18613 20420
rect 18647 20448 18659 20451
rect 20346 20448 20352 20460
rect 18647 20420 20352 20448
rect 18647 20417 18659 20420
rect 18601 20411 18659 20417
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 18116 20383 18174 20389
rect 18116 20349 18128 20383
rect 18162 20349 18174 20383
rect 18116 20343 18174 20349
rect 19112 20383 19170 20389
rect 19112 20349 19124 20383
rect 19158 20380 19170 20383
rect 19518 20380 19524 20392
rect 19158 20352 19524 20380
rect 19158 20349 19170 20352
rect 19112 20343 19170 20349
rect 19518 20340 19524 20352
rect 19576 20340 19582 20392
rect 2746 20284 4108 20312
rect 5905 20315 5963 20321
rect 5905 20281 5917 20315
rect 5951 20312 5963 20315
rect 7006 20312 7012 20324
rect 5951 20284 7012 20312
rect 5951 20281 5963 20284
rect 5905 20275 5963 20281
rect 7006 20272 7012 20284
rect 7064 20272 7070 20324
rect 7187 20315 7245 20321
rect 7187 20281 7199 20315
rect 7233 20281 7245 20315
rect 7187 20275 7245 20281
rect 8757 20315 8815 20321
rect 8757 20281 8769 20315
rect 8803 20312 8815 20315
rect 9122 20312 9128 20324
rect 8803 20284 9128 20312
rect 8803 20281 8815 20284
rect 8757 20275 8815 20281
rect 1811 20247 1869 20253
rect 1811 20244 1823 20247
rect 1452 20216 1823 20244
rect 1452 20204 1458 20216
rect 1811 20213 1823 20216
rect 1857 20213 1869 20247
rect 1811 20207 1869 20213
rect 2225 20247 2283 20253
rect 2225 20213 2237 20247
rect 2271 20244 2283 20247
rect 2498 20244 2504 20256
rect 2271 20216 2504 20244
rect 2271 20213 2283 20216
rect 2225 20207 2283 20213
rect 2498 20204 2504 20216
rect 2556 20204 2562 20256
rect 2915 20247 2973 20253
rect 2915 20213 2927 20247
rect 2961 20244 2973 20247
rect 3510 20244 3516 20256
rect 2961 20216 3516 20244
rect 2961 20213 2973 20216
rect 2915 20207 2973 20213
rect 3510 20204 3516 20216
rect 3568 20204 3574 20256
rect 3786 20204 3792 20256
rect 3844 20244 3850 20256
rect 3927 20247 3985 20253
rect 3927 20244 3939 20247
rect 3844 20216 3939 20244
rect 3844 20204 3850 20216
rect 3927 20213 3939 20216
rect 3973 20213 3985 20247
rect 6178 20244 6184 20256
rect 6139 20216 6184 20244
rect 3927 20207 3985 20213
rect 6178 20204 6184 20216
rect 6236 20204 6242 20256
rect 6546 20244 6552 20256
rect 6507 20216 6552 20244
rect 6546 20204 6552 20216
rect 6604 20244 6610 20256
rect 7202 20244 7230 20275
rect 9122 20272 9128 20284
rect 9180 20272 9186 20324
rect 10321 20315 10379 20321
rect 10321 20281 10333 20315
rect 10367 20281 10379 20315
rect 10321 20275 10379 20281
rect 13586 20315 13644 20321
rect 13586 20281 13598 20315
rect 13632 20281 13644 20315
rect 13586 20275 13644 20281
rect 8021 20247 8079 20253
rect 8021 20244 8033 20247
rect 6604 20216 8033 20244
rect 6604 20204 6610 20216
rect 8021 20213 8033 20216
rect 8067 20213 8079 20247
rect 8021 20207 8079 20213
rect 10134 20204 10140 20256
rect 10192 20244 10198 20256
rect 10336 20244 10364 20275
rect 13170 20244 13176 20256
rect 10192 20216 10364 20244
rect 13131 20216 13176 20244
rect 10192 20204 10198 20216
rect 13170 20204 13176 20216
rect 13228 20244 13234 20256
rect 13601 20244 13629 20275
rect 16298 20272 16304 20324
rect 16356 20312 16362 20324
rect 19199 20315 19257 20321
rect 19199 20312 19211 20315
rect 16356 20284 16401 20312
rect 18064 20284 19211 20312
rect 16356 20272 16362 20284
rect 18064 20256 18092 20284
rect 19199 20281 19211 20284
rect 19245 20281 19257 20315
rect 19199 20275 19257 20281
rect 14458 20244 14464 20256
rect 13228 20216 13629 20244
rect 14419 20216 14464 20244
rect 13228 20204 13234 20216
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 15151 20247 15209 20253
rect 15151 20213 15163 20247
rect 15197 20244 15209 20247
rect 15378 20244 15384 20256
rect 15197 20216 15384 20244
rect 15197 20213 15209 20216
rect 15151 20207 15209 20213
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 15562 20244 15568 20256
rect 15523 20216 15568 20244
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 18046 20204 18052 20256
rect 18104 20204 18110 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 6822 20000 6828 20052
rect 6880 20040 6886 20052
rect 7285 20043 7343 20049
rect 7285 20040 7297 20043
rect 6880 20012 7297 20040
rect 6880 20000 6886 20012
rect 7285 20009 7297 20012
rect 7331 20009 7343 20043
rect 7285 20003 7343 20009
rect 8711 20043 8769 20049
rect 8711 20009 8723 20043
rect 8757 20040 8769 20043
rect 9030 20040 9036 20052
rect 8757 20012 9036 20040
rect 8757 20009 8769 20012
rect 8711 20003 8769 20009
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 9122 20000 9128 20052
rect 9180 20040 9186 20052
rect 9858 20040 9864 20052
rect 9180 20012 9864 20040
rect 9180 20000 9186 20012
rect 9858 20000 9864 20012
rect 9916 20040 9922 20052
rect 10597 20043 10655 20049
rect 10597 20040 10609 20043
rect 9916 20012 10609 20040
rect 9916 20000 9922 20012
rect 10597 20009 10609 20012
rect 10643 20009 10655 20043
rect 10597 20003 10655 20009
rect 10778 20000 10784 20052
rect 10836 20040 10842 20052
rect 11563 20043 11621 20049
rect 11563 20040 11575 20043
rect 10836 20012 11575 20040
rect 10836 20000 10842 20012
rect 11563 20009 11575 20012
rect 11609 20009 11621 20043
rect 11563 20003 11621 20009
rect 13170 20000 13176 20052
rect 13228 20040 13234 20052
rect 13265 20043 13323 20049
rect 13265 20040 13277 20043
rect 13228 20012 13277 20040
rect 13228 20000 13234 20012
rect 13265 20009 13277 20012
rect 13311 20009 13323 20043
rect 13265 20003 13323 20009
rect 13722 20000 13728 20052
rect 13780 20040 13786 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 13780 20012 14105 20040
rect 13780 20000 13786 20012
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 15838 20040 15844 20052
rect 15799 20012 15844 20040
rect 14093 20003 14151 20009
rect 15838 20000 15844 20012
rect 15896 20000 15902 20052
rect 16040 20012 17816 20040
rect 5537 19975 5595 19981
rect 5537 19941 5549 19975
rect 5583 19972 5595 19975
rect 6270 19972 6276 19984
rect 5583 19944 6276 19972
rect 5583 19941 5595 19944
rect 5537 19935 5595 19941
rect 6270 19932 6276 19944
rect 6328 19932 6334 19984
rect 6546 19932 6552 19984
rect 6604 19972 6610 19984
rect 6686 19975 6744 19981
rect 6686 19972 6698 19975
rect 6604 19944 6698 19972
rect 6604 19932 6610 19944
rect 6686 19941 6698 19944
rect 6732 19941 6744 19975
rect 6686 19935 6744 19941
rect 9582 19932 9588 19984
rect 9640 19972 9646 19984
rect 9998 19975 10056 19981
rect 9998 19972 10010 19975
rect 9640 19944 10010 19972
rect 9640 19932 9646 19944
rect 9998 19941 10010 19944
rect 10044 19941 10056 19975
rect 9998 19935 10056 19941
rect 15746 19932 15752 19984
rect 15804 19972 15810 19984
rect 16040 19972 16068 20012
rect 17788 19984 17816 20012
rect 16206 19972 16212 19984
rect 15804 19944 16068 19972
rect 16167 19944 16212 19972
rect 15804 19932 15810 19944
rect 16206 19932 16212 19944
rect 16264 19932 16270 19984
rect 16761 19975 16819 19981
rect 16761 19941 16773 19975
rect 16807 19972 16819 19975
rect 16850 19972 16856 19984
rect 16807 19944 16856 19972
rect 16807 19941 16819 19944
rect 16761 19935 16819 19941
rect 16850 19932 16856 19944
rect 16908 19932 16914 19984
rect 17770 19972 17776 19984
rect 17683 19944 17776 19972
rect 17770 19932 17776 19944
rect 17828 19932 17834 19984
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 1486 19904 1492 19916
rect 1443 19876 1492 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 1486 19864 1492 19876
rect 1544 19864 1550 19916
rect 2682 19864 2688 19916
rect 2740 19904 2746 19916
rect 2961 19907 3019 19913
rect 2961 19904 2973 19907
rect 2740 19876 2973 19904
rect 2740 19864 2746 19876
rect 2961 19873 2973 19876
rect 3007 19904 3019 19907
rect 4614 19904 4620 19916
rect 3007 19876 4620 19904
rect 3007 19873 3019 19876
rect 2961 19867 3019 19873
rect 4614 19864 4620 19876
rect 4672 19864 4678 19916
rect 5077 19907 5135 19913
rect 5077 19873 5089 19907
rect 5123 19873 5135 19907
rect 5258 19904 5264 19916
rect 5219 19876 5264 19904
rect 5077 19867 5135 19873
rect 4706 19796 4712 19848
rect 4764 19836 4770 19848
rect 5092 19836 5120 19867
rect 5258 19864 5264 19876
rect 5316 19904 5322 19916
rect 5442 19904 5448 19916
rect 5316 19876 5448 19904
rect 5316 19864 5322 19876
rect 5442 19864 5448 19876
rect 5500 19904 5506 19916
rect 5813 19907 5871 19913
rect 5813 19904 5825 19907
rect 5500 19876 5825 19904
rect 5500 19864 5506 19876
rect 5813 19873 5825 19876
rect 5859 19873 5871 19907
rect 5813 19867 5871 19873
rect 8640 19907 8698 19913
rect 8640 19873 8652 19907
rect 8686 19904 8698 19907
rect 8938 19904 8944 19916
rect 8686 19876 8944 19904
rect 8686 19873 8698 19876
rect 8640 19867 8698 19873
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 11492 19907 11550 19913
rect 11492 19873 11504 19907
rect 11538 19904 11550 19907
rect 11882 19904 11888 19916
rect 11538 19876 11888 19904
rect 11538 19873 11550 19876
rect 11492 19867 11550 19873
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 13814 19864 13820 19916
rect 13872 19904 13878 19916
rect 14458 19904 14464 19916
rect 13872 19876 14464 19904
rect 13872 19864 13878 19876
rect 14458 19864 14464 19876
rect 14516 19864 14522 19916
rect 18874 19864 18880 19916
rect 18932 19904 18938 19916
rect 19188 19907 19246 19913
rect 19188 19904 19200 19907
rect 18932 19876 19200 19904
rect 18932 19864 18938 19876
rect 19188 19873 19200 19876
rect 19234 19873 19246 19907
rect 19188 19867 19246 19873
rect 6362 19836 6368 19848
rect 4764 19808 6040 19836
rect 6323 19808 6368 19836
rect 4764 19796 4770 19808
rect 6012 19768 6040 19808
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 7006 19796 7012 19848
rect 7064 19836 7070 19848
rect 9677 19839 9735 19845
rect 9677 19836 9689 19839
rect 7064 19808 9689 19836
rect 7064 19796 7070 19808
rect 9677 19805 9689 19808
rect 9723 19836 9735 19839
rect 10594 19836 10600 19848
rect 9723 19808 10600 19836
rect 9723 19805 9735 19808
rect 9677 19799 9735 19805
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 12802 19796 12808 19848
rect 12860 19836 12866 19848
rect 12897 19839 12955 19845
rect 12897 19836 12909 19839
rect 12860 19808 12909 19836
rect 12860 19796 12866 19808
rect 12897 19805 12909 19808
rect 12943 19805 12955 19839
rect 12897 19799 12955 19805
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19836 16175 19839
rect 16390 19836 16396 19848
rect 16163 19808 16396 19836
rect 16163 19805 16175 19808
rect 16117 19799 16175 19805
rect 16390 19796 16396 19808
rect 16448 19796 16454 19848
rect 17678 19836 17684 19848
rect 17639 19808 17684 19836
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 17954 19836 17960 19848
rect 17915 19808 17960 19836
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 12066 19768 12072 19780
rect 6012 19740 12072 19768
rect 12066 19728 12072 19740
rect 12124 19728 12130 19780
rect 1535 19703 1593 19709
rect 1535 19669 1547 19703
rect 1581 19700 1593 19703
rect 1670 19700 1676 19712
rect 1581 19672 1676 19700
rect 1581 19669 1593 19672
rect 1535 19663 1593 19669
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 2406 19660 2412 19712
rect 2464 19700 2470 19712
rect 3145 19703 3203 19709
rect 3145 19700 3157 19703
rect 2464 19672 3157 19700
rect 2464 19660 2470 19672
rect 3145 19669 3157 19672
rect 3191 19669 3203 19703
rect 7742 19700 7748 19712
rect 7703 19672 7748 19700
rect 3145 19663 3203 19669
rect 7742 19660 7748 19672
rect 7800 19660 7806 19712
rect 12526 19700 12532 19712
rect 12487 19672 12532 19700
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 19291 19703 19349 19709
rect 19291 19700 19303 19703
rect 16632 19672 19303 19700
rect 16632 19660 16638 19672
rect 19291 19669 19303 19672
rect 19337 19669 19349 19703
rect 19291 19663 19349 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 4706 19496 4712 19508
rect 4667 19468 4712 19496
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 10134 19456 10140 19508
rect 10192 19496 10198 19508
rect 10413 19499 10471 19505
rect 10413 19496 10425 19499
rect 10192 19468 10425 19496
rect 10192 19456 10198 19468
rect 10413 19465 10425 19468
rect 10459 19465 10471 19499
rect 10413 19459 10471 19465
rect 10594 19456 10600 19508
rect 10652 19496 10658 19508
rect 10689 19499 10747 19505
rect 10689 19496 10701 19499
rect 10652 19468 10701 19496
rect 10652 19456 10658 19468
rect 10689 19465 10701 19468
rect 10735 19465 10747 19499
rect 10689 19459 10747 19465
rect 15841 19499 15899 19505
rect 15841 19465 15853 19499
rect 15887 19496 15899 19499
rect 16206 19496 16212 19508
rect 15887 19468 16212 19496
rect 15887 19465 15899 19468
rect 15841 19459 15899 19465
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 16390 19456 16396 19508
rect 16448 19496 16454 19508
rect 16577 19499 16635 19505
rect 16577 19496 16589 19499
rect 16448 19468 16589 19496
rect 16448 19456 16454 19468
rect 16577 19465 16589 19468
rect 16623 19496 16635 19499
rect 17954 19496 17960 19508
rect 16623 19468 17960 19496
rect 16623 19465 16635 19468
rect 16577 19459 16635 19465
rect 17954 19456 17960 19468
rect 18012 19456 18018 19508
rect 24762 19496 24768 19508
rect 18064 19468 19334 19496
rect 24723 19468 24768 19496
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 8665 19431 8723 19437
rect 8665 19428 8677 19431
rect 8628 19400 8677 19428
rect 8628 19388 8634 19400
rect 8665 19397 8677 19400
rect 8711 19397 8723 19431
rect 8665 19391 8723 19397
rect 5905 19363 5963 19369
rect 5905 19329 5917 19363
rect 5951 19360 5963 19363
rect 6362 19360 6368 19372
rect 5951 19332 6368 19360
rect 5951 19329 5963 19332
rect 5905 19323 5963 19329
rect 6362 19320 6368 19332
rect 6420 19360 6426 19372
rect 7009 19363 7067 19369
rect 7009 19360 7021 19363
rect 6420 19332 7021 19360
rect 6420 19320 6426 19332
rect 7009 19329 7021 19332
rect 7055 19329 7067 19363
rect 8680 19360 8708 19391
rect 11330 19388 11336 19440
rect 11388 19428 11394 19440
rect 11517 19431 11575 19437
rect 11517 19428 11529 19431
rect 11388 19400 11529 19428
rect 11388 19388 11394 19400
rect 11517 19397 11529 19400
rect 11563 19428 11575 19431
rect 12434 19428 12440 19440
rect 11563 19400 12440 19428
rect 11563 19397 11575 19400
rect 11517 19391 11575 19397
rect 12434 19388 12440 19400
rect 12492 19388 12498 19440
rect 17681 19431 17739 19437
rect 17681 19397 17693 19431
rect 17727 19428 17739 19431
rect 17770 19428 17776 19440
rect 17727 19400 17776 19428
rect 17727 19397 17739 19400
rect 17681 19391 17739 19397
rect 17770 19388 17776 19400
rect 17828 19388 17834 19440
rect 10134 19360 10140 19372
rect 8680 19332 10140 19360
rect 7009 19323 7067 19329
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 10238 19332 12173 19360
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19261 1455 19295
rect 1397 19255 1455 19261
rect 2660 19295 2718 19301
rect 2660 19261 2672 19295
rect 2706 19292 2718 19295
rect 2706 19264 3188 19292
rect 2706 19261 2718 19264
rect 2660 19255 2718 19261
rect 1412 19224 1440 19255
rect 2038 19224 2044 19236
rect 1412 19196 2044 19224
rect 2038 19184 2044 19196
rect 2096 19184 2102 19236
rect 3160 19233 3188 19264
rect 3418 19252 3424 19304
rect 3476 19292 3482 19304
rect 3605 19295 3663 19301
rect 3605 19292 3617 19295
rect 3476 19264 3617 19292
rect 3476 19252 3482 19264
rect 3605 19261 3617 19264
rect 3651 19261 3663 19295
rect 4062 19292 4068 19304
rect 4023 19264 4068 19292
rect 3605 19255 3663 19261
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5258 19292 5264 19304
rect 5123 19264 5264 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 5442 19252 5448 19304
rect 5500 19292 5506 19304
rect 5629 19295 5687 19301
rect 5629 19292 5641 19295
rect 5500 19264 5641 19292
rect 5500 19252 5506 19264
rect 5629 19261 5641 19264
rect 5675 19261 5687 19295
rect 7742 19292 7748 19304
rect 7703 19264 7748 19292
rect 5629 19255 5687 19261
rect 7742 19252 7748 19264
rect 7800 19252 7806 19304
rect 9398 19292 9404 19304
rect 7944 19264 9404 19292
rect 3145 19227 3203 19233
rect 3145 19193 3157 19227
rect 3191 19224 3203 19227
rect 4246 19224 4252 19236
rect 3191 19196 4252 19224
rect 3191 19193 3203 19196
rect 3145 19187 3203 19193
rect 4246 19184 4252 19196
rect 4304 19184 4310 19236
rect 4341 19227 4399 19233
rect 4341 19193 4353 19227
rect 4387 19224 4399 19227
rect 7944 19224 7972 19264
rect 9398 19252 9404 19264
rect 9456 19292 9462 19304
rect 9493 19295 9551 19301
rect 9493 19292 9505 19295
rect 9456 19264 9505 19292
rect 9456 19252 9462 19264
rect 9493 19261 9505 19264
rect 9539 19261 9551 19295
rect 10238 19292 10266 19332
rect 12161 19329 12173 19332
rect 12207 19329 12219 19363
rect 12161 19323 12219 19329
rect 11333 19295 11391 19301
rect 11333 19292 11345 19295
rect 9493 19255 9551 19261
rect 10152 19264 10266 19292
rect 11164 19264 11345 19292
rect 8938 19224 8944 19236
rect 4387 19196 7972 19224
rect 8899 19196 8944 19224
rect 4387 19193 4399 19196
rect 4341 19187 4399 19193
rect 8938 19184 8944 19196
rect 8996 19184 9002 19236
rect 9814 19227 9872 19233
rect 9814 19224 9826 19227
rect 9600 19196 9826 19224
rect 9600 19168 9628 19196
rect 9814 19193 9826 19196
rect 9860 19224 9872 19227
rect 10152 19224 10180 19264
rect 9860 19196 10180 19224
rect 9860 19193 9872 19196
rect 9814 19187 9872 19193
rect 11164 19168 11192 19264
rect 11333 19261 11345 19264
rect 11379 19261 11391 19295
rect 11333 19255 11391 19261
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2590 19156 2596 19168
rect 2547 19128 2596 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 2731 19159 2789 19165
rect 2731 19125 2743 19159
rect 2777 19156 2789 19159
rect 3234 19156 3240 19168
rect 2777 19128 3240 19156
rect 2777 19125 2789 19128
rect 2731 19119 2789 19125
rect 3234 19116 3240 19128
rect 3292 19116 3298 19168
rect 3418 19156 3424 19168
rect 3379 19128 3424 19156
rect 3418 19116 3424 19128
rect 3476 19116 3482 19168
rect 6362 19156 6368 19168
rect 6323 19128 6368 19156
rect 6362 19116 6368 19128
rect 6420 19156 6426 19168
rect 6546 19156 6552 19168
rect 6420 19128 6552 19156
rect 6420 19116 6426 19128
rect 6546 19116 6552 19128
rect 6604 19156 6610 19168
rect 7561 19159 7619 19165
rect 7561 19156 7573 19159
rect 6604 19128 7573 19156
rect 6604 19116 6610 19128
rect 7561 19125 7573 19128
rect 7607 19156 7619 19159
rect 7926 19156 7932 19168
rect 7607 19128 7932 19156
rect 7607 19125 7619 19128
rect 7561 19119 7619 19125
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 8018 19116 8024 19168
rect 8076 19156 8082 19168
rect 8113 19159 8171 19165
rect 8113 19156 8125 19159
rect 8076 19128 8125 19156
rect 8076 19116 8082 19128
rect 8113 19125 8125 19128
rect 8159 19125 8171 19159
rect 8113 19119 8171 19125
rect 9401 19159 9459 19165
rect 9401 19125 9413 19159
rect 9447 19156 9459 19159
rect 9582 19156 9588 19168
rect 9447 19128 9588 19156
rect 9447 19125 9459 19128
rect 9401 19119 9459 19125
rect 9582 19116 9588 19128
rect 9640 19116 9646 19168
rect 11146 19156 11152 19168
rect 11107 19128 11152 19156
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 11882 19156 11888 19168
rect 11843 19128 11888 19156
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12176 19156 12204 19323
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 18064 19360 18092 19468
rect 13872 19332 18092 19360
rect 19306 19360 19334 19468
rect 24762 19456 24768 19468
rect 24820 19456 24826 19508
rect 20073 19363 20131 19369
rect 20073 19360 20085 19363
rect 19306 19332 20085 19360
rect 13872 19320 13878 19332
rect 20073 19329 20085 19332
rect 20119 19329 20131 19363
rect 20073 19323 20131 19329
rect 12526 19292 12532 19304
rect 12487 19264 12532 19292
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 12802 19252 12808 19304
rect 12860 19292 12866 19304
rect 13262 19292 13268 19304
rect 12860 19264 13268 19292
rect 12860 19252 12866 19264
rect 13262 19252 13268 19264
rect 13320 19252 13326 19304
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19292 13507 19295
rect 13906 19292 13912 19304
rect 13495 19264 13912 19292
rect 13495 19261 13507 19264
rect 13449 19255 13507 19261
rect 13906 19252 13912 19264
rect 13964 19252 13970 19304
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14792 19264 14933 19292
rect 14792 19252 14798 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 16720 19295 16778 19301
rect 16720 19261 16732 19295
rect 16766 19292 16778 19295
rect 17126 19292 17132 19304
rect 16766 19264 17132 19292
rect 16766 19261 16778 19264
rect 16720 19255 16778 19261
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 17310 19252 17316 19304
rect 17368 19292 17374 19304
rect 18084 19295 18142 19301
rect 18084 19292 18096 19295
rect 17368 19264 18096 19292
rect 17368 19252 17374 19264
rect 18084 19261 18096 19264
rect 18130 19292 18142 19295
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 18130 19264 18521 19292
rect 18130 19261 18142 19264
rect 18084 19255 18142 19261
rect 18509 19261 18521 19264
rect 18555 19292 18567 19295
rect 18966 19292 18972 19304
rect 18555 19264 18972 19292
rect 18555 19261 18567 19264
rect 18509 19255 18567 19261
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19087 19295 19145 19301
rect 19087 19261 19099 19295
rect 19133 19292 19145 19295
rect 19426 19292 19432 19304
rect 19133 19264 19432 19292
rect 19133 19261 19145 19264
rect 19087 19255 19145 19261
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 20530 19252 20536 19304
rect 20588 19292 20594 19304
rect 23106 19292 23112 19304
rect 20588 19264 23112 19292
rect 20588 19252 20594 19264
rect 23106 19252 23112 19264
rect 23164 19292 23170 19304
rect 24581 19295 24639 19301
rect 24581 19292 24593 19295
rect 23164 19264 24593 19292
rect 23164 19252 23170 19264
rect 24581 19261 24593 19264
rect 24627 19292 24639 19295
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 24627 19264 25145 19292
rect 24627 19261 24639 19264
rect 24581 19255 24639 19261
rect 25133 19261 25145 19264
rect 25179 19261 25191 19295
rect 25133 19255 25191 19261
rect 13170 19184 13176 19236
rect 13228 19224 13234 19236
rect 13817 19227 13875 19233
rect 13817 19224 13829 19227
rect 13228 19196 13829 19224
rect 13228 19184 13234 19196
rect 13817 19193 13829 19196
rect 13863 19224 13875 19227
rect 16807 19227 16865 19233
rect 13863 19196 14872 19224
rect 13863 19193 13875 19196
rect 13817 19187 13875 19193
rect 12897 19159 12955 19165
rect 12897 19156 12909 19159
rect 12176 19128 12909 19156
rect 12897 19125 12909 19128
rect 12943 19156 12955 19159
rect 13188 19156 13216 19184
rect 12943 19128 13216 19156
rect 12943 19125 12955 19128
rect 12897 19119 12955 19125
rect 13262 19116 13268 19168
rect 13320 19156 13326 19168
rect 14844 19165 14872 19196
rect 16807 19193 16819 19227
rect 16853 19224 16865 19227
rect 17678 19224 17684 19236
rect 16853 19196 17684 19224
rect 16853 19193 16865 19196
rect 16807 19187 16865 19193
rect 17678 19184 17684 19196
rect 17736 19184 17742 19236
rect 18874 19184 18880 19236
rect 18932 19224 18938 19236
rect 19521 19227 19579 19233
rect 19521 19224 19533 19227
rect 18932 19196 19533 19224
rect 18932 19184 18938 19196
rect 19521 19193 19533 19196
rect 19567 19193 19579 19227
rect 19521 19187 19579 19193
rect 14093 19159 14151 19165
rect 14093 19156 14105 19159
rect 13320 19128 14105 19156
rect 13320 19116 13326 19128
rect 14093 19125 14105 19128
rect 14139 19125 14151 19159
rect 14093 19119 14151 19125
rect 14829 19159 14887 19165
rect 14829 19125 14841 19159
rect 14875 19156 14887 19159
rect 15289 19159 15347 19165
rect 15289 19156 15301 19159
rect 14875 19128 15301 19156
rect 14875 19125 14887 19128
rect 14829 19119 14887 19125
rect 15289 19125 15301 19128
rect 15335 19125 15347 19159
rect 15289 19119 15347 19125
rect 17770 19116 17776 19168
rect 17828 19156 17834 19168
rect 18187 19159 18245 19165
rect 18187 19156 18199 19159
rect 17828 19128 18199 19156
rect 17828 19116 17834 19128
rect 18187 19125 18199 19128
rect 18233 19125 18245 19159
rect 18187 19119 18245 19125
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 19245 19159 19303 19165
rect 19245 19156 19257 19159
rect 19116 19128 19257 19156
rect 19116 19116 19122 19128
rect 19245 19125 19257 19128
rect 19291 19125 19303 19159
rect 19245 19119 19303 19125
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 19889 19159 19947 19165
rect 19889 19156 19901 19159
rect 19484 19128 19901 19156
rect 19484 19116 19490 19128
rect 19889 19125 19901 19128
rect 19935 19125 19947 19159
rect 19889 19119 19947 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 4246 18912 4252 18964
rect 4304 18952 4310 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 4304 18924 8493 18952
rect 4304 18912 4310 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 9398 18952 9404 18964
rect 9359 18924 9404 18952
rect 8481 18915 8539 18921
rect 9398 18912 9404 18924
rect 9456 18912 9462 18964
rect 12434 18952 12440 18964
rect 12395 18924 12440 18952
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 13170 18952 13176 18964
rect 13131 18924 13176 18952
rect 13170 18912 13176 18924
rect 13228 18912 13234 18964
rect 13538 18912 13544 18964
rect 13596 18952 13602 18964
rect 13725 18955 13783 18961
rect 13725 18952 13737 18955
rect 13596 18924 13737 18952
rect 13596 18912 13602 18924
rect 13725 18921 13737 18924
rect 13771 18921 13783 18955
rect 13725 18915 13783 18921
rect 16209 18955 16267 18961
rect 16209 18921 16221 18955
rect 16255 18952 16267 18955
rect 16298 18952 16304 18964
rect 16255 18924 16304 18952
rect 16255 18921 16267 18924
rect 16209 18915 16267 18921
rect 16298 18912 16304 18924
rect 16356 18912 16362 18964
rect 16574 18952 16580 18964
rect 16535 18924 16580 18952
rect 16574 18912 16580 18924
rect 16632 18912 16638 18964
rect 17126 18952 17132 18964
rect 17087 18924 17132 18952
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 18049 18955 18107 18961
rect 18049 18952 18061 18955
rect 17736 18924 18061 18952
rect 17736 18912 17742 18924
rect 18049 18921 18061 18924
rect 18095 18921 18107 18955
rect 18049 18915 18107 18921
rect 24210 18912 24216 18964
rect 24268 18952 24274 18964
rect 24765 18955 24823 18961
rect 24765 18952 24777 18955
rect 24268 18924 24777 18952
rect 24268 18912 24274 18924
rect 24765 18921 24777 18924
rect 24811 18921 24823 18955
rect 24765 18915 24823 18921
rect 4893 18887 4951 18893
rect 4893 18853 4905 18887
rect 4939 18884 4951 18887
rect 6086 18884 6092 18896
rect 4939 18856 5488 18884
rect 6047 18856 6092 18884
rect 4939 18853 4951 18856
rect 4893 18847 4951 18853
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 1946 18816 1952 18828
rect 1903 18788 1952 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 1946 18776 1952 18788
rect 2004 18816 2010 18828
rect 2958 18816 2964 18828
rect 3016 18825 3022 18828
rect 3016 18819 3054 18825
rect 2004 18788 2964 18816
rect 2004 18776 2010 18788
rect 2958 18776 2964 18788
rect 3042 18785 3054 18819
rect 3016 18779 3054 18785
rect 3016 18776 3022 18779
rect 3694 18708 3700 18760
rect 3752 18748 3758 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3752 18720 4077 18748
rect 3752 18708 3758 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 2087 18683 2145 18689
rect 2087 18649 2099 18683
rect 2133 18680 2145 18683
rect 4522 18680 4528 18692
rect 2133 18652 4528 18680
rect 2133 18649 2145 18652
rect 2087 18643 2145 18649
rect 4522 18640 4528 18652
rect 4580 18640 4586 18692
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 1581 18615 1639 18621
rect 1581 18612 1593 18615
rect 1544 18584 1593 18612
rect 1544 18572 1550 18584
rect 1581 18581 1593 18584
rect 1627 18581 1639 18615
rect 1581 18575 1639 18581
rect 3099 18615 3157 18621
rect 3099 18581 3111 18615
rect 3145 18612 3157 18615
rect 3602 18612 3608 18624
rect 3145 18584 3608 18612
rect 3145 18581 3157 18584
rect 3099 18575 3157 18581
rect 3602 18572 3608 18584
rect 3660 18572 3666 18624
rect 3697 18615 3755 18621
rect 3697 18581 3709 18615
rect 3743 18612 3755 18615
rect 4062 18612 4068 18624
rect 3743 18584 4068 18612
rect 3743 18581 3755 18584
rect 3697 18575 3755 18581
rect 4062 18572 4068 18584
rect 4120 18612 4126 18624
rect 4908 18612 4936 18847
rect 5460 18828 5488 18856
rect 6086 18844 6092 18856
rect 6144 18844 6150 18896
rect 10226 18844 10232 18896
rect 10284 18884 10290 18896
rect 10321 18887 10379 18893
rect 10321 18884 10333 18887
rect 10284 18856 10333 18884
rect 10284 18844 10290 18856
rect 10321 18853 10333 18856
rect 10367 18853 10379 18887
rect 10870 18884 10876 18896
rect 10831 18856 10876 18884
rect 10321 18847 10379 18853
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 15610 18887 15668 18893
rect 15610 18884 15622 18887
rect 15528 18856 15622 18884
rect 15528 18844 15534 18856
rect 15610 18853 15622 18856
rect 15656 18853 15668 18887
rect 15610 18847 15668 18853
rect 5350 18816 5356 18828
rect 5311 18788 5356 18816
rect 5350 18776 5356 18788
rect 5408 18776 5414 18828
rect 5442 18776 5448 18828
rect 5500 18816 5506 18828
rect 5813 18819 5871 18825
rect 5813 18816 5825 18819
rect 5500 18788 5825 18816
rect 5500 18776 5506 18788
rect 5813 18785 5825 18788
rect 5859 18785 5871 18819
rect 7006 18816 7012 18828
rect 6967 18788 7012 18816
rect 5813 18779 5871 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 7190 18776 7196 18828
rect 7248 18816 7254 18828
rect 7377 18819 7435 18825
rect 7377 18816 7389 18819
rect 7248 18788 7389 18816
rect 7248 18776 7254 18788
rect 7377 18785 7389 18788
rect 7423 18785 7435 18819
rect 7377 18779 7435 18785
rect 11701 18819 11759 18825
rect 11701 18785 11713 18819
rect 11747 18816 11759 18819
rect 11790 18816 11796 18828
rect 11747 18788 11796 18816
rect 11747 18785 11759 18788
rect 11701 18779 11759 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 11882 18776 11888 18828
rect 11940 18816 11946 18828
rect 17034 18816 17040 18828
rect 11940 18788 15654 18816
rect 16995 18788 17040 18816
rect 11940 18776 11946 18788
rect 7653 18751 7711 18757
rect 7653 18717 7665 18751
rect 7699 18748 7711 18751
rect 8018 18748 8024 18760
rect 7699 18720 8024 18748
rect 7699 18717 7711 18720
rect 7653 18711 7711 18717
rect 8018 18708 8024 18720
rect 8076 18708 8082 18760
rect 8481 18751 8539 18757
rect 8481 18717 8493 18751
rect 8527 18748 8539 18751
rect 8662 18748 8668 18760
rect 8527 18720 8668 18748
rect 8527 18717 8539 18720
rect 8481 18711 8539 18717
rect 8662 18708 8668 18720
rect 8720 18708 8726 18760
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18748 10287 18751
rect 12805 18751 12863 18757
rect 10275 18720 11284 18748
rect 10275 18717 10287 18720
rect 10229 18711 10287 18717
rect 5074 18640 5080 18692
rect 5132 18680 5138 18692
rect 9030 18680 9036 18692
rect 5132 18652 9036 18680
rect 5132 18640 5138 18652
rect 9030 18640 9036 18652
rect 9088 18640 9094 18692
rect 11256 18689 11284 18720
rect 12805 18717 12817 18751
rect 12851 18748 12863 18751
rect 13170 18748 13176 18760
rect 12851 18720 13176 18748
rect 12851 18717 12863 18720
rect 12805 18711 12863 18717
rect 13170 18708 13176 18720
rect 13228 18708 13234 18760
rect 15286 18748 15292 18760
rect 15247 18720 15292 18748
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 15626 18748 15654 18788
rect 17034 18776 17040 18788
rect 17092 18776 17098 18828
rect 17402 18776 17408 18828
rect 17460 18816 17466 18828
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 17460 18788 17509 18816
rect 17460 18776 17466 18788
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 18668 18819 18726 18825
rect 18668 18785 18680 18819
rect 18714 18816 18726 18819
rect 18782 18816 18788 18828
rect 18714 18788 18788 18816
rect 18714 18785 18726 18788
rect 18668 18779 18726 18785
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 18966 18776 18972 18828
rect 19024 18816 19030 18828
rect 19648 18819 19706 18825
rect 19648 18816 19660 18819
rect 19024 18788 19660 18816
rect 19024 18776 19030 18788
rect 19648 18785 19660 18788
rect 19694 18816 19706 18819
rect 20070 18816 20076 18828
rect 19694 18788 20076 18816
rect 19694 18785 19706 18788
rect 19648 18779 19706 18785
rect 20070 18776 20076 18788
rect 20128 18776 20134 18828
rect 24118 18776 24124 18828
rect 24176 18816 24182 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 24176 18788 24593 18816
rect 24176 18776 24182 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 18506 18748 18512 18760
rect 15626 18720 18512 18748
rect 18506 18708 18512 18720
rect 18564 18708 18570 18760
rect 20438 18708 20444 18760
rect 20496 18748 20502 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20496 18720 20913 18748
rect 20496 18708 20502 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 11241 18683 11299 18689
rect 11241 18649 11253 18683
rect 11287 18680 11299 18683
rect 17770 18680 17776 18692
rect 11287 18652 17776 18680
rect 11287 18649 11299 18652
rect 11241 18643 11299 18649
rect 17770 18640 17776 18652
rect 17828 18640 17834 18692
rect 18414 18640 18420 18692
rect 18472 18680 18478 18692
rect 19751 18683 19809 18689
rect 19751 18680 19763 18683
rect 18472 18652 19763 18680
rect 18472 18640 18478 18652
rect 19751 18649 19763 18652
rect 19797 18649 19809 18683
rect 19751 18643 19809 18649
rect 5258 18612 5264 18624
rect 4120 18584 4936 18612
rect 5219 18584 5264 18612
rect 4120 18572 4126 18584
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 8021 18615 8079 18621
rect 8021 18581 8033 18615
rect 8067 18612 8079 18615
rect 8294 18612 8300 18624
rect 8067 18584 8300 18612
rect 8067 18581 8079 18584
rect 8021 18575 8079 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 8711 18615 8769 18621
rect 8711 18581 8723 18615
rect 8757 18612 8769 18615
rect 9214 18612 9220 18624
rect 8757 18584 9220 18612
rect 8757 18581 8769 18584
rect 8711 18575 8769 18581
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 9582 18572 9588 18624
rect 9640 18612 9646 18624
rect 9861 18615 9919 18621
rect 9861 18612 9873 18615
rect 9640 18584 9873 18612
rect 9640 18572 9646 18584
rect 9861 18581 9873 18584
rect 9907 18581 9919 18615
rect 9861 18575 9919 18581
rect 11839 18615 11897 18621
rect 11839 18581 11851 18615
rect 11885 18612 11897 18615
rect 12158 18612 12164 18624
rect 11885 18584 12164 18612
rect 11885 18581 11897 18584
rect 11839 18575 11897 18581
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 14090 18612 14096 18624
rect 14051 18584 14096 18612
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 14734 18572 14740 18624
rect 14792 18612 14798 18624
rect 14921 18615 14979 18621
rect 14921 18612 14933 18615
rect 14792 18584 14933 18612
rect 14792 18572 14798 18584
rect 14921 18581 14933 18584
rect 14967 18581 14979 18615
rect 14921 18575 14979 18581
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 18739 18615 18797 18621
rect 18739 18612 18751 18615
rect 18656 18584 18751 18612
rect 18656 18572 18662 18584
rect 18739 18581 18751 18584
rect 18785 18581 18797 18615
rect 18739 18575 18797 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 2041 18411 2099 18417
rect 2041 18408 2053 18411
rect 2004 18380 2053 18408
rect 2004 18368 2010 18380
rect 2041 18377 2053 18380
rect 2087 18377 2099 18411
rect 2041 18371 2099 18377
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 4890 18408 4896 18420
rect 2547 18380 4896 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 1648 18207 1706 18213
rect 1648 18173 1660 18207
rect 1694 18204 1706 18207
rect 2516 18204 2544 18371
rect 4890 18368 4896 18380
rect 4948 18368 4954 18420
rect 5077 18411 5135 18417
rect 5077 18377 5089 18411
rect 5123 18408 5135 18411
rect 5166 18408 5172 18420
rect 5123 18380 5172 18408
rect 5123 18377 5135 18380
rect 5077 18371 5135 18377
rect 5166 18368 5172 18380
rect 5224 18408 5230 18420
rect 7006 18408 7012 18420
rect 5224 18380 7012 18408
rect 5224 18368 5230 18380
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 9030 18408 9036 18420
rect 8991 18380 9036 18408
rect 9030 18368 9036 18380
rect 9088 18408 9094 18420
rect 12069 18411 12127 18417
rect 12069 18408 12081 18411
rect 9088 18380 12081 18408
rect 9088 18368 9094 18380
rect 12069 18377 12081 18380
rect 12115 18408 12127 18411
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 12115 18380 12173 18408
rect 12115 18377 12127 18380
rect 12069 18371 12127 18377
rect 12161 18377 12173 18380
rect 12207 18377 12219 18411
rect 12161 18371 12219 18377
rect 13262 18368 13268 18420
rect 13320 18408 13326 18420
rect 13449 18411 13507 18417
rect 13449 18408 13461 18411
rect 13320 18380 13461 18408
rect 13320 18368 13326 18380
rect 13449 18377 13461 18380
rect 13495 18377 13507 18411
rect 13449 18371 13507 18377
rect 13906 18368 13912 18420
rect 13964 18408 13970 18420
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 13964 18380 15761 18408
rect 13964 18368 13970 18380
rect 15749 18377 15761 18380
rect 15795 18408 15807 18411
rect 17034 18408 17040 18420
rect 15795 18380 15884 18408
rect 16995 18380 17040 18408
rect 15795 18377 15807 18380
rect 15749 18371 15807 18377
rect 2958 18300 2964 18352
rect 3016 18340 3022 18352
rect 3053 18343 3111 18349
rect 3053 18340 3065 18343
rect 3016 18312 3065 18340
rect 3016 18300 3022 18312
rect 3053 18309 3065 18312
rect 3099 18309 3111 18343
rect 3053 18303 3111 18309
rect 3068 18272 3096 18303
rect 4430 18300 4436 18352
rect 4488 18340 4494 18352
rect 6549 18343 6607 18349
rect 6549 18340 6561 18343
rect 4488 18312 6561 18340
rect 4488 18300 4494 18312
rect 6549 18309 6561 18312
rect 6595 18340 6607 18343
rect 7190 18340 7196 18352
rect 6595 18312 7196 18340
rect 6595 18309 6607 18312
rect 6549 18303 6607 18309
rect 7190 18300 7196 18312
rect 7248 18300 7254 18352
rect 12434 18300 12440 18352
rect 12492 18340 12498 18352
rect 12492 18312 12934 18340
rect 12492 18300 12498 18312
rect 4341 18275 4399 18281
rect 3068 18244 3740 18272
rect 1694 18176 2544 18204
rect 3513 18207 3571 18213
rect 1694 18173 1706 18176
rect 1648 18167 1706 18173
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 3605 18207 3663 18213
rect 3605 18204 3617 18207
rect 3559 18176 3617 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 3605 18173 3617 18176
rect 3651 18173 3663 18207
rect 3605 18167 3663 18173
rect 1719 18071 1777 18077
rect 1719 18037 1731 18071
rect 1765 18068 1777 18071
rect 1946 18068 1952 18080
rect 1765 18040 1952 18068
rect 1765 18037 1777 18040
rect 1719 18031 1777 18037
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2593 18071 2651 18077
rect 2593 18037 2605 18071
rect 2639 18068 2651 18071
rect 2958 18068 2964 18080
rect 2639 18040 2964 18068
rect 2639 18037 2651 18040
rect 2593 18031 2651 18037
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 3620 18068 3648 18167
rect 3712 18136 3740 18244
rect 4341 18241 4353 18275
rect 4387 18272 4399 18275
rect 7742 18272 7748 18284
rect 4387 18244 7748 18272
rect 4387 18241 4399 18244
rect 4341 18235 4399 18241
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 8021 18275 8079 18281
rect 8021 18241 8033 18275
rect 8067 18272 8079 18275
rect 8110 18272 8116 18284
rect 8067 18244 8116 18272
rect 8067 18241 8079 18244
rect 8021 18235 8079 18241
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 11517 18275 11575 18281
rect 10367 18244 11376 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 11348 18216 11376 18244
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 12802 18272 12808 18284
rect 11563 18244 12808 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 12906 18272 12934 18312
rect 14734 18272 14740 18284
rect 12906 18244 14136 18272
rect 14695 18244 14740 18272
rect 4062 18204 4068 18216
rect 4023 18176 4068 18204
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 5166 18204 5172 18216
rect 5127 18176 5172 18204
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 5721 18207 5779 18213
rect 5721 18204 5733 18207
rect 5316 18176 5733 18204
rect 5316 18164 5322 18176
rect 5721 18173 5733 18176
rect 5767 18204 5779 18207
rect 6086 18204 6092 18216
rect 5767 18176 6092 18204
rect 5767 18173 5779 18176
rect 5721 18167 5779 18173
rect 6086 18164 6092 18176
rect 6144 18164 6150 18216
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 9217 18207 9275 18213
rect 9217 18204 9229 18207
rect 9088 18176 9229 18204
rect 9088 18164 9094 18176
rect 9217 18173 9229 18176
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 10781 18207 10839 18213
rect 9732 18176 9777 18204
rect 9732 18164 9738 18176
rect 10781 18173 10793 18207
rect 10827 18173 10839 18207
rect 11330 18204 11336 18216
rect 11291 18176 11336 18204
rect 10781 18167 10839 18173
rect 5442 18136 5448 18148
rect 3712 18108 5448 18136
rect 5442 18096 5448 18108
rect 5500 18096 5506 18148
rect 5905 18139 5963 18145
rect 5905 18105 5917 18139
rect 5951 18136 5963 18139
rect 6730 18136 6736 18148
rect 5951 18108 6736 18136
rect 5951 18105 5963 18108
rect 5905 18099 5963 18105
rect 6730 18096 6736 18108
rect 6788 18096 6794 18148
rect 7377 18139 7435 18145
rect 7377 18105 7389 18139
rect 7423 18105 7435 18139
rect 7377 18099 7435 18105
rect 4430 18068 4436 18080
rect 3620 18040 4436 18068
rect 4430 18028 4436 18040
rect 4488 18028 4494 18080
rect 6273 18071 6331 18077
rect 6273 18037 6285 18071
rect 6319 18068 6331 18071
rect 6546 18068 6552 18080
rect 6319 18040 6552 18068
rect 6319 18037 6331 18040
rect 6273 18031 6331 18037
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 7392 18068 7420 18099
rect 7466 18096 7472 18148
rect 7524 18136 7530 18148
rect 9950 18136 9956 18148
rect 7524 18108 7569 18136
rect 9911 18108 9956 18136
rect 7524 18096 7530 18108
rect 9950 18096 9956 18108
rect 10008 18096 10014 18148
rect 8294 18068 8300 18080
rect 7392 18040 8300 18068
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 8662 18068 8668 18080
rect 8623 18040 8668 18068
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 10689 18071 10747 18077
rect 10689 18037 10701 18071
rect 10735 18068 10747 18071
rect 10796 18068 10824 18167
rect 11330 18164 11336 18176
rect 11388 18164 11394 18216
rect 12906 18213 12934 18244
rect 14108 18216 14136 18244
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18204 12127 18207
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12115 18176 12449 18204
rect 12115 18173 12127 18176
rect 12069 18167 12127 18173
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18173 12955 18207
rect 13909 18207 13967 18213
rect 13909 18204 13921 18207
rect 12897 18167 12955 18173
rect 13786 18176 13921 18204
rect 13170 18136 13176 18148
rect 13131 18108 13176 18136
rect 13170 18096 13176 18108
rect 13228 18096 13234 18148
rect 11330 18068 11336 18080
rect 10735 18040 11336 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 11790 18068 11796 18080
rect 11751 18040 11796 18068
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 13786 18068 13814 18176
rect 13909 18173 13921 18176
rect 13955 18204 13967 18207
rect 14001 18207 14059 18213
rect 14001 18204 14013 18207
rect 13955 18176 14013 18204
rect 13955 18173 13967 18176
rect 13909 18167 13967 18173
rect 14001 18173 14013 18176
rect 14047 18173 14059 18207
rect 14001 18167 14059 18173
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 14148 18176 14473 18204
rect 14148 18164 14154 18176
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 14461 18167 14519 18173
rect 15856 18136 15884 18380
rect 17034 18368 17040 18380
rect 17092 18368 17098 18420
rect 18782 18368 18788 18420
rect 18840 18408 18846 18420
rect 19061 18411 19119 18417
rect 19061 18408 19073 18411
rect 18840 18380 19073 18408
rect 18840 18368 18846 18380
rect 19061 18377 19073 18380
rect 19107 18408 19119 18411
rect 19518 18408 19524 18420
rect 19107 18380 19524 18408
rect 19107 18377 19119 18380
rect 19061 18371 19119 18377
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 20070 18408 20076 18420
rect 20031 18380 20076 18408
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 16574 18340 16580 18352
rect 16040 18312 16580 18340
rect 16040 18281 16068 18312
rect 16574 18300 16580 18312
rect 16632 18300 16638 18352
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18241 16083 18275
rect 16482 18272 16488 18284
rect 16443 18244 16488 18272
rect 16025 18235 16083 18241
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 16666 18232 16672 18284
rect 16724 18272 16730 18284
rect 16724 18244 19564 18272
rect 16724 18232 16730 18244
rect 18668 18207 18726 18213
rect 18668 18173 18680 18207
rect 18714 18204 18726 18207
rect 18782 18204 18788 18216
rect 18714 18176 18788 18204
rect 18714 18173 18726 18176
rect 18668 18167 18726 18173
rect 18782 18164 18788 18176
rect 18840 18204 18846 18216
rect 19429 18207 19487 18213
rect 19429 18204 19441 18207
rect 18840 18176 19441 18204
rect 18840 18164 18846 18176
rect 19429 18173 19441 18176
rect 19475 18173 19487 18207
rect 19536 18204 19564 18244
rect 19648 18207 19706 18213
rect 19648 18204 19660 18207
rect 19536 18176 19660 18204
rect 19429 18167 19487 18173
rect 19648 18173 19660 18176
rect 19694 18204 19706 18207
rect 20441 18207 20499 18213
rect 20441 18204 20453 18207
rect 19694 18176 20453 18204
rect 19694 18173 19706 18176
rect 19648 18167 19706 18173
rect 20441 18173 20453 18176
rect 20487 18204 20499 18207
rect 20530 18204 20536 18216
rect 20487 18176 20536 18204
rect 20487 18173 20499 18176
rect 20441 18167 20499 18173
rect 20530 18164 20536 18176
rect 20588 18164 20594 18216
rect 16117 18139 16175 18145
rect 16117 18136 16129 18139
rect 15856 18108 16129 18136
rect 16117 18105 16129 18108
rect 16163 18105 16175 18139
rect 16117 18099 16175 18105
rect 17954 18096 17960 18148
rect 18012 18136 18018 18148
rect 19751 18139 19809 18145
rect 19751 18136 19763 18139
rect 18012 18108 19763 18136
rect 18012 18096 18018 18108
rect 19751 18105 19763 18108
rect 19797 18105 19809 18139
rect 19751 18099 19809 18105
rect 13596 18040 13814 18068
rect 15381 18071 15439 18077
rect 13596 18028 13602 18040
rect 15381 18037 15393 18071
rect 15427 18068 15439 18071
rect 15470 18068 15476 18080
rect 15427 18040 15476 18068
rect 15427 18037 15439 18040
rect 15381 18031 15439 18037
rect 15470 18028 15476 18040
rect 15528 18028 15534 18080
rect 17402 18068 17408 18080
rect 17363 18040 17408 18068
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 18739 18071 18797 18077
rect 18739 18037 18751 18071
rect 18785 18068 18797 18071
rect 18966 18068 18972 18080
rect 18785 18040 18972 18068
rect 18785 18037 18797 18040
rect 18739 18031 18797 18037
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 20622 18068 20628 18080
rect 20583 18040 20628 18068
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 21174 18028 21180 18080
rect 21232 18068 21238 18080
rect 21637 18071 21695 18077
rect 21637 18068 21649 18071
rect 21232 18040 21649 18068
rect 21232 18028 21238 18040
rect 21637 18037 21649 18040
rect 21683 18037 21695 18071
rect 21637 18031 21695 18037
rect 24118 18028 24124 18080
rect 24176 18068 24182 18080
rect 24581 18071 24639 18077
rect 24581 18068 24593 18071
rect 24176 18040 24593 18068
rect 24176 18028 24182 18040
rect 24581 18037 24593 18040
rect 24627 18037 24639 18071
rect 24581 18031 24639 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 3697 17867 3755 17873
rect 3697 17833 3709 17867
rect 3743 17864 3755 17867
rect 4062 17864 4068 17876
rect 3743 17836 4068 17864
rect 3743 17833 3755 17836
rect 3697 17827 3755 17833
rect 4062 17824 4068 17836
rect 4120 17864 4126 17876
rect 5445 17867 5503 17873
rect 5445 17864 5457 17867
rect 4120 17836 5457 17864
rect 4120 17824 4126 17836
rect 5445 17833 5457 17836
rect 5491 17833 5503 17867
rect 6362 17864 6368 17876
rect 6323 17836 6368 17864
rect 5445 17827 5503 17833
rect 6362 17824 6368 17836
rect 6420 17824 6426 17876
rect 6917 17867 6975 17873
rect 6917 17833 6929 17867
rect 6963 17864 6975 17867
rect 7377 17867 7435 17873
rect 7377 17864 7389 17867
rect 6963 17836 7389 17864
rect 6963 17833 6975 17836
rect 6917 17827 6975 17833
rect 7377 17833 7389 17836
rect 7423 17864 7435 17867
rect 7466 17864 7472 17876
rect 7423 17836 7472 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 10134 17864 10140 17876
rect 10095 17836 10140 17864
rect 10134 17824 10140 17836
rect 10192 17824 10198 17876
rect 13081 17867 13139 17873
rect 13081 17833 13093 17867
rect 13127 17864 13139 17867
rect 13170 17864 13176 17876
rect 13127 17836 13176 17864
rect 13127 17833 13139 17836
rect 13081 17827 13139 17833
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 16485 17867 16543 17873
rect 16485 17864 16497 17867
rect 16172 17836 16497 17864
rect 16172 17824 16178 17836
rect 16485 17833 16497 17836
rect 16531 17864 16543 17867
rect 18417 17867 18475 17873
rect 18417 17864 18429 17867
rect 16531 17836 18429 17864
rect 16531 17833 16543 17836
rect 16485 17827 16543 17833
rect 18417 17833 18429 17836
rect 18463 17833 18475 17867
rect 18417 17827 18475 17833
rect 5166 17796 5172 17808
rect 4724 17768 5172 17796
rect 4724 17740 4752 17768
rect 5166 17756 5172 17768
rect 5224 17756 5230 17808
rect 7926 17796 7932 17808
rect 7887 17768 7932 17796
rect 7926 17756 7932 17768
rect 7984 17756 7990 17808
rect 8110 17756 8116 17808
rect 8168 17796 8174 17808
rect 8481 17799 8539 17805
rect 8481 17796 8493 17799
rect 8168 17768 8493 17796
rect 8168 17756 8174 17768
rect 8481 17765 8493 17768
rect 8527 17765 8539 17799
rect 8481 17759 8539 17765
rect 10597 17799 10655 17805
rect 10597 17765 10609 17799
rect 10643 17796 10655 17799
rect 10778 17796 10784 17808
rect 10643 17768 10784 17796
rect 10643 17765 10655 17768
rect 10597 17759 10655 17765
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 14277 17799 14335 17805
rect 14277 17765 14289 17799
rect 14323 17796 14335 17799
rect 15286 17796 15292 17808
rect 14323 17768 15292 17796
rect 14323 17765 14335 17768
rect 14277 17759 14335 17765
rect 15286 17756 15292 17768
rect 15344 17796 15350 17808
rect 16025 17799 16083 17805
rect 16025 17796 16037 17799
rect 15344 17768 16037 17796
rect 15344 17756 15350 17768
rect 16025 17765 16037 17768
rect 16071 17765 16083 17799
rect 16850 17796 16856 17808
rect 16811 17768 16856 17796
rect 16025 17759 16083 17765
rect 16850 17756 16856 17768
rect 16908 17756 16914 17808
rect 17402 17756 17408 17808
rect 17460 17796 17466 17808
rect 17460 17768 18828 17796
rect 17460 17756 17466 17768
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 2314 17728 2320 17740
rect 1995 17700 2320 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 4706 17728 4712 17740
rect 4619 17700 4712 17728
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 4985 17731 5043 17737
rect 4985 17697 4997 17731
rect 5031 17728 5043 17731
rect 5350 17728 5356 17740
rect 5031 17700 5356 17728
rect 5031 17697 5043 17700
rect 4985 17691 5043 17697
rect 5350 17688 5356 17700
rect 5408 17728 5414 17740
rect 6546 17728 6552 17740
rect 5408 17700 6552 17728
rect 5408 17688 5414 17700
rect 6546 17688 6552 17700
rect 6604 17688 6610 17740
rect 11974 17728 11980 17740
rect 11935 17700 11980 17728
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 12434 17728 12440 17740
rect 12395 17700 12440 17728
rect 12434 17688 12440 17700
rect 12492 17688 12498 17740
rect 13817 17731 13875 17737
rect 13817 17697 13829 17731
rect 13863 17697 13875 17731
rect 14090 17728 14096 17740
rect 14051 17700 14096 17728
rect 13817 17691 13875 17697
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 3326 17660 3332 17672
rect 3007 17632 3332 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 3326 17620 3332 17632
rect 3384 17620 3390 17672
rect 5169 17663 5227 17669
rect 5169 17629 5181 17663
rect 5215 17660 5227 17663
rect 5997 17663 6055 17669
rect 5997 17660 6009 17663
rect 5215 17632 6009 17660
rect 5215 17629 5227 17632
rect 5169 17623 5227 17629
rect 5997 17629 6009 17632
rect 6043 17660 6055 17663
rect 6822 17660 6828 17672
rect 6043 17632 6828 17660
rect 6043 17629 6055 17632
rect 5997 17623 6055 17629
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17660 7895 17663
rect 8662 17660 8668 17672
rect 7883 17632 8668 17660
rect 7883 17629 7895 17632
rect 7837 17623 7895 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17660 10563 17663
rect 10686 17660 10692 17672
rect 10551 17632 10692 17660
rect 10551 17629 10563 17632
rect 10505 17623 10563 17629
rect 10686 17620 10692 17632
rect 10744 17620 10750 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17629 10839 17663
rect 12526 17660 12532 17672
rect 12487 17632 12532 17660
rect 10781 17623 10839 17629
rect 8294 17552 8300 17604
rect 8352 17592 8358 17604
rect 10796 17592 10824 17623
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 13832 17660 13860 17691
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 15632 17731 15690 17737
rect 15632 17697 15644 17731
rect 15678 17728 15690 17731
rect 15930 17728 15936 17740
rect 15678 17700 15936 17728
rect 15678 17697 15690 17700
rect 15632 17691 15690 17697
rect 15930 17688 15936 17700
rect 15988 17688 15994 17740
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 16666 17728 16672 17740
rect 16623 17700 16672 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 16666 17688 16672 17700
rect 16724 17728 16730 17740
rect 17126 17728 17132 17740
rect 16724 17700 17132 17728
rect 16724 17688 16730 17700
rect 17126 17688 17132 17700
rect 17184 17688 17190 17740
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17728 18659 17731
rect 18690 17728 18696 17740
rect 18647 17700 18696 17728
rect 18647 17697 18659 17700
rect 18601 17691 18659 17697
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 18800 17737 18828 17768
rect 20990 17737 20996 17740
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17697 18843 17731
rect 20936 17731 20996 17737
rect 20936 17728 20948 17731
rect 18785 17691 18843 17697
rect 20869 17700 20948 17728
rect 13906 17660 13912 17672
rect 13819 17632 13912 17660
rect 13906 17620 13912 17632
rect 13964 17660 13970 17672
rect 16758 17660 16764 17672
rect 13964 17632 16764 17660
rect 13964 17620 13970 17632
rect 16758 17620 16764 17632
rect 16816 17660 16822 17672
rect 17034 17660 17040 17672
rect 16816 17632 17040 17660
rect 16816 17620 16822 17632
rect 17034 17620 17040 17632
rect 17092 17620 17098 17672
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 20869 17660 20897 17700
rect 20936 17697 20948 17700
rect 20982 17697 20996 17731
rect 20936 17691 20996 17697
rect 20990 17688 20996 17691
rect 21048 17688 21054 17740
rect 22256 17731 22314 17737
rect 22256 17697 22268 17731
rect 22302 17728 22314 17731
rect 22554 17728 22560 17740
rect 22302 17700 22560 17728
rect 22302 17697 22314 17700
rect 22256 17691 22314 17697
rect 22554 17688 22560 17700
rect 22612 17688 22618 17740
rect 23268 17731 23326 17737
rect 23268 17697 23280 17731
rect 23314 17728 23326 17731
rect 23566 17728 23572 17740
rect 23314 17700 23572 17728
rect 23314 17697 23326 17700
rect 23268 17691 23326 17697
rect 23566 17688 23572 17700
rect 23624 17688 23630 17740
rect 17276 17632 20897 17660
rect 17276 17620 17282 17632
rect 11698 17592 11704 17604
rect 8352 17564 11704 17592
rect 8352 17552 8358 17564
rect 11698 17552 11704 17564
rect 11756 17552 11762 17604
rect 15703 17595 15761 17601
rect 15703 17561 15715 17595
rect 15749 17592 15761 17595
rect 19242 17592 19248 17604
rect 15749 17564 19248 17592
rect 15749 17561 15761 17564
rect 15703 17555 15761 17561
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 1762 17484 1768 17536
rect 1820 17524 1826 17536
rect 2133 17527 2191 17533
rect 2133 17524 2145 17527
rect 1820 17496 2145 17524
rect 1820 17484 1826 17496
rect 2133 17493 2145 17496
rect 2179 17493 2191 17527
rect 2133 17487 2191 17493
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 4798 17524 4804 17536
rect 4387 17496 4804 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 9309 17527 9367 17533
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9674 17524 9680 17536
rect 9355 17496 9680 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9674 17484 9680 17496
rect 9732 17524 9738 17536
rect 10134 17524 10140 17536
rect 9732 17496 10140 17524
rect 9732 17484 9738 17496
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 14366 17484 14372 17536
rect 14424 17524 14430 17536
rect 14553 17527 14611 17533
rect 14553 17524 14565 17527
rect 14424 17496 14565 17524
rect 14424 17484 14430 17496
rect 14553 17493 14565 17496
rect 14599 17493 14611 17527
rect 14553 17487 14611 17493
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 17218 17524 17224 17536
rect 15620 17496 17224 17524
rect 15620 17484 15626 17496
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 17494 17524 17500 17536
rect 17455 17496 17500 17524
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 18141 17527 18199 17533
rect 18141 17493 18153 17527
rect 18187 17524 18199 17527
rect 18230 17524 18236 17536
rect 18187 17496 18236 17524
rect 18187 17493 18199 17496
rect 18141 17487 18199 17493
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 20254 17484 20260 17536
rect 20312 17524 20318 17536
rect 21039 17527 21097 17533
rect 21039 17524 21051 17527
rect 20312 17496 21051 17524
rect 20312 17484 20318 17496
rect 21039 17493 21051 17496
rect 21085 17493 21097 17527
rect 21039 17487 21097 17493
rect 21726 17484 21732 17536
rect 21784 17524 21790 17536
rect 22327 17527 22385 17533
rect 22327 17524 22339 17527
rect 21784 17496 22339 17524
rect 21784 17484 21790 17496
rect 22327 17493 22339 17496
rect 22373 17493 22385 17527
rect 22327 17487 22385 17493
rect 22462 17484 22468 17536
rect 22520 17524 22526 17536
rect 23339 17527 23397 17533
rect 23339 17524 23351 17527
rect 22520 17496 23351 17524
rect 22520 17484 22526 17496
rect 23339 17493 23351 17496
rect 23385 17493 23397 17527
rect 23339 17487 23397 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 4525 17323 4583 17329
rect 4525 17289 4537 17323
rect 4571 17320 4583 17323
rect 4706 17320 4712 17332
rect 4571 17292 4712 17320
rect 4571 17289 4583 17292
rect 4525 17283 4583 17289
rect 4706 17280 4712 17292
rect 4764 17280 4770 17332
rect 7745 17323 7803 17329
rect 7745 17289 7757 17323
rect 7791 17320 7803 17323
rect 7926 17320 7932 17332
rect 7791 17292 7932 17320
rect 7791 17289 7803 17292
rect 7745 17283 7803 17289
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 11701 17323 11759 17329
rect 8076 17292 8121 17320
rect 8076 17280 8082 17292
rect 11701 17289 11713 17323
rect 11747 17320 11759 17323
rect 12434 17320 12440 17332
rect 11747 17292 12440 17320
rect 11747 17289 11759 17292
rect 11701 17283 11759 17289
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 13262 17280 13268 17332
rect 13320 17320 13326 17332
rect 13906 17320 13912 17332
rect 13320 17292 13814 17320
rect 13867 17292 13912 17320
rect 13320 17280 13326 17292
rect 2041 17255 2099 17261
rect 2041 17221 2053 17255
rect 2087 17252 2099 17255
rect 6178 17252 6184 17264
rect 2087 17224 6184 17252
rect 2087 17221 2099 17224
rect 2041 17215 2099 17221
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2056 17116 2084 17215
rect 6178 17212 6184 17224
rect 6236 17252 6242 17264
rect 7837 17255 7895 17261
rect 7837 17252 7849 17255
rect 6236 17224 7849 17252
rect 6236 17212 6242 17224
rect 7837 17221 7849 17224
rect 7883 17221 7895 17255
rect 7837 17215 7895 17221
rect 2958 17144 2964 17196
rect 3016 17184 3022 17196
rect 5721 17187 5779 17193
rect 3016 17156 4568 17184
rect 3016 17144 3022 17156
rect 1443 17088 2084 17116
rect 2593 17119 2651 17125
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2593 17085 2605 17119
rect 2639 17116 2651 17119
rect 3672 17119 3730 17125
rect 2639 17088 3004 17116
rect 2639 17085 2651 17088
rect 2593 17079 2651 17085
rect 2976 16992 3004 17088
rect 3672 17085 3684 17119
rect 3718 17116 3730 17119
rect 4154 17116 4160 17128
rect 3718 17088 4160 17116
rect 3718 17085 3730 17088
rect 3672 17079 3730 17085
rect 4154 17076 4160 17088
rect 4212 17116 4218 17128
rect 4212 17088 4305 17116
rect 4212 17076 4218 17088
rect 3881 17051 3939 17057
rect 3881 17017 3893 17051
rect 3927 17048 3939 17051
rect 4338 17048 4344 17060
rect 3927 17020 4344 17048
rect 3927 17017 3939 17020
rect 3881 17011 3939 17017
rect 4338 17008 4344 17020
rect 4396 17008 4402 17060
rect 4540 17048 4568 17156
rect 5721 17153 5733 17187
rect 5767 17184 5779 17187
rect 6546 17184 6552 17196
rect 5767 17156 6552 17184
rect 5767 17153 5779 17156
rect 5721 17147 5779 17153
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6788 17156 6837 17184
rect 6788 17144 6794 17156
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 8036 17184 8064 17280
rect 13786 17252 13814 17292
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 17402 17320 17408 17332
rect 16960 17292 17408 17320
rect 16960 17252 16988 17292
rect 17402 17280 17408 17292
rect 17460 17320 17466 17332
rect 17773 17323 17831 17329
rect 17773 17320 17785 17323
rect 17460 17292 17785 17320
rect 17460 17280 17466 17292
rect 17773 17289 17785 17292
rect 17819 17289 17831 17323
rect 24762 17320 24768 17332
rect 24723 17292 24768 17320
rect 17773 17283 17831 17289
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 13786 17224 16988 17252
rect 17037 17255 17095 17261
rect 17037 17221 17049 17255
rect 17083 17252 17095 17255
rect 18230 17252 18236 17264
rect 17083 17224 18236 17252
rect 17083 17221 17095 17224
rect 17037 17215 17095 17221
rect 18230 17212 18236 17224
rect 18288 17212 18294 17264
rect 18506 17212 18512 17264
rect 18564 17252 18570 17264
rect 18564 17224 21864 17252
rect 18564 17212 18570 17224
rect 21836 17196 21864 17224
rect 8573 17187 8631 17193
rect 8573 17184 8585 17187
rect 8036 17156 8585 17184
rect 6825 17147 6883 17153
rect 8573 17153 8585 17156
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 10413 17187 10471 17193
rect 10413 17153 10425 17187
rect 10459 17184 10471 17187
rect 11238 17184 11244 17196
rect 10459 17156 11244 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 14366 17184 14372 17196
rect 13587 17156 14372 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 16114 17184 16120 17196
rect 16075 17156 16120 17184
rect 16114 17144 16120 17156
rect 16172 17144 16178 17196
rect 18322 17144 18328 17196
rect 18380 17184 18386 17196
rect 20763 17187 20821 17193
rect 20763 17184 20775 17187
rect 18380 17156 20775 17184
rect 18380 17144 18386 17156
rect 20763 17153 20775 17156
rect 20809 17153 20821 17187
rect 20763 17147 20821 17153
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 21048 17156 21097 17184
rect 21048 17144 21054 17156
rect 21085 17153 21097 17156
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 21818 17144 21824 17196
rect 21876 17184 21882 17196
rect 22097 17187 22155 17193
rect 22097 17184 22109 17187
rect 21876 17156 22109 17184
rect 21876 17144 21882 17156
rect 22097 17153 22109 17156
rect 22143 17153 22155 17187
rect 22097 17147 22155 17153
rect 5994 17076 6000 17128
rect 6052 17116 6058 17128
rect 9122 17116 9128 17128
rect 6052 17088 9128 17116
rect 6052 17076 6058 17088
rect 9122 17076 9128 17088
rect 9180 17076 9186 17128
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17085 12863 17119
rect 13262 17116 13268 17128
rect 13223 17088 13268 17116
rect 12805 17079 12863 17085
rect 4706 17048 4712 17060
rect 4540 17020 4712 17048
rect 4706 17008 4712 17020
rect 4764 17008 4770 17060
rect 4798 17008 4804 17060
rect 4856 17048 4862 17060
rect 5350 17048 5356 17060
rect 4856 17020 4901 17048
rect 5311 17020 5356 17048
rect 4856 17008 4862 17020
rect 5350 17008 5356 17020
rect 5408 17008 5414 17060
rect 7146 17051 7204 17057
rect 7146 17017 7158 17051
rect 7192 17017 7204 17051
rect 7146 17011 7204 17017
rect 7837 17051 7895 17057
rect 7837 17017 7849 17051
rect 7883 17048 7895 17051
rect 8570 17048 8576 17060
rect 7883 17020 8576 17048
rect 7883 17017 7895 17020
rect 7837 17011 7895 17017
rect 2314 16980 2320 16992
rect 2275 16952 2320 16980
rect 2314 16940 2320 16952
rect 2372 16940 2378 16992
rect 2774 16980 2780 16992
rect 2735 16952 2780 16980
rect 2774 16940 2780 16952
rect 2832 16940 2838 16992
rect 2958 16940 2964 16992
rect 3016 16980 3022 16992
rect 3053 16983 3111 16989
rect 3053 16980 3065 16983
rect 3016 16952 3065 16980
rect 3016 16940 3022 16952
rect 3053 16949 3065 16952
rect 3099 16949 3111 16983
rect 3053 16943 3111 16949
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 5997 16983 6055 16989
rect 5997 16980 6009 16983
rect 4304 16952 6009 16980
rect 4304 16940 4310 16952
rect 5997 16949 6009 16952
rect 6043 16980 6055 16983
rect 6362 16980 6368 16992
rect 6043 16952 6368 16980
rect 6043 16949 6055 16952
rect 5997 16943 6055 16949
rect 6362 16940 6368 16952
rect 6420 16980 6426 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6420 16952 6561 16980
rect 6420 16940 6426 16952
rect 6549 16949 6561 16952
rect 6595 16980 6607 16983
rect 7006 16980 7012 16992
rect 6595 16952 7012 16980
rect 6595 16949 6607 16952
rect 6549 16943 6607 16949
rect 7006 16940 7012 16952
rect 7064 16980 7070 16992
rect 7161 16980 7189 17011
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 8894 17051 8952 17057
rect 8894 17017 8906 17051
rect 8940 17048 8952 17051
rect 9674 17048 9680 17060
rect 8940 17020 9680 17048
rect 8940 17017 8952 17020
rect 8894 17011 8952 17017
rect 8389 16983 8447 16989
rect 8389 16980 8401 16983
rect 7064 16952 8401 16980
rect 7064 16940 7070 16952
rect 8389 16949 8401 16952
rect 8435 16980 8447 16983
rect 8909 16980 8937 17011
rect 9674 17008 9680 17020
rect 9732 17008 9738 17060
rect 10505 17051 10563 17057
rect 10505 17017 10517 17051
rect 10551 17048 10563 17051
rect 10778 17048 10784 17060
rect 10551 17020 10784 17048
rect 10551 17017 10563 17020
rect 10505 17011 10563 17017
rect 9490 16980 9496 16992
rect 8435 16952 8937 16980
rect 9451 16952 9496 16980
rect 8435 16949 8447 16952
rect 8389 16943 8447 16949
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 9861 16983 9919 16989
rect 9861 16949 9873 16983
rect 9907 16980 9919 16983
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 9907 16952 10241 16980
rect 9907 16949 9919 16952
rect 9861 16943 9919 16949
rect 10229 16949 10241 16952
rect 10275 16980 10287 16983
rect 10520 16980 10548 17011
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 10870 17008 10876 17060
rect 10928 17048 10934 17060
rect 11057 17051 11115 17057
rect 11057 17048 11069 17051
rect 10928 17020 11069 17048
rect 10928 17008 10934 17020
rect 11057 17017 11069 17020
rect 11103 17017 11115 17051
rect 11057 17011 11115 17017
rect 12820 17048 12848 17079
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 15657 17119 15715 17125
rect 15657 17085 15669 17119
rect 15703 17116 15715 17119
rect 15930 17116 15936 17128
rect 15703 17088 15936 17116
rect 15703 17085 15715 17088
rect 15657 17079 15715 17085
rect 15930 17076 15936 17088
rect 15988 17076 15994 17128
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 19648 17119 19706 17125
rect 19648 17116 19660 17119
rect 19484 17088 19660 17116
rect 19484 17076 19490 17088
rect 19648 17085 19660 17088
rect 19694 17116 19706 17119
rect 20073 17119 20131 17125
rect 20073 17116 20085 17119
rect 19694 17088 20085 17116
rect 19694 17085 19706 17088
rect 19648 17079 19706 17085
rect 20073 17085 20085 17088
rect 20119 17085 20131 17119
rect 20073 17079 20131 17085
rect 20346 17076 20352 17128
rect 20404 17116 20410 17128
rect 20660 17119 20718 17125
rect 20660 17116 20672 17119
rect 20404 17088 20672 17116
rect 20404 17076 20410 17088
rect 20660 17085 20672 17088
rect 20706 17116 20718 17119
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 20706 17088 21465 17116
rect 20706 17085 20718 17088
rect 20660 17079 20718 17085
rect 21453 17085 21465 17088
rect 21499 17085 21511 17119
rect 21453 17079 21511 17085
rect 21688 17119 21746 17125
rect 21688 17085 21700 17119
rect 21734 17116 21746 17119
rect 21836 17116 21864 17144
rect 22554 17116 22560 17128
rect 21734 17088 21864 17116
rect 22467 17088 22560 17116
rect 21734 17085 21746 17088
rect 21688 17079 21746 17085
rect 22554 17076 22560 17088
rect 22612 17116 22618 17128
rect 23290 17116 23296 17128
rect 22612 17088 23296 17116
rect 22612 17076 22618 17088
rect 23290 17076 23296 17088
rect 23348 17076 23354 17128
rect 24578 17116 24584 17128
rect 24539 17088 24584 17116
rect 24578 17076 24584 17088
rect 24636 17116 24642 17128
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24636 17088 25145 17116
rect 24636 17076 24642 17088
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 13538 17048 13544 17060
rect 12820 17020 13544 17048
rect 12820 16992 12848 17020
rect 13538 17008 13544 17020
rect 13596 17008 13602 17060
rect 14690 17051 14748 17057
rect 14690 17048 14702 17051
rect 14200 17020 14702 17048
rect 14200 16992 14228 17020
rect 14690 17017 14702 17020
rect 14736 17048 14748 17051
rect 15470 17048 15476 17060
rect 14736 17020 15476 17048
rect 14736 17017 14748 17020
rect 14690 17011 14748 17017
rect 15470 17008 15476 17020
rect 15528 17048 15534 17060
rect 16025 17051 16083 17057
rect 16025 17048 16037 17051
rect 15528 17020 16037 17048
rect 15528 17008 15534 17020
rect 16025 17017 16037 17020
rect 16071 17048 16083 17051
rect 16438 17051 16496 17057
rect 16438 17048 16450 17051
rect 16071 17020 16450 17048
rect 16071 17017 16083 17020
rect 16025 17011 16083 17017
rect 16438 17017 16450 17020
rect 16484 17048 16496 17051
rect 16850 17048 16856 17060
rect 16484 17020 16856 17048
rect 16484 17017 16496 17020
rect 16438 17011 16496 17017
rect 16850 17008 16856 17020
rect 16908 17048 16914 17060
rect 17313 17051 17371 17057
rect 17313 17048 17325 17051
rect 16908 17020 17325 17048
rect 16908 17008 16914 17020
rect 17313 17017 17325 17020
rect 17359 17017 17371 17051
rect 18138 17048 18144 17060
rect 18099 17020 18144 17048
rect 17313 17011 17371 17017
rect 18138 17008 18144 17020
rect 18196 17008 18202 17060
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 18782 17048 18788 17060
rect 18288 17020 18333 17048
rect 18743 17020 18788 17048
rect 18288 17008 18294 17020
rect 18782 17008 18788 17020
rect 18840 17008 18846 17060
rect 21358 17008 21364 17060
rect 21416 17048 21422 17060
rect 21775 17051 21833 17057
rect 21775 17048 21787 17051
rect 21416 17020 21787 17048
rect 21416 17008 21422 17020
rect 21775 17017 21787 17020
rect 21821 17017 21833 17051
rect 21775 17011 21833 17017
rect 10275 16952 10548 16980
rect 10275 16949 10287 16952
rect 10229 16943 10287 16949
rect 10962 16940 10968 16992
rect 11020 16980 11026 16992
rect 11974 16980 11980 16992
rect 11020 16952 11980 16980
rect 11020 16940 11026 16952
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12713 16983 12771 16989
rect 12713 16949 12725 16983
rect 12759 16980 12771 16983
rect 12802 16980 12808 16992
rect 12759 16952 12808 16980
rect 12759 16949 12771 16952
rect 12713 16943 12771 16949
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 14182 16980 14188 16992
rect 14143 16952 14188 16980
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 15286 16980 15292 16992
rect 15247 16952 15292 16980
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 18690 16940 18696 16992
rect 18748 16980 18754 16992
rect 19061 16983 19119 16989
rect 19061 16980 19073 16983
rect 18748 16952 19073 16980
rect 18748 16940 18754 16952
rect 19061 16949 19073 16952
rect 19107 16949 19119 16983
rect 19061 16943 19119 16949
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 19751 16983 19809 16989
rect 19751 16980 19763 16983
rect 19576 16952 19763 16980
rect 19576 16940 19582 16952
rect 19751 16949 19763 16952
rect 19797 16949 19809 16983
rect 19751 16943 19809 16949
rect 23293 16983 23351 16989
rect 23293 16949 23305 16983
rect 23339 16980 23351 16983
rect 23566 16980 23572 16992
rect 23339 16952 23572 16980
rect 23339 16949 23351 16952
rect 23293 16943 23351 16949
rect 23566 16940 23572 16952
rect 23624 16940 23630 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 4985 16779 5043 16785
rect 4985 16745 4997 16779
rect 5031 16776 5043 16779
rect 6822 16776 6828 16788
rect 5031 16748 6040 16776
rect 6783 16748 6828 16776
rect 5031 16745 5043 16748
rect 4985 16739 5043 16745
rect 6012 16720 6040 16748
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 7561 16779 7619 16785
rect 7561 16745 7573 16779
rect 7607 16776 7619 16779
rect 7926 16776 7932 16788
rect 7607 16748 7932 16776
rect 7607 16745 7619 16748
rect 7561 16739 7619 16745
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8662 16776 8668 16788
rect 8623 16748 8668 16776
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 9490 16736 9496 16788
rect 9548 16776 9554 16788
rect 10686 16776 10692 16788
rect 9548 16748 9904 16776
rect 10647 16748 10692 16776
rect 9548 16736 9554 16748
rect 4246 16668 4252 16720
rect 4304 16708 4310 16720
rect 4427 16711 4485 16717
rect 4427 16708 4439 16711
rect 4304 16680 4439 16708
rect 4304 16668 4310 16680
rect 4427 16677 4439 16680
rect 4473 16677 4485 16711
rect 4427 16671 4485 16677
rect 4706 16668 4712 16720
rect 4764 16708 4770 16720
rect 5261 16711 5319 16717
rect 5261 16708 5273 16711
rect 4764 16680 5273 16708
rect 4764 16668 4770 16680
rect 5261 16677 5273 16680
rect 5307 16677 5319 16711
rect 5994 16708 6000 16720
rect 5907 16680 6000 16708
rect 5261 16671 5319 16677
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 7834 16708 7840 16720
rect 7795 16680 7840 16708
rect 7834 16668 7840 16680
rect 7892 16668 7898 16720
rect 9214 16668 9220 16720
rect 9272 16708 9278 16720
rect 9876 16717 9904 16748
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 14090 16736 14096 16788
rect 14148 16776 14154 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 14148 16748 14381 16776
rect 14148 16736 14154 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 16666 16776 16672 16788
rect 16627 16748 16672 16776
rect 14369 16739 14427 16745
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 18601 16779 18659 16785
rect 18601 16776 18613 16779
rect 18196 16748 18613 16776
rect 18196 16736 18202 16748
rect 18601 16745 18613 16748
rect 18647 16776 18659 16779
rect 21082 16776 21088 16788
rect 18647 16748 19932 16776
rect 21043 16748 21088 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 9769 16711 9827 16717
rect 9769 16708 9781 16711
rect 9272 16680 9781 16708
rect 9272 16668 9278 16680
rect 9769 16677 9781 16680
rect 9815 16677 9827 16711
rect 9769 16671 9827 16677
rect 9861 16711 9919 16717
rect 9861 16677 9873 16711
rect 9907 16677 9919 16711
rect 11422 16708 11428 16720
rect 11383 16680 11428 16708
rect 9861 16671 9919 16677
rect 11422 16668 11428 16680
rect 11480 16668 11486 16720
rect 13535 16711 13593 16717
rect 13535 16677 13547 16711
rect 13581 16708 13593 16711
rect 13722 16708 13728 16720
rect 13581 16680 13728 16708
rect 13581 16677 13593 16680
rect 13535 16671 13593 16677
rect 13722 16668 13728 16680
rect 13780 16708 13786 16720
rect 14182 16708 14188 16720
rect 13780 16680 14188 16708
rect 13780 16668 13786 16680
rect 14182 16668 14188 16680
rect 14240 16668 14246 16720
rect 15286 16668 15292 16720
rect 15344 16708 15350 16720
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 15344 16680 15761 16708
rect 15344 16668 15350 16680
rect 15749 16677 15761 16680
rect 15795 16708 15807 16711
rect 15838 16708 15844 16720
rect 15795 16680 15844 16708
rect 15795 16677 15807 16680
rect 15749 16671 15807 16677
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 17494 16668 17500 16720
rect 17552 16708 17558 16720
rect 17773 16711 17831 16717
rect 17773 16708 17785 16711
rect 17552 16680 17785 16708
rect 17552 16668 17558 16680
rect 17773 16677 17785 16680
rect 17819 16677 17831 16711
rect 19334 16708 19340 16720
rect 19295 16680 19340 16708
rect 17773 16671 17831 16677
rect 19334 16668 19340 16680
rect 19392 16668 19398 16720
rect 19904 16717 19932 16748
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 19889 16711 19947 16717
rect 19889 16677 19901 16711
rect 19935 16708 19947 16711
rect 19978 16708 19984 16720
rect 19935 16680 19984 16708
rect 19935 16677 19947 16680
rect 19889 16671 19947 16677
rect 19978 16668 19984 16680
rect 20036 16668 20042 16720
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16640 2007 16643
rect 2590 16640 2596 16652
rect 1995 16612 2596 16640
rect 1995 16609 2007 16612
rect 1949 16603 2007 16609
rect 2590 16600 2596 16612
rect 2648 16600 2654 16652
rect 3028 16643 3086 16649
rect 3028 16609 3040 16643
rect 3074 16640 3086 16643
rect 3142 16640 3148 16652
rect 3074 16612 3148 16640
rect 3074 16609 3086 16612
rect 3028 16603 3086 16609
rect 3142 16600 3148 16612
rect 3200 16600 3206 16652
rect 4338 16600 4344 16652
rect 4396 16640 4402 16652
rect 20968 16643 21026 16649
rect 4396 16612 4844 16640
rect 4396 16600 4402 16612
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 4614 16572 4620 16584
rect 4111 16544 4620 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 4614 16532 4620 16544
rect 4672 16532 4678 16584
rect 4816 16572 4844 16612
rect 20968 16609 20980 16643
rect 21014 16640 21026 16643
rect 21082 16640 21088 16652
rect 21014 16612 21088 16640
rect 21014 16609 21026 16612
rect 20968 16603 21026 16609
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 21980 16643 22038 16649
rect 21980 16609 21992 16643
rect 22026 16640 22038 16643
rect 22094 16640 22100 16652
rect 22026 16612 22100 16640
rect 22026 16609 22038 16612
rect 21980 16603 22038 16609
rect 22094 16600 22100 16612
rect 22152 16600 22158 16652
rect 22922 16640 22928 16652
rect 22883 16612 22928 16640
rect 22922 16600 22928 16612
rect 22980 16600 22986 16652
rect 25016 16643 25074 16649
rect 25016 16609 25028 16643
rect 25062 16640 25074 16643
rect 25222 16640 25228 16652
rect 25062 16612 25228 16640
rect 25062 16609 25074 16612
rect 25016 16603 25074 16609
rect 25222 16600 25228 16612
rect 25280 16600 25286 16652
rect 5905 16575 5963 16581
rect 5905 16572 5917 16575
rect 4816 16544 5917 16572
rect 5905 16541 5917 16544
rect 5951 16572 5963 16575
rect 6178 16572 6184 16584
rect 5951 16544 6184 16572
rect 5951 16541 5963 16544
rect 5905 16535 5963 16541
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 7742 16572 7748 16584
rect 7703 16544 7748 16572
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 8662 16532 8668 16584
rect 8720 16572 8726 16584
rect 10045 16575 10103 16581
rect 10045 16572 10057 16575
rect 8720 16544 10057 16572
rect 8720 16532 8726 16544
rect 10045 16541 10057 16544
rect 10091 16572 10103 16575
rect 10870 16572 10876 16584
rect 10091 16544 10876 16572
rect 10091 16541 10103 16544
rect 10045 16535 10103 16541
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16572 11391 16575
rect 11606 16572 11612 16584
rect 11379 16544 11612 16572
rect 11379 16541 11391 16544
rect 11333 16535 11391 16541
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 13170 16572 13176 16584
rect 11756 16544 11801 16572
rect 13131 16544 13176 16572
rect 11756 16532 11762 16544
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 15105 16575 15163 16581
rect 15105 16541 15117 16575
rect 15151 16572 15163 16575
rect 15470 16572 15476 16584
rect 15151 16544 15476 16572
rect 15151 16541 15163 16544
rect 15105 16535 15163 16541
rect 15470 16532 15476 16544
rect 15528 16572 15534 16584
rect 15657 16575 15715 16581
rect 15657 16572 15669 16575
rect 15528 16544 15669 16572
rect 15528 16532 15534 16544
rect 15657 16541 15669 16544
rect 15703 16541 15715 16575
rect 15657 16535 15715 16541
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16572 17555 16575
rect 17678 16572 17684 16584
rect 17543 16544 17684 16572
rect 17543 16541 17555 16544
rect 17497 16535 17555 16541
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16572 18015 16575
rect 18782 16572 18788 16584
rect 18003 16544 18788 16572
rect 18003 16541 18015 16544
rect 17957 16535 18015 16541
rect 5350 16464 5356 16516
rect 5408 16504 5414 16516
rect 6457 16507 6515 16513
rect 6457 16504 6469 16507
rect 5408 16476 6469 16504
rect 5408 16464 5414 16476
rect 6457 16473 6469 16476
rect 6503 16504 6515 16507
rect 8110 16504 8116 16516
rect 6503 16476 8116 16504
rect 6503 16473 6515 16476
rect 6457 16467 6515 16473
rect 8110 16464 8116 16476
rect 8168 16464 8174 16516
rect 8294 16504 8300 16516
rect 8255 16476 8300 16504
rect 8294 16464 8300 16476
rect 8352 16464 8358 16516
rect 16209 16507 16267 16513
rect 16209 16473 16221 16507
rect 16255 16504 16267 16507
rect 17972 16504 18000 16535
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 19242 16572 19248 16584
rect 19203 16544 19248 16572
rect 19242 16532 19248 16544
rect 19300 16532 19306 16584
rect 22646 16532 22652 16584
rect 22704 16572 22710 16584
rect 23937 16575 23995 16581
rect 23937 16572 23949 16575
rect 22704 16544 23949 16572
rect 22704 16532 22710 16544
rect 23937 16541 23949 16544
rect 23983 16541 23995 16575
rect 23937 16535 23995 16541
rect 16255 16476 18000 16504
rect 22051 16507 22109 16513
rect 16255 16473 16267 16476
rect 16209 16467 16267 16473
rect 22051 16473 22063 16507
rect 22097 16504 22109 16507
rect 24670 16504 24676 16516
rect 22097 16476 24676 16504
rect 22097 16473 22109 16476
rect 22051 16467 22109 16473
rect 24670 16464 24676 16476
rect 24728 16464 24734 16516
rect 2130 16436 2136 16448
rect 2091 16408 2136 16436
rect 2130 16396 2136 16408
rect 2188 16396 2194 16448
rect 3099 16439 3157 16445
rect 3099 16405 3111 16439
rect 3145 16436 3157 16439
rect 7558 16436 7564 16448
rect 3145 16408 7564 16436
rect 3145 16405 3157 16408
rect 3099 16399 3157 16405
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 9030 16396 9036 16448
rect 9088 16436 9094 16448
rect 10870 16436 10876 16448
rect 9088 16408 10876 16436
rect 9088 16396 9094 16408
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11149 16439 11207 16445
rect 11149 16405 11161 16439
rect 11195 16436 11207 16439
rect 11238 16436 11244 16448
rect 11195 16408 11244 16436
rect 11195 16405 11207 16408
rect 11149 16399 11207 16405
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 11882 16396 11888 16448
rect 11940 16436 11946 16448
rect 12805 16439 12863 16445
rect 12805 16436 12817 16439
rect 11940 16408 12817 16436
rect 11940 16396 11946 16408
rect 12805 16405 12817 16408
rect 12851 16436 12863 16439
rect 13262 16436 13268 16448
rect 12851 16408 13268 16436
rect 12851 16405 12863 16408
rect 12805 16399 12863 16405
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 14090 16436 14096 16448
rect 14051 16408 14096 16436
rect 14090 16396 14096 16408
rect 14148 16396 14154 16448
rect 15286 16396 15292 16448
rect 15344 16436 15350 16448
rect 20622 16436 20628 16448
rect 15344 16408 20628 16436
rect 15344 16396 15350 16408
rect 20622 16396 20628 16408
rect 20680 16396 20686 16448
rect 22278 16396 22284 16448
rect 22336 16436 22342 16448
rect 23063 16439 23121 16445
rect 23063 16436 23075 16439
rect 22336 16408 23075 16436
rect 22336 16396 22342 16408
rect 23063 16405 23075 16408
rect 23109 16405 23121 16439
rect 23063 16399 23121 16405
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 25087 16439 25145 16445
rect 25087 16436 25099 16439
rect 24912 16408 25099 16436
rect 24912 16396 24918 16408
rect 25087 16405 25099 16408
rect 25133 16405 25145 16439
rect 25087 16399 25145 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 4798 16192 4804 16244
rect 4856 16232 4862 16244
rect 5077 16235 5135 16241
rect 5077 16232 5089 16235
rect 4856 16204 5089 16232
rect 4856 16192 4862 16204
rect 5077 16201 5089 16204
rect 5123 16201 5135 16235
rect 5077 16195 5135 16201
rect 5905 16235 5963 16241
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 5994 16232 6000 16244
rect 5951 16204 6000 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 6178 16232 6184 16244
rect 6139 16204 6184 16232
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 6641 16235 6699 16241
rect 6641 16201 6653 16235
rect 6687 16232 6699 16235
rect 6730 16232 6736 16244
rect 6687 16204 6736 16232
rect 6687 16201 6699 16204
rect 6641 16195 6699 16201
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 7193 16235 7251 16241
rect 7193 16201 7205 16235
rect 7239 16232 7251 16235
rect 7561 16235 7619 16241
rect 7561 16232 7573 16235
rect 7239 16204 7573 16232
rect 7239 16201 7251 16204
rect 7193 16195 7251 16201
rect 7561 16201 7573 16204
rect 7607 16232 7619 16235
rect 7834 16232 7840 16244
rect 7607 16204 7840 16232
rect 7607 16201 7619 16204
rect 7561 16195 7619 16201
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 9033 16235 9091 16241
rect 9033 16201 9045 16235
rect 9079 16232 9091 16235
rect 9490 16232 9496 16244
rect 9079 16204 9496 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 9674 16232 9680 16244
rect 9635 16204 9680 16232
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10778 16232 10784 16244
rect 10739 16204 10784 16232
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 14001 16235 14059 16241
rect 14001 16201 14013 16235
rect 14047 16232 14059 16235
rect 15657 16235 15715 16241
rect 15657 16232 15669 16235
rect 14047 16204 15669 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 15657 16201 15669 16204
rect 15703 16201 15715 16235
rect 15838 16232 15844 16244
rect 15799 16204 15844 16232
rect 15657 16195 15715 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 17494 16232 17500 16244
rect 16163 16204 17055 16232
rect 17455 16204 17500 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 9508 16164 9536 16192
rect 11241 16167 11299 16173
rect 11241 16164 11253 16167
rect 9508 16136 11253 16164
rect 11241 16133 11253 16136
rect 11287 16164 11299 16167
rect 11422 16164 11428 16176
rect 11287 16136 11428 16164
rect 11287 16133 11299 16136
rect 11241 16127 11299 16133
rect 11422 16124 11428 16136
rect 11480 16124 11486 16176
rect 15470 16164 15476 16176
rect 15431 16136 15476 16164
rect 15470 16124 15476 16136
rect 15528 16164 15534 16176
rect 17027 16164 17055 16204
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 19242 16192 19248 16244
rect 19300 16232 19306 16244
rect 20625 16235 20683 16241
rect 20625 16232 20637 16235
rect 19300 16204 20637 16232
rect 19300 16192 19306 16204
rect 20625 16201 20637 16204
rect 20671 16201 20683 16235
rect 21082 16232 21088 16244
rect 21043 16204 21088 16232
rect 20625 16195 20683 16201
rect 21082 16192 21088 16204
rect 21140 16192 21146 16244
rect 22002 16232 22008 16244
rect 21963 16204 22008 16232
rect 22002 16192 22008 16204
rect 22060 16192 22066 16244
rect 24762 16232 24768 16244
rect 24723 16204 24768 16232
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 17773 16167 17831 16173
rect 17773 16164 17785 16167
rect 15528 16136 16804 16164
rect 17027 16136 17785 16164
rect 15528 16124 15534 16136
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 6730 16096 6736 16108
rect 5592 16068 6736 16096
rect 5592 16056 5598 16068
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 7558 16056 7564 16108
rect 7616 16096 7622 16108
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7616 16068 7757 16096
rect 7616 16056 7622 16068
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 8389 16099 8447 16105
rect 8389 16065 8401 16099
rect 8435 16096 8447 16099
rect 8662 16096 8668 16108
rect 8435 16068 8668 16096
rect 8435 16065 8447 16068
rect 8389 16059 8447 16065
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 10778 16096 10784 16108
rect 9824 16068 10784 16096
rect 9824 16056 9830 16068
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16096 14795 16099
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14783 16068 14933 16096
rect 14783 16065 14795 16068
rect 14737 16059 14795 16065
rect 14921 16065 14933 16068
rect 14967 16096 14979 16099
rect 15286 16096 15292 16108
rect 14967 16068 15292 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15378 16056 15384 16108
rect 15436 16096 15442 16108
rect 16482 16096 16488 16108
rect 15436 16068 16488 16096
rect 15436 16056 15442 16068
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 16776 16105 16804 16136
rect 17773 16133 17785 16136
rect 17819 16133 17831 16167
rect 17773 16127 17831 16133
rect 16761 16099 16819 16105
rect 16761 16065 16773 16099
rect 16807 16065 16819 16099
rect 16761 16059 16819 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 2038 16028 2044 16040
rect 1443 16000 2044 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 16028 2559 16031
rect 2593 16031 2651 16037
rect 2593 16028 2605 16031
rect 2547 16000 2605 16028
rect 2547 15997 2559 16000
rect 2501 15991 2559 15997
rect 2593 15997 2605 16000
rect 2639 16028 2651 16031
rect 2866 16028 2872 16040
rect 2639 16000 2872 16028
rect 2639 15997 2651 16000
rect 2593 15991 2651 15997
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 16028 3111 16031
rect 3418 16028 3424 16040
rect 3099 16000 3424 16028
rect 3099 15997 3111 16000
rect 3053 15991 3111 15997
rect 2222 15920 2228 15972
rect 2280 15960 2286 15972
rect 3068 15960 3096 15991
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 4157 16031 4215 16037
rect 4157 15997 4169 16031
rect 4203 16028 4215 16031
rect 9861 16031 9919 16037
rect 4203 16000 5396 16028
rect 4203 15997 4215 16000
rect 4157 15991 4215 15997
rect 2280 15932 3096 15960
rect 3329 15963 3387 15969
rect 2280 15920 2286 15932
rect 3329 15929 3341 15963
rect 3375 15960 3387 15963
rect 5258 15960 5264 15972
rect 3375 15932 5264 15960
rect 3375 15929 3387 15932
rect 3329 15923 3387 15929
rect 5258 15920 5264 15932
rect 5316 15920 5322 15972
rect 5368 15904 5396 16000
rect 9861 15997 9873 16031
rect 9907 15997 9919 16031
rect 13078 16028 13084 16040
rect 13039 16000 13084 16028
rect 9861 15991 9919 15997
rect 7834 15920 7840 15972
rect 7892 15960 7898 15972
rect 7892 15932 7937 15960
rect 7892 15920 7898 15932
rect 8478 15920 8484 15972
rect 8536 15960 8542 15972
rect 9309 15963 9367 15969
rect 9309 15960 9321 15963
rect 8536 15932 9321 15960
rect 8536 15920 8542 15932
rect 9309 15929 9321 15932
rect 9355 15960 9367 15963
rect 9876 15960 9904 15991
rect 13078 15988 13084 16000
rect 13136 16028 13142 16040
rect 14277 16031 14335 16037
rect 14277 16028 14289 16031
rect 13136 16000 14289 16028
rect 13136 15988 13142 16000
rect 14277 15997 14289 16000
rect 14323 15997 14335 16031
rect 14277 15991 14335 15997
rect 15657 16031 15715 16037
rect 15657 15997 15669 16031
rect 15703 16028 15715 16031
rect 16209 16031 16267 16037
rect 16209 16028 16221 16031
rect 15703 16000 16221 16028
rect 15703 15997 15715 16000
rect 15657 15991 15715 15997
rect 16209 15997 16221 16000
rect 16255 15997 16267 16031
rect 16209 15991 16267 15997
rect 10182 15963 10240 15969
rect 10182 15960 10194 15963
rect 9355 15932 9904 15960
rect 10013 15932 10194 15960
rect 9355 15929 9367 15932
rect 9309 15923 9367 15929
rect 1210 15852 1216 15904
rect 1268 15892 1274 15904
rect 3142 15892 3148 15904
rect 1268 15864 3148 15892
rect 1268 15852 1274 15864
rect 3142 15852 3148 15864
rect 3200 15892 3206 15904
rect 3605 15895 3663 15901
rect 3605 15892 3617 15895
rect 3200 15864 3617 15892
rect 3200 15852 3206 15864
rect 3605 15861 3617 15864
rect 3651 15861 3663 15895
rect 3605 15855 3663 15861
rect 4065 15895 4123 15901
rect 4065 15861 4077 15895
rect 4111 15892 4123 15895
rect 4246 15892 4252 15904
rect 4111 15864 4252 15892
rect 4111 15861 4123 15864
rect 4065 15855 4123 15861
rect 4246 15852 4252 15864
rect 4304 15892 4310 15904
rect 4525 15895 4583 15901
rect 4525 15892 4537 15895
rect 4304 15864 4537 15892
rect 4304 15852 4310 15864
rect 4525 15861 4537 15864
rect 4571 15861 4583 15895
rect 5350 15892 5356 15904
rect 5311 15864 5356 15892
rect 4525 15855 4583 15861
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 10013 15892 10041 15932
rect 10182 15929 10194 15932
rect 10228 15960 10240 15963
rect 12161 15963 12219 15969
rect 12161 15960 12173 15963
rect 10228 15932 12173 15960
rect 10228 15929 10240 15932
rect 10182 15923 10240 15929
rect 12161 15929 12173 15932
rect 12207 15960 12219 15963
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 12207 15932 12909 15960
rect 12207 15929 12219 15932
rect 12161 15923 12219 15929
rect 12897 15929 12909 15932
rect 12943 15960 12955 15963
rect 12986 15960 12992 15972
rect 12943 15932 12992 15960
rect 12943 15929 12955 15932
rect 12897 15923 12955 15929
rect 12986 15920 12992 15932
rect 13044 15960 13050 15972
rect 13262 15960 13268 15972
rect 13044 15932 13268 15960
rect 13044 15920 13050 15932
rect 13262 15920 13268 15932
rect 13320 15960 13326 15972
rect 13402 15963 13460 15969
rect 13402 15960 13414 15963
rect 13320 15932 13414 15960
rect 13320 15920 13326 15932
rect 13402 15929 13414 15932
rect 13448 15960 13460 15963
rect 13722 15960 13728 15972
rect 13448 15932 13728 15960
rect 13448 15929 13460 15932
rect 13402 15923 13460 15929
rect 13722 15920 13728 15932
rect 13780 15920 13786 15972
rect 14090 15920 14096 15972
rect 14148 15960 14154 15972
rect 14918 15960 14924 15972
rect 14148 15932 14924 15960
rect 14148 15920 14154 15932
rect 14918 15920 14924 15932
rect 14976 15960 14982 15972
rect 15013 15963 15071 15969
rect 15013 15960 15025 15963
rect 14976 15932 15025 15960
rect 14976 15920 14982 15932
rect 15013 15929 15025 15932
rect 15059 15960 15071 15963
rect 16117 15963 16175 15969
rect 16117 15960 16129 15963
rect 15059 15932 16129 15960
rect 15059 15929 15071 15932
rect 15013 15923 15071 15929
rect 16117 15929 16129 15932
rect 16163 15929 16175 15963
rect 16224 15960 16252 15991
rect 16574 15960 16580 15972
rect 16224 15932 16580 15960
rect 16117 15923 16175 15929
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 17788 15960 17816 16127
rect 20070 16124 20076 16176
rect 20128 16164 20134 16176
rect 21315 16167 21373 16173
rect 21315 16164 21327 16167
rect 20128 16136 21327 16164
rect 20128 16124 20134 16136
rect 21315 16133 21327 16136
rect 21361 16133 21373 16167
rect 21315 16127 21373 16133
rect 18141 16099 18199 16105
rect 18141 16065 18153 16099
rect 18187 16096 18199 16099
rect 18598 16096 18604 16108
rect 18187 16068 18604 16096
rect 18187 16065 18199 16068
rect 18141 16059 18199 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19576 16068 19717 16096
rect 19576 16056 19582 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19978 16096 19984 16108
rect 19939 16068 19984 16096
rect 19705 16059 19763 16065
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 20162 16056 20168 16108
rect 20220 16096 20226 16108
rect 22327 16099 22385 16105
rect 22327 16096 22339 16099
rect 20220 16068 22339 16096
rect 20220 16056 20226 16068
rect 22327 16065 22339 16068
rect 22373 16065 22385 16099
rect 22327 16059 22385 16065
rect 21244 16031 21302 16037
rect 21244 15997 21256 16031
rect 21290 16028 21302 16031
rect 21290 16000 21772 16028
rect 21290 15997 21302 16000
rect 21244 15991 21302 15997
rect 18233 15963 18291 15969
rect 18233 15960 18245 15963
rect 17788 15932 18245 15960
rect 18233 15929 18245 15932
rect 18279 15929 18291 15963
rect 18782 15960 18788 15972
rect 18743 15932 18788 15960
rect 18233 15923 18291 15929
rect 11606 15892 11612 15904
rect 9732 15864 10041 15892
rect 11567 15864 11612 15892
rect 9732 15852 9738 15864
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 16298 15892 16304 15904
rect 15620 15864 16304 15892
rect 15620 15852 15626 15864
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 18248 15892 18276 15923
rect 18782 15920 18788 15932
rect 18840 15920 18846 15972
rect 19242 15920 19248 15972
rect 19300 15960 19306 15972
rect 19429 15963 19487 15969
rect 19429 15960 19441 15963
rect 19300 15932 19441 15960
rect 19300 15920 19306 15932
rect 19429 15929 19441 15932
rect 19475 15960 19487 15963
rect 19797 15963 19855 15969
rect 19797 15960 19809 15963
rect 19475 15932 19809 15960
rect 19475 15929 19487 15932
rect 19429 15923 19487 15929
rect 19797 15929 19809 15932
rect 19843 15929 19855 15963
rect 19797 15923 19855 15929
rect 19061 15895 19119 15901
rect 19061 15892 19073 15895
rect 18248 15864 19073 15892
rect 19061 15861 19073 15864
rect 19107 15892 19119 15895
rect 19334 15892 19340 15904
rect 19107 15864 19340 15892
rect 19107 15861 19119 15864
rect 19061 15855 19119 15861
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 21744 15901 21772 16000
rect 22002 15988 22008 16040
rect 22060 16028 22066 16040
rect 22224 16031 22282 16037
rect 22224 16028 22236 16031
rect 22060 16000 22236 16028
rect 22060 15988 22066 16000
rect 22224 15997 22236 16000
rect 22270 15997 22282 16031
rect 22224 15991 22282 15997
rect 22922 15988 22928 16040
rect 22980 16028 22986 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 22980 16000 24593 16028
rect 22980 15988 22986 16000
rect 24581 15997 24593 16000
rect 24627 16028 24639 16031
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24627 16000 25145 16028
rect 24627 15997 24639 16000
rect 24581 15991 24639 15997
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 21729 15895 21787 15901
rect 21729 15861 21741 15895
rect 21775 15892 21787 15895
rect 22186 15892 22192 15904
rect 21775 15864 22192 15892
rect 21775 15861 21787 15864
rect 21729 15855 21787 15861
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 22922 15892 22928 15904
rect 22883 15864 22928 15892
rect 22922 15852 22928 15864
rect 22980 15852 22986 15904
rect 25222 15852 25228 15904
rect 25280 15892 25286 15904
rect 25501 15895 25559 15901
rect 25501 15892 25513 15895
rect 25280 15864 25513 15892
rect 25280 15852 25286 15864
rect 25501 15861 25513 15864
rect 25547 15861 25559 15895
rect 25501 15855 25559 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1118 15648 1124 15700
rect 1176 15688 1182 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1176 15660 1593 15688
rect 1176 15648 1182 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 1581 15651 1639 15657
rect 2866 15648 2872 15700
rect 2924 15688 2930 15700
rect 3142 15688 3148 15700
rect 2924 15660 3148 15688
rect 2924 15648 2930 15660
rect 3142 15648 3148 15660
rect 3200 15648 3206 15700
rect 3510 15648 3516 15700
rect 3568 15688 3574 15700
rect 4614 15688 4620 15700
rect 3568 15660 4429 15688
rect 4575 15660 4620 15688
rect 3568 15648 3574 15660
rect 4246 15620 4252 15632
rect 4207 15592 4252 15620
rect 4246 15580 4252 15592
rect 4304 15580 4310 15632
rect 4401 15620 4429 15660
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 5074 15648 5080 15700
rect 5132 15688 5138 15700
rect 5534 15688 5540 15700
rect 5132 15660 5540 15688
rect 5132 15648 5138 15660
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 7469 15691 7527 15697
rect 7469 15657 7481 15691
rect 7515 15688 7527 15691
rect 7834 15688 7840 15700
rect 7515 15660 7840 15688
rect 7515 15657 7527 15660
rect 7469 15651 7527 15657
rect 7834 15648 7840 15660
rect 7892 15648 7898 15700
rect 9214 15648 9220 15700
rect 9272 15688 9278 15700
rect 9401 15691 9459 15697
rect 9401 15688 9413 15691
rect 9272 15660 9413 15688
rect 9272 15648 9278 15660
rect 9401 15657 9413 15660
rect 9447 15657 9459 15691
rect 9401 15651 9459 15657
rect 11514 15648 11520 15700
rect 11572 15688 11578 15700
rect 12529 15691 12587 15697
rect 12529 15688 12541 15691
rect 11572 15660 12541 15688
rect 11572 15648 11578 15660
rect 12529 15657 12541 15660
rect 12575 15688 12587 15691
rect 13170 15688 13176 15700
rect 12575 15660 13176 15688
rect 12575 15657 12587 15660
rect 12529 15651 12587 15657
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 13262 15648 13268 15700
rect 13320 15688 13326 15700
rect 13357 15691 13415 15697
rect 13357 15688 13369 15691
rect 13320 15660 13369 15688
rect 13320 15648 13326 15660
rect 13357 15657 13369 15660
rect 13403 15657 13415 15691
rect 14918 15688 14924 15700
rect 14879 15660 14924 15688
rect 13357 15651 13415 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 16482 15688 16488 15700
rect 16443 15660 16488 15688
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 18233 15691 18291 15697
rect 18233 15657 18245 15691
rect 18279 15688 18291 15691
rect 18322 15688 18328 15700
rect 18279 15660 18328 15688
rect 18279 15657 18291 15660
rect 18233 15651 18291 15657
rect 18322 15648 18328 15660
rect 18380 15648 18386 15700
rect 18598 15688 18604 15700
rect 18559 15660 18604 15688
rect 18598 15648 18604 15660
rect 18656 15648 18662 15700
rect 19518 15648 19524 15700
rect 19576 15688 19582 15700
rect 19705 15691 19763 15697
rect 19705 15688 19717 15691
rect 19576 15660 19717 15688
rect 19576 15648 19582 15660
rect 19705 15657 19717 15660
rect 19751 15657 19763 15691
rect 19705 15651 19763 15657
rect 20806 15648 20812 15700
rect 20864 15688 20870 15700
rect 22002 15688 22008 15700
rect 20864 15660 22008 15688
rect 20864 15648 20870 15660
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 23842 15648 23848 15700
rect 23900 15688 23906 15700
rect 24811 15691 24869 15697
rect 24811 15688 24823 15691
rect 23900 15660 24823 15688
rect 23900 15648 23906 15660
rect 24811 15657 24823 15660
rect 24857 15657 24869 15691
rect 24811 15651 24869 15657
rect 6178 15620 6184 15632
rect 4401 15592 6184 15620
rect 6178 15580 6184 15592
rect 6236 15580 6242 15632
rect 6911 15623 6969 15629
rect 6911 15589 6923 15623
rect 6957 15620 6969 15623
rect 7006 15620 7012 15632
rect 6957 15592 7012 15620
rect 6957 15589 6969 15592
rect 6911 15583 6969 15589
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 7558 15580 7564 15632
rect 7616 15620 7622 15632
rect 8113 15623 8171 15629
rect 8113 15620 8125 15623
rect 7616 15592 8125 15620
rect 7616 15580 7622 15592
rect 8113 15589 8125 15592
rect 8159 15589 8171 15623
rect 8113 15583 8171 15589
rect 8711 15623 8769 15629
rect 8711 15589 8723 15623
rect 8757 15620 8769 15623
rect 11606 15620 11612 15632
rect 8757 15592 11612 15620
rect 8757 15589 8769 15592
rect 8711 15583 8769 15589
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 12161 15623 12219 15629
rect 12161 15589 12173 15623
rect 12207 15620 12219 15623
rect 13078 15620 13084 15632
rect 12207 15592 13084 15620
rect 12207 15589 12219 15592
rect 12161 15583 12219 15589
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 14734 15580 14740 15632
rect 14792 15620 14798 15632
rect 15473 15623 15531 15629
rect 15473 15620 15485 15623
rect 14792 15592 15485 15620
rect 14792 15580 14798 15592
rect 15473 15589 15485 15592
rect 15519 15589 15531 15623
rect 17310 15620 17316 15632
rect 17271 15592 17316 15620
rect 15473 15583 15531 15589
rect 17310 15580 17316 15592
rect 17368 15580 17374 15632
rect 17678 15580 17684 15632
rect 17736 15620 17742 15632
rect 17865 15623 17923 15629
rect 17865 15620 17877 15623
rect 17736 15592 17877 15620
rect 17736 15580 17742 15592
rect 17865 15589 17877 15592
rect 17911 15620 17923 15623
rect 18782 15620 18788 15632
rect 17911 15592 18788 15620
rect 17911 15589 17923 15592
rect 17865 15583 17923 15589
rect 18782 15580 18788 15592
rect 18840 15580 18846 15632
rect 18877 15623 18935 15629
rect 18877 15589 18889 15623
rect 18923 15620 18935 15623
rect 18966 15620 18972 15632
rect 18923 15592 18972 15620
rect 18923 15589 18935 15592
rect 18877 15583 18935 15589
rect 18966 15580 18972 15592
rect 19024 15580 19030 15632
rect 19429 15623 19487 15629
rect 19429 15589 19441 15623
rect 19475 15620 19487 15623
rect 19978 15620 19984 15632
rect 19475 15592 19984 15620
rect 19475 15589 19487 15592
rect 19429 15583 19487 15589
rect 19978 15580 19984 15592
rect 20036 15580 20042 15632
rect 21266 15620 21272 15632
rect 21227 15592 21272 15620
rect 21266 15580 21272 15592
rect 21324 15580 21330 15632
rect 21450 15580 21456 15632
rect 21508 15620 21514 15632
rect 21508 15592 23474 15620
rect 21508 15580 21514 15592
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 2961 15555 3019 15561
rect 2961 15521 2973 15555
rect 3007 15552 3019 15555
rect 3418 15552 3424 15564
rect 3007 15524 3424 15552
rect 3007 15521 3019 15524
rect 2961 15515 3019 15521
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 5074 15552 5080 15564
rect 5035 15524 5080 15552
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 5534 15552 5540 15564
rect 5495 15524 5540 15552
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 8478 15552 8484 15564
rect 5767 15524 8484 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 8478 15512 8484 15524
rect 8536 15512 8542 15564
rect 8570 15512 8576 15564
rect 8628 15552 8634 15564
rect 9861 15555 9919 15561
rect 8628 15524 8673 15552
rect 8628 15512 8634 15524
rect 9861 15521 9873 15555
rect 9907 15521 9919 15555
rect 9861 15515 9919 15521
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15484 2099 15487
rect 2590 15484 2596 15496
rect 2087 15456 2596 15484
rect 2087 15453 2099 15456
rect 2041 15447 2099 15453
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 5258 15444 5264 15496
rect 5316 15484 5322 15496
rect 6549 15487 6607 15493
rect 6549 15484 6561 15487
rect 5316 15456 6561 15484
rect 5316 15444 5322 15456
rect 6549 15453 6561 15456
rect 6595 15484 6607 15487
rect 8018 15484 8024 15496
rect 6595 15456 8024 15484
rect 6595 15453 6607 15456
rect 6549 15447 6607 15453
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 9870 15428 9898 15515
rect 10134 15512 10140 15564
rect 10192 15552 10198 15564
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 10192 15524 10333 15552
rect 10192 15512 10198 15524
rect 10321 15521 10333 15524
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 10870 15512 10876 15564
rect 10928 15552 10934 15564
rect 11422 15552 11428 15564
rect 10928 15524 11428 15552
rect 10928 15512 10934 15524
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 11882 15552 11888 15564
rect 11843 15524 11888 15552
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 22716 15555 22774 15561
rect 22716 15521 22728 15555
rect 22762 15552 22774 15555
rect 22922 15552 22928 15564
rect 22762 15524 22928 15552
rect 22762 15521 22774 15524
rect 22716 15515 22774 15521
rect 22922 15512 22928 15524
rect 22980 15512 22986 15564
rect 23446 15552 23474 15592
rect 23728 15555 23786 15561
rect 23728 15552 23740 15555
rect 23446 15524 23740 15552
rect 23728 15521 23740 15524
rect 23774 15552 23786 15555
rect 24210 15552 24216 15564
rect 23774 15524 24216 15552
rect 23774 15521 23786 15524
rect 23728 15515 23786 15521
rect 24210 15512 24216 15524
rect 24268 15512 24274 15564
rect 24740 15555 24798 15561
rect 24740 15521 24752 15555
rect 24786 15552 24798 15555
rect 25130 15552 25136 15564
rect 24786 15524 25136 15552
rect 24786 15521 24798 15524
rect 24740 15515 24798 15521
rect 25130 15512 25136 15524
rect 25188 15512 25194 15564
rect 10597 15487 10655 15493
rect 10597 15453 10609 15487
rect 10643 15484 10655 15487
rect 12342 15484 12348 15496
rect 10643 15456 12348 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 12989 15487 13047 15493
rect 12989 15484 13001 15487
rect 12820 15456 13001 15484
rect 9858 15416 9864 15428
rect 2608 15388 9864 15416
rect 2222 15308 2228 15360
rect 2280 15348 2286 15360
rect 2608 15357 2636 15388
rect 9858 15376 9864 15388
rect 9916 15376 9922 15428
rect 2593 15351 2651 15357
rect 2593 15348 2605 15351
rect 2280 15320 2605 15348
rect 2280 15308 2286 15320
rect 2593 15317 2605 15320
rect 2639 15317 2651 15351
rect 2593 15311 2651 15317
rect 3697 15351 3755 15357
rect 3697 15317 3709 15351
rect 3743 15348 3755 15351
rect 4062 15348 4068 15360
rect 3743 15320 4068 15348
rect 3743 15317 3755 15320
rect 3697 15311 3755 15317
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 6362 15348 6368 15360
rect 6323 15320 6368 15348
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 7834 15348 7840 15360
rect 7795 15320 7840 15348
rect 7834 15308 7840 15320
rect 7892 15308 7898 15360
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 12820 15357 12848 15456
rect 12989 15453 13001 15456
rect 13035 15453 13047 15487
rect 15378 15484 15384 15496
rect 15339 15456 15384 15484
rect 12989 15447 13047 15453
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 15470 15444 15476 15496
rect 15528 15484 15534 15496
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15528 15456 15669 15484
rect 15528 15444 15534 15456
rect 15657 15453 15669 15456
rect 15703 15453 15715 15487
rect 17210 15487 17268 15493
rect 17210 15484 17222 15487
rect 15657 15447 15715 15453
rect 17144 15456 17222 15484
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 12676 15320 12817 15348
rect 12676 15308 12682 15320
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 12805 15311 12863 15317
rect 13909 15351 13967 15357
rect 13909 15317 13921 15351
rect 13955 15348 13967 15351
rect 14734 15348 14740 15360
rect 13955 15320 14740 15348
rect 13955 15317 13967 15320
rect 13909 15311 13967 15317
rect 14734 15308 14740 15320
rect 14792 15308 14798 15360
rect 17144 15348 17172 15456
rect 17210 15453 17222 15456
rect 17256 15453 17268 15487
rect 17210 15447 17268 15453
rect 18598 15444 18604 15496
rect 18656 15484 18662 15496
rect 18785 15487 18843 15493
rect 18785 15484 18797 15487
rect 18656 15456 18797 15484
rect 18656 15444 18662 15456
rect 18785 15453 18797 15456
rect 18831 15453 18843 15487
rect 21174 15484 21180 15496
rect 21135 15456 21180 15484
rect 18785 15447 18843 15453
rect 21174 15444 21180 15456
rect 21232 15444 21238 15496
rect 21453 15487 21511 15493
rect 21453 15453 21465 15487
rect 21499 15453 21511 15487
rect 22094 15484 22100 15496
rect 22055 15456 22100 15484
rect 21453 15447 21511 15453
rect 20162 15416 20168 15428
rect 17328 15388 20168 15416
rect 17218 15348 17224 15360
rect 17131 15320 17224 15348
rect 17218 15308 17224 15320
rect 17276 15348 17282 15360
rect 17328 15348 17356 15388
rect 20162 15376 20168 15388
rect 20220 15376 20226 15428
rect 21082 15376 21088 15428
rect 21140 15416 21146 15428
rect 21468 15416 21496 15447
rect 22094 15444 22100 15456
rect 22152 15444 22158 15496
rect 21634 15416 21640 15428
rect 21140 15388 21640 15416
rect 21140 15376 21146 15388
rect 21634 15376 21640 15388
rect 21692 15376 21698 15428
rect 22787 15419 22845 15425
rect 22787 15416 22799 15419
rect 21744 15388 22799 15416
rect 17276 15320 17356 15348
rect 17276 15308 17282 15320
rect 17494 15308 17500 15360
rect 17552 15348 17558 15360
rect 21744 15348 21772 15388
rect 22787 15385 22799 15388
rect 22833 15385 22845 15419
rect 22787 15379 22845 15385
rect 17552 15320 21772 15348
rect 17552 15308 17558 15320
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 23799 15351 23857 15357
rect 23799 15348 23811 15351
rect 21968 15320 23811 15348
rect 21968 15308 21974 15320
rect 23799 15317 23811 15320
rect 23845 15317 23857 15351
rect 23799 15311 23857 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2130 15144 2136 15156
rect 2091 15116 2136 15144
rect 2130 15104 2136 15116
rect 2188 15104 2194 15156
rect 3050 15144 3056 15156
rect 3011 15116 3056 15144
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 3418 15144 3424 15156
rect 3379 15116 3424 15144
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4890 15144 4896 15156
rect 4755 15116 4896 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 6181 15147 6239 15153
rect 6181 15113 6193 15147
rect 6227 15144 6239 15147
rect 6457 15147 6515 15153
rect 6457 15144 6469 15147
rect 6227 15116 6469 15144
rect 6227 15113 6239 15116
rect 6181 15107 6239 15113
rect 6457 15113 6469 15116
rect 6503 15144 6515 15147
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 6503 15116 6561 15144
rect 6503 15113 6515 15116
rect 6457 15107 6515 15113
rect 6549 15113 6561 15116
rect 6595 15113 6607 15147
rect 6549 15107 6607 15113
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 8018 15144 8024 15156
rect 7156 15116 7788 15144
rect 7979 15116 8024 15144
rect 7156 15104 7162 15116
rect 1394 15036 1400 15088
rect 1452 15076 1458 15088
rect 2409 15079 2467 15085
rect 2409 15076 2421 15079
rect 1452 15048 2421 15076
rect 1452 15036 1458 15048
rect 2409 15045 2421 15048
rect 2455 15045 2467 15079
rect 2409 15039 2467 15045
rect 2731 15079 2789 15085
rect 2731 15045 2743 15079
rect 2777 15076 2789 15079
rect 7558 15076 7564 15088
rect 2777 15048 7564 15076
rect 2777 15045 2789 15048
rect 2731 15039 2789 15045
rect 7558 15036 7564 15048
rect 7616 15036 7622 15088
rect 7760 15076 7788 15116
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 9858 15144 9864 15156
rect 9819 15116 9864 15144
rect 9858 15104 9864 15116
rect 9916 15144 9922 15156
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 9916 15116 10609 15144
rect 9916 15104 9922 15116
rect 10597 15113 10609 15116
rect 10643 15144 10655 15147
rect 10962 15144 10968 15156
rect 10643 15116 10968 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 9674 15076 9680 15088
rect 7760 15048 9680 15076
rect 9674 15036 9680 15048
rect 9732 15036 9738 15088
rect 10134 15036 10140 15088
rect 10192 15076 10198 15088
rect 10229 15079 10287 15085
rect 10229 15076 10241 15079
rect 10192 15048 10241 15076
rect 10192 15036 10198 15048
rect 10229 15045 10241 15048
rect 10275 15045 10287 15079
rect 10229 15039 10287 15045
rect 4341 15011 4399 15017
rect 3620 14980 4292 15008
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14940 1639 14943
rect 2130 14940 2136 14952
rect 1627 14912 2136 14940
rect 1627 14909 1639 14912
rect 1581 14903 1639 14909
rect 2130 14900 2136 14912
rect 2188 14900 2194 14952
rect 2660 14943 2718 14949
rect 2660 14909 2672 14943
rect 2706 14940 2718 14943
rect 3050 14940 3056 14952
rect 2706 14912 3056 14940
rect 2706 14909 2718 14912
rect 2660 14903 2718 14909
rect 3050 14900 3056 14912
rect 3108 14900 3114 14952
rect 3142 14900 3148 14952
rect 3200 14940 3206 14952
rect 3510 14940 3516 14952
rect 3200 14912 3516 14940
rect 3200 14900 3206 14912
rect 3510 14900 3516 14912
rect 3568 14940 3574 14952
rect 3620 14949 3648 14980
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3568 14912 3617 14940
rect 3568 14900 3574 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 4062 14940 4068 14952
rect 4023 14912 4068 14940
rect 3605 14903 3663 14909
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4264 14940 4292 14980
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 4614 15008 4620 15020
rect 4387 14980 4620 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 4614 14968 4620 14980
rect 4672 14968 4678 15020
rect 4890 14968 4896 15020
rect 4948 15008 4954 15020
rect 5905 15011 5963 15017
rect 4948 14980 5672 15008
rect 4948 14968 4954 14980
rect 5166 14940 5172 14952
rect 4264 14912 5172 14940
rect 5166 14900 5172 14912
rect 5224 14900 5230 14952
rect 5644 14949 5672 14980
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 6362 15008 6368 15020
rect 5951 14980 6368 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6362 14968 6368 14980
rect 6420 15008 6426 15020
rect 6825 15011 6883 15017
rect 6825 15008 6837 15011
rect 6420 14980 6837 15008
rect 6420 14968 6426 14980
rect 6825 14977 6837 14980
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 8662 14968 8668 15020
rect 8720 15008 8726 15020
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8720 14980 8953 15008
rect 8720 14968 8726 14980
rect 8941 14977 8953 14980
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 5629 14943 5687 14949
rect 5629 14909 5641 14943
rect 5675 14940 5687 14943
rect 8018 14940 8024 14952
rect 5675 14912 8024 14940
rect 5675 14909 5687 14912
rect 5629 14903 5687 14909
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 10612 14940 10640 15107
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 12575 15147 12633 15153
rect 12575 15144 12587 15147
rect 11296 15116 12587 15144
rect 11296 15104 11302 15116
rect 12575 15113 12587 15116
rect 12621 15113 12633 15147
rect 12575 15107 12633 15113
rect 12986 15104 12992 15156
rect 13044 15144 13050 15156
rect 13265 15147 13323 15153
rect 13265 15144 13277 15147
rect 13044 15116 13277 15144
rect 13044 15104 13050 15116
rect 13265 15113 13277 15116
rect 13311 15113 13323 15147
rect 14734 15144 14740 15156
rect 14695 15116 14740 15144
rect 13265 15107 13323 15113
rect 14734 15104 14740 15116
rect 14792 15144 14798 15156
rect 16761 15147 16819 15153
rect 16761 15144 16773 15147
rect 14792 15116 16773 15144
rect 14792 15104 14798 15116
rect 16761 15113 16773 15116
rect 16807 15144 16819 15147
rect 17310 15144 17316 15156
rect 16807 15116 17316 15144
rect 16807 15113 16819 15116
rect 16761 15107 16819 15113
rect 17310 15104 17316 15116
rect 17368 15144 17374 15156
rect 18966 15144 18972 15156
rect 17368 15116 18972 15144
rect 17368 15104 17374 15116
rect 18966 15104 18972 15116
rect 19024 15144 19030 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 19024 15116 19073 15144
rect 19024 15104 19030 15116
rect 19061 15113 19073 15116
rect 19107 15113 19119 15147
rect 19061 15107 19119 15113
rect 21266 15104 21272 15156
rect 21324 15144 21330 15156
rect 21453 15147 21511 15153
rect 21453 15144 21465 15147
rect 21324 15116 21465 15144
rect 21324 15104 21330 15116
rect 21453 15113 21465 15116
rect 21499 15144 21511 15147
rect 22097 15147 22155 15153
rect 22097 15144 22109 15147
rect 21499 15116 22109 15144
rect 21499 15113 21511 15116
rect 21453 15107 21511 15113
rect 22097 15113 22109 15116
rect 22143 15113 22155 15147
rect 22097 15107 22155 15113
rect 22833 15147 22891 15153
rect 22833 15113 22845 15147
rect 22879 15144 22891 15147
rect 22922 15144 22928 15156
rect 22879 15116 22928 15144
rect 22879 15113 22891 15116
rect 22833 15107 22891 15113
rect 22922 15104 22928 15116
rect 22980 15104 22986 15156
rect 23106 15144 23112 15156
rect 23067 15116 23112 15144
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 25130 15144 25136 15156
rect 25091 15116 25136 15144
rect 25130 15104 25136 15116
rect 25188 15104 25194 15156
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 11793 15079 11851 15085
rect 11793 15076 11805 15079
rect 11480 15048 11805 15076
rect 11480 15036 11486 15048
rect 11793 15045 11805 15048
rect 11839 15045 11851 15079
rect 11793 15039 11851 15045
rect 17126 15036 17132 15088
rect 17184 15076 17190 15088
rect 18598 15076 18604 15088
rect 17184 15048 18604 15076
rect 17184 15036 17190 15048
rect 18598 15036 18604 15048
rect 18656 15076 18662 15088
rect 19429 15079 19487 15085
rect 19429 15076 19441 15079
rect 18656 15048 19441 15076
rect 18656 15036 18662 15048
rect 19429 15045 19441 15048
rect 19475 15045 19487 15079
rect 19429 15039 19487 15045
rect 21174 15036 21180 15088
rect 21232 15076 21238 15088
rect 21729 15079 21787 15085
rect 21729 15076 21741 15079
rect 21232 15048 21741 15076
rect 21232 15036 21238 15048
rect 21729 15045 21741 15048
rect 21775 15045 21787 15079
rect 21729 15039 21787 15045
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 11514 15008 11520 15020
rect 10744 14980 11284 15008
rect 11475 14980 11520 15008
rect 10744 14968 10750 14980
rect 11256 14949 11284 14980
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 13814 15008 13820 15020
rect 13775 14980 13820 15008
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14090 15008 14096 15020
rect 14051 14980 14096 15008
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 15838 15008 15844 15020
rect 15799 14980 15844 15008
rect 15838 14968 15844 14980
rect 15896 14968 15902 15020
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 16632 14980 17785 15008
rect 16632 14968 16638 14980
rect 17773 14977 17785 14980
rect 17819 14977 17831 15011
rect 17773 14971 17831 14977
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 15008 18199 15011
rect 18322 15008 18328 15020
rect 18187 14980 18328 15008
rect 18187 14977 18199 14980
rect 18141 14971 18199 14977
rect 10781 14943 10839 14949
rect 10781 14940 10793 14943
rect 10612 14912 10793 14940
rect 10781 14909 10793 14912
rect 10827 14909 10839 14943
rect 10781 14903 10839 14909
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 11882 14940 11888 14952
rect 11287 14912 11888 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 11882 14900 11888 14912
rect 11940 14940 11946 14952
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 11940 14912 12173 14940
rect 11940 14900 11946 14912
rect 12161 14909 12173 14912
rect 12207 14909 12219 14943
rect 12161 14903 12219 14909
rect 12504 14943 12562 14949
rect 12504 14909 12516 14943
rect 12550 14940 12562 14943
rect 12894 14940 12900 14952
rect 12550 14912 12900 14940
rect 12550 14909 12562 14912
rect 12504 14903 12562 14909
rect 12894 14900 12900 14912
rect 12952 14940 12958 14952
rect 12952 14912 13032 14940
rect 12952 14900 12958 14912
rect 2774 14872 2780 14884
rect 1964 14844 2780 14872
rect 1765 14807 1823 14813
rect 1765 14773 1777 14807
rect 1811 14804 1823 14807
rect 1964 14804 1992 14844
rect 2774 14832 2780 14844
rect 2832 14832 2838 14884
rect 3418 14832 3424 14884
rect 3476 14872 3482 14884
rect 6457 14875 6515 14881
rect 3476 14844 5120 14872
rect 3476 14832 3482 14844
rect 5092 14816 5120 14844
rect 6457 14841 6469 14875
rect 6503 14872 6515 14875
rect 6822 14872 6828 14884
rect 6503 14844 6828 14872
rect 6503 14841 6515 14844
rect 6457 14835 6515 14841
rect 6822 14832 6828 14844
rect 6880 14872 6886 14884
rect 7146 14875 7204 14881
rect 7146 14872 7158 14875
rect 6880 14844 7158 14872
rect 6880 14832 6886 14844
rect 7146 14841 7158 14844
rect 7192 14841 7204 14875
rect 8662 14872 8668 14884
rect 8623 14844 8668 14872
rect 7146 14835 7204 14841
rect 8662 14832 8668 14844
rect 8720 14832 8726 14884
rect 8754 14832 8760 14884
rect 8812 14872 8818 14884
rect 8812 14844 8857 14872
rect 8812 14832 8818 14844
rect 1811 14776 1992 14804
rect 1811 14773 1823 14776
rect 1765 14767 1823 14773
rect 3878 14764 3884 14816
rect 3936 14804 3942 14816
rect 4154 14804 4160 14816
rect 3936 14776 4160 14804
rect 3936 14764 3942 14776
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 5074 14804 5080 14816
rect 4987 14776 5080 14804
rect 5074 14764 5080 14776
rect 5132 14804 5138 14816
rect 5258 14804 5264 14816
rect 5132 14776 5264 14804
rect 5132 14764 5138 14776
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 7742 14804 7748 14816
rect 7703 14776 7748 14804
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 8570 14804 8576 14816
rect 8527 14776 8576 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 8570 14764 8576 14776
rect 8628 14764 8634 14816
rect 13004 14813 13032 14912
rect 16482 14900 16488 14952
rect 16540 14940 16546 14952
rect 17012 14943 17070 14949
rect 17012 14940 17024 14943
rect 16540 14912 17024 14940
rect 16540 14900 16546 14912
rect 17012 14909 17024 14912
rect 17058 14940 17070 14943
rect 17058 14912 17540 14940
rect 17058 14909 17070 14912
rect 17012 14903 17070 14909
rect 13909 14875 13967 14881
rect 13909 14841 13921 14875
rect 13955 14872 13967 14875
rect 14182 14872 14188 14884
rect 13955 14844 14188 14872
rect 13955 14841 13967 14844
rect 13909 14835 13967 14841
rect 14182 14832 14188 14844
rect 14240 14832 14246 14884
rect 15381 14875 15439 14881
rect 15381 14841 15393 14875
rect 15427 14841 15439 14875
rect 15381 14835 15439 14841
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14804 13047 14807
rect 13170 14804 13176 14816
rect 13035 14776 13176 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 15197 14807 15255 14813
rect 15197 14773 15209 14807
rect 15243 14804 15255 14807
rect 15286 14804 15292 14816
rect 15243 14776 15292 14804
rect 15243 14773 15255 14776
rect 15197 14767 15255 14773
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 15396 14804 15424 14835
rect 15470 14832 15476 14884
rect 15528 14872 15534 14884
rect 15528 14844 15573 14872
rect 15528 14832 15534 14844
rect 16390 14804 16396 14816
rect 15396 14776 16396 14804
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 17083 14807 17141 14813
rect 17083 14773 17095 14807
rect 17129 14804 17141 14807
rect 17310 14804 17316 14816
rect 17129 14776 17316 14804
rect 17129 14773 17141 14776
rect 17083 14767 17141 14773
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 17512 14813 17540 14912
rect 17788 14872 17816 14971
rect 18322 14968 18328 14980
rect 18380 14968 18386 15020
rect 18782 15008 18788 15020
rect 18743 14980 18788 15008
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 20162 14968 20168 15020
rect 20220 15008 20226 15020
rect 22462 15008 22468 15020
rect 20220 14980 22468 15008
rect 20220 14968 20226 14980
rect 22462 14968 22468 14980
rect 22520 14968 22526 15020
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 20349 14943 20407 14949
rect 20349 14940 20361 14943
rect 19484 14912 20361 14940
rect 19484 14900 19490 14912
rect 20349 14909 20361 14912
rect 20395 14909 20407 14943
rect 20530 14940 20536 14952
rect 20491 14912 20536 14940
rect 20349 14903 20407 14909
rect 18233 14875 18291 14881
rect 18233 14872 18245 14875
rect 17788 14844 18245 14872
rect 18233 14841 18245 14844
rect 18279 14872 18291 14875
rect 19242 14872 19248 14884
rect 18279 14844 19248 14872
rect 18279 14841 18291 14844
rect 18233 14835 18291 14841
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 20364 14872 20392 14903
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 20714 14900 20720 14952
rect 20772 14940 20778 14952
rect 22348 14943 22406 14949
rect 22348 14940 22360 14943
rect 20772 14912 22360 14940
rect 20772 14900 20778 14912
rect 22348 14909 22360 14912
rect 22394 14940 22406 14943
rect 23106 14940 23112 14952
rect 22394 14912 23112 14940
rect 22394 14909 22406 14912
rect 22348 14903 22406 14909
rect 23106 14900 23112 14912
rect 23164 14900 23170 14952
rect 23728 14943 23786 14949
rect 23728 14940 23740 14943
rect 23446 14912 23740 14940
rect 20854 14875 20912 14881
rect 20854 14872 20866 14875
rect 20364 14844 20866 14872
rect 20854 14841 20866 14844
rect 20900 14841 20912 14875
rect 20854 14835 20912 14841
rect 21174 14832 21180 14884
rect 21232 14872 21238 14884
rect 23446 14872 23474 14912
rect 23728 14909 23740 14912
rect 23774 14940 23786 14943
rect 24121 14943 24179 14949
rect 24121 14940 24133 14943
rect 23774 14912 24133 14940
rect 23774 14909 23786 14912
rect 23728 14903 23786 14909
rect 24121 14909 24133 14912
rect 24167 14909 24179 14943
rect 24121 14903 24179 14909
rect 21232 14844 23474 14872
rect 21232 14832 21238 14844
rect 24026 14832 24032 14884
rect 24084 14872 24090 14884
rect 24673 14875 24731 14881
rect 24673 14872 24685 14875
rect 24084 14844 24685 14872
rect 24084 14832 24090 14844
rect 24673 14841 24685 14844
rect 24719 14841 24731 14875
rect 24673 14835 24731 14841
rect 17497 14807 17555 14813
rect 17497 14773 17509 14807
rect 17543 14804 17555 14807
rect 18506 14804 18512 14816
rect 17543 14776 18512 14804
rect 17543 14773 17555 14776
rect 17497 14767 17555 14773
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 20990 14764 20996 14816
rect 21048 14804 21054 14816
rect 22419 14807 22477 14813
rect 22419 14804 22431 14807
rect 21048 14776 22431 14804
rect 21048 14764 21054 14776
rect 22419 14773 22431 14776
rect 22465 14773 22477 14807
rect 22419 14767 22477 14773
rect 23198 14764 23204 14816
rect 23256 14804 23262 14816
rect 23799 14807 23857 14813
rect 23799 14804 23811 14807
rect 23256 14776 23811 14804
rect 23256 14764 23262 14776
rect 23799 14773 23811 14776
rect 23845 14773 23857 14807
rect 23799 14767 23857 14773
rect 24210 14764 24216 14816
rect 24268 14804 24274 14816
rect 24489 14807 24547 14813
rect 24489 14804 24501 14807
rect 24268 14776 24501 14804
rect 24268 14764 24274 14776
rect 24489 14773 24501 14776
rect 24535 14773 24547 14807
rect 24489 14767 24547 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 3418 14600 3424 14612
rect 2740 14572 3424 14600
rect 2740 14560 2746 14572
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 3510 14560 3516 14612
rect 3568 14600 3574 14612
rect 3605 14603 3663 14609
rect 3605 14600 3617 14603
rect 3568 14572 3617 14600
rect 3568 14560 3574 14572
rect 3605 14569 3617 14572
rect 3651 14569 3663 14603
rect 3605 14563 3663 14569
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 8662 14600 8668 14612
rect 4212 14572 4257 14600
rect 4448 14572 8668 14600
rect 4212 14560 4218 14572
rect 3099 14535 3157 14541
rect 3099 14501 3111 14535
rect 3145 14532 3157 14535
rect 4448 14532 4476 14572
rect 8662 14560 8668 14572
rect 8720 14600 8726 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 8720 14572 8953 14600
rect 8720 14560 8726 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 8941 14563 8999 14569
rect 10686 14560 10692 14612
rect 10744 14600 10750 14612
rect 10781 14603 10839 14609
rect 10781 14600 10793 14603
rect 10744 14572 10793 14600
rect 10744 14560 10750 14572
rect 10781 14569 10793 14572
rect 10827 14569 10839 14603
rect 13814 14600 13820 14612
rect 13775 14572 13820 14600
rect 10781 14563 10839 14569
rect 7742 14532 7748 14544
rect 3145 14504 4476 14532
rect 4540 14504 6316 14532
rect 7703 14504 7748 14532
rect 3145 14501 3157 14504
rect 3099 14495 3157 14501
rect 4540 14476 4568 14504
rect 6288 14476 6316 14504
rect 7742 14492 7748 14504
rect 7800 14532 7806 14544
rect 8110 14532 8116 14544
rect 7800 14504 8116 14532
rect 7800 14492 7806 14504
rect 8110 14492 8116 14504
rect 8168 14532 8174 14544
rect 8573 14535 8631 14541
rect 8573 14532 8585 14535
rect 8168 14504 8585 14532
rect 8168 14492 8174 14504
rect 8573 14501 8585 14504
rect 8619 14532 8631 14535
rect 8754 14532 8760 14544
rect 8619 14504 8760 14532
rect 8619 14501 8631 14504
rect 8573 14495 8631 14501
rect 8754 14492 8760 14504
rect 8812 14492 8818 14544
rect 10796 14532 10824 14563
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 14182 14600 14188 14612
rect 14143 14572 14188 14600
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14884 14572 15117 14600
rect 14884 14560 14890 14572
rect 15105 14569 15117 14572
rect 15151 14600 15163 14603
rect 15378 14600 15384 14612
rect 15151 14572 15384 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 15378 14560 15384 14572
rect 15436 14560 15442 14612
rect 17218 14600 17224 14612
rect 17179 14572 17224 14600
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 19426 14600 19432 14612
rect 19387 14572 19432 14600
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 20530 14560 20536 14612
rect 20588 14600 20594 14612
rect 20625 14603 20683 14609
rect 20625 14600 20637 14603
rect 20588 14572 20637 14600
rect 20588 14560 20594 14572
rect 20625 14569 20637 14572
rect 20671 14600 20683 14603
rect 22557 14603 22615 14609
rect 22557 14600 22569 14603
rect 20671 14572 22569 14600
rect 20671 14569 20683 14572
rect 20625 14563 20683 14569
rect 22557 14569 22569 14572
rect 22603 14569 22615 14603
rect 24762 14600 24768 14612
rect 24723 14572 24768 14600
rect 22557 14563 22615 14569
rect 24762 14560 24768 14572
rect 24820 14560 24826 14612
rect 11977 14535 12035 14541
rect 10796 14504 11744 14532
rect 11716 14476 11744 14504
rect 11977 14501 11989 14535
rect 12023 14532 12035 14535
rect 12618 14532 12624 14544
rect 12023 14504 12624 14532
rect 12023 14501 12035 14504
rect 11977 14495 12035 14501
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 12986 14532 12992 14544
rect 12947 14504 12992 14532
rect 12986 14492 12992 14504
rect 13044 14492 13050 14544
rect 13541 14535 13599 14541
rect 13541 14501 13553 14535
rect 13587 14532 13599 14535
rect 14090 14532 14096 14544
rect 13587 14504 14096 14532
rect 13587 14501 13599 14504
rect 13541 14495 13599 14501
rect 14090 14492 14096 14504
rect 14148 14492 14154 14544
rect 14200 14532 14228 14560
rect 15473 14535 15531 14541
rect 15473 14532 15485 14535
rect 14200 14504 15485 14532
rect 15473 14501 15485 14504
rect 15519 14501 15531 14535
rect 17586 14532 17592 14544
rect 17547 14504 17592 14532
rect 15473 14495 15531 14501
rect 17586 14492 17592 14504
rect 17644 14492 17650 14544
rect 17681 14535 17739 14541
rect 17681 14501 17693 14535
rect 17727 14532 17739 14535
rect 18230 14532 18236 14544
rect 17727 14504 18236 14532
rect 17727 14501 17739 14504
rect 17681 14495 17739 14501
rect 18230 14492 18236 14504
rect 18288 14492 18294 14544
rect 21082 14532 21088 14544
rect 21043 14504 21088 14532
rect 21082 14492 21088 14504
rect 21140 14492 21146 14544
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 1578 14464 1584 14476
rect 1443 14436 1584 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 1578 14424 1584 14436
rect 1636 14424 1642 14476
rect 2682 14424 2688 14476
rect 2740 14464 2746 14476
rect 2996 14467 3054 14473
rect 2996 14464 3008 14467
rect 2740 14436 3008 14464
rect 2740 14424 2746 14436
rect 2996 14433 3008 14436
rect 3042 14433 3054 14467
rect 4062 14464 4068 14476
rect 4023 14436 4068 14464
rect 2996 14427 3054 14433
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 4522 14464 4528 14476
rect 4483 14436 4528 14464
rect 4522 14424 4528 14436
rect 4580 14424 4586 14476
rect 5166 14464 5172 14476
rect 5127 14436 5172 14464
rect 5166 14424 5172 14436
rect 5224 14424 5230 14476
rect 5534 14464 5540 14476
rect 5495 14436 5540 14464
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 6086 14464 6092 14476
rect 6047 14436 6092 14464
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 6270 14464 6276 14476
rect 6183 14436 6276 14464
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 9858 14464 9864 14476
rect 9819 14436 9864 14464
rect 9858 14424 9864 14436
rect 9916 14424 9922 14476
rect 10042 14424 10048 14476
rect 10100 14464 10106 14476
rect 10137 14467 10195 14473
rect 10137 14464 10149 14467
rect 10100 14436 10149 14464
rect 10100 14424 10106 14436
rect 10137 14433 10149 14436
rect 10183 14433 10195 14467
rect 11238 14464 11244 14476
rect 11199 14436 11244 14464
rect 10137 14427 10195 14433
rect 11238 14424 11244 14436
rect 11296 14424 11302 14476
rect 11698 14464 11704 14476
rect 11611 14436 11704 14464
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 20530 14424 20536 14476
rect 20588 14464 20594 14476
rect 20714 14464 20720 14476
rect 20588 14436 20720 14464
rect 20588 14424 20594 14436
rect 20714 14424 20720 14436
rect 20772 14424 20778 14476
rect 22462 14464 22468 14476
rect 22423 14436 22468 14464
rect 22462 14424 22468 14436
rect 22520 14424 22526 14476
rect 23014 14464 23020 14476
rect 22975 14436 23020 14464
rect 23014 14424 23020 14436
rect 23072 14424 23078 14476
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24854 14464 24860 14476
rect 24627 14436 24860 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 6362 14396 6368 14408
rect 6323 14368 6368 14396
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14396 7711 14399
rect 7926 14396 7932 14408
rect 7699 14368 7932 14396
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8294 14396 8300 14408
rect 8255 14368 8300 14396
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 9398 14356 9404 14408
rect 9456 14396 9462 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 9456 14368 10425 14396
rect 9456 14356 9462 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 12158 14356 12164 14408
rect 12216 14396 12222 14408
rect 12897 14399 12955 14405
rect 12897 14396 12909 14399
rect 12216 14368 12909 14396
rect 12216 14356 12222 14368
rect 12897 14365 12909 14368
rect 12943 14396 12955 14399
rect 13998 14396 14004 14408
rect 12943 14368 14004 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 13998 14356 14004 14368
rect 14056 14356 14062 14408
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 2314 14288 2320 14340
rect 2372 14328 2378 14340
rect 2372 14300 7788 14328
rect 2372 14288 2378 14300
rect 5166 14220 5172 14272
rect 5224 14260 5230 14272
rect 5534 14260 5540 14272
rect 5224 14232 5540 14260
rect 5224 14220 5230 14232
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 7193 14263 7251 14269
rect 7193 14229 7205 14263
rect 7239 14260 7251 14263
rect 7282 14260 7288 14272
rect 7239 14232 7288 14260
rect 7239 14229 7251 14232
rect 7193 14223 7251 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 7760 14260 7788 14300
rect 8202 14288 8208 14340
rect 8260 14328 8266 14340
rect 10962 14328 10968 14340
rect 8260 14300 10968 14328
rect 8260 14288 8266 14300
rect 10962 14288 10968 14300
rect 11020 14288 11026 14340
rect 15396 14328 15424 14359
rect 15562 14356 15568 14408
rect 15620 14396 15626 14408
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 15620 14368 15669 14396
rect 15620 14356 15626 14368
rect 15657 14365 15669 14368
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 19061 14399 19119 14405
rect 19061 14365 19073 14399
rect 19107 14396 19119 14399
rect 19150 14396 19156 14408
rect 19107 14368 19156 14396
rect 19107 14365 19119 14368
rect 19061 14359 19119 14365
rect 19150 14356 19156 14368
rect 19208 14356 19214 14408
rect 20990 14396 20996 14408
rect 20951 14368 20996 14396
rect 20990 14356 20996 14368
rect 21048 14356 21054 14408
rect 21450 14396 21456 14408
rect 21411 14368 21456 14396
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 15470 14328 15476 14340
rect 15383 14300 15476 14328
rect 15470 14288 15476 14300
rect 15528 14328 15534 14340
rect 17494 14328 17500 14340
rect 15528 14300 17500 14328
rect 15528 14288 15534 14300
rect 17494 14288 17500 14300
rect 17552 14288 17558 14340
rect 18141 14331 18199 14337
rect 18141 14297 18153 14331
rect 18187 14328 18199 14331
rect 19242 14328 19248 14340
rect 18187 14300 19248 14328
rect 18187 14297 18199 14300
rect 18141 14291 18199 14297
rect 19242 14288 19248 14300
rect 19300 14288 19306 14340
rect 20346 14328 20352 14340
rect 19438 14300 20352 14328
rect 8938 14260 8944 14272
rect 7760 14232 8944 14260
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 9490 14260 9496 14272
rect 9451 14232 9496 14260
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 16666 14220 16672 14272
rect 16724 14260 16730 14272
rect 19438 14260 19466 14300
rect 20346 14288 20352 14300
rect 20404 14288 20410 14340
rect 21542 14288 21548 14340
rect 21600 14328 21606 14340
rect 22281 14331 22339 14337
rect 22281 14328 22293 14331
rect 21600 14300 22293 14328
rect 21600 14288 21606 14300
rect 22281 14297 22293 14300
rect 22327 14328 22339 14331
rect 22922 14328 22928 14340
rect 22327 14300 22928 14328
rect 22327 14297 22339 14300
rect 22281 14291 22339 14297
rect 22922 14288 22928 14300
rect 22980 14288 22986 14340
rect 19978 14260 19984 14272
rect 16724 14232 19466 14260
rect 19939 14232 19984 14260
rect 16724 14220 16730 14232
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 21913 14263 21971 14269
rect 21913 14260 21925 14263
rect 21876 14232 21925 14260
rect 21876 14220 21882 14232
rect 21913 14229 21925 14232
rect 21959 14229 21971 14263
rect 23658 14260 23664 14272
rect 23619 14232 23664 14260
rect 21913 14223 21971 14229
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1762 14056 1768 14068
rect 1723 14028 1768 14056
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 4062 14056 4068 14068
rect 3476 14028 4068 14056
rect 3476 14016 3482 14028
rect 4062 14016 4068 14028
rect 4120 14056 4126 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 4120 14028 5641 14056
rect 4120 14016 4126 14028
rect 5629 14025 5641 14028
rect 5675 14025 5687 14059
rect 5629 14019 5687 14025
rect 6270 14016 6276 14068
rect 6328 14056 6334 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 6328 14028 6377 14056
rect 6328 14016 6334 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 8110 14056 8116 14068
rect 8071 14028 8116 14056
rect 6365 14019 6423 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 9858 14056 9864 14068
rect 9815 14028 9864 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 9950 14016 9956 14068
rect 10008 14056 10014 14068
rect 10008 14028 12480 14056
rect 10008 14016 10014 14028
rect 1780 13988 1808 14016
rect 5534 13988 5540 14000
rect 1780 13960 5540 13988
rect 1780 13852 1808 13960
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 6546 13948 6552 14000
rect 6604 13988 6610 14000
rect 6822 13988 6828 14000
rect 6604 13960 6828 13988
rect 6604 13948 6610 13960
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 7161 13960 7788 13988
rect 2682 13920 2688 13932
rect 2643 13892 2688 13920
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 5350 13920 5356 13932
rect 4203 13892 5212 13920
rect 5311 13892 5356 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 1857 13855 1915 13861
rect 1857 13852 1869 13855
rect 1780 13824 1869 13852
rect 1857 13821 1869 13824
rect 1903 13821 1915 13855
rect 2866 13852 2872 13864
rect 2827 13824 2872 13852
rect 1857 13815 1915 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 4890 13852 4896 13864
rect 4571 13824 4896 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5184 13861 5212 13892
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 7161 13920 7189 13960
rect 7466 13920 7472 13932
rect 5500 13892 7189 13920
rect 7427 13892 7472 13920
rect 5500 13880 5506 13892
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 7760 13920 7788 13960
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 8803 13991 8861 13997
rect 8803 13988 8815 13991
rect 7892 13960 8815 13988
rect 7892 13948 7898 13960
rect 8803 13957 8815 13960
rect 8849 13957 8861 13991
rect 8803 13951 8861 13957
rect 9030 13948 9036 14000
rect 9088 13988 9094 14000
rect 10134 13988 10140 14000
rect 9088 13960 10140 13988
rect 9088 13948 9094 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 11698 13988 11704 14000
rect 11659 13960 11704 13988
rect 11698 13948 11704 13960
rect 11756 13948 11762 14000
rect 10152 13920 10180 13948
rect 12452 13932 12480 14028
rect 12986 14016 12992 14068
rect 13044 14056 13050 14068
rect 13357 14059 13415 14065
rect 13357 14056 13369 14059
rect 13044 14028 13369 14056
rect 13044 14016 13050 14028
rect 13357 14025 13369 14028
rect 13403 14056 13415 14059
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 13403 14028 13645 14056
rect 13403 14025 13415 14028
rect 13357 14019 13415 14025
rect 13633 14025 13645 14028
rect 13679 14056 13691 14059
rect 13998 14056 14004 14068
rect 13679 14028 13814 14056
rect 13959 14028 14004 14056
rect 13679 14025 13691 14028
rect 13633 14019 13691 14025
rect 13786 13988 13814 14028
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 14829 14059 14887 14065
rect 14829 14056 14841 14059
rect 14240 14028 14841 14056
rect 14240 14016 14246 14028
rect 14829 14025 14841 14028
rect 14875 14056 14887 14059
rect 14921 14059 14979 14065
rect 14921 14056 14933 14059
rect 14875 14028 14933 14056
rect 14875 14025 14887 14028
rect 14829 14019 14887 14025
rect 14921 14025 14933 14028
rect 14967 14025 14979 14059
rect 14921 14019 14979 14025
rect 16853 14059 16911 14065
rect 16853 14025 16865 14059
rect 16899 14056 16911 14059
rect 18230 14056 18236 14068
rect 16899 14028 18236 14056
rect 16899 14025 16911 14028
rect 16853 14019 16911 14025
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 19978 14016 19984 14068
rect 20036 14056 20042 14068
rect 20901 14059 20959 14065
rect 20901 14056 20913 14059
rect 20036 14028 20913 14056
rect 20036 14016 20042 14028
rect 20901 14025 20913 14028
rect 20947 14056 20959 14059
rect 21082 14056 21088 14068
rect 20947 14028 21088 14056
rect 20947 14025 20959 14028
rect 20901 14019 20959 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 22462 14056 22468 14068
rect 22423 14028 22468 14056
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 24765 14059 24823 14065
rect 24765 14025 24777 14059
rect 24811 14056 24823 14059
rect 24854 14056 24860 14068
rect 24811 14028 24860 14056
rect 24811 14025 24823 14028
rect 24765 14019 24823 14025
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 15378 13988 15384 14000
rect 13786 13960 15384 13988
rect 15378 13948 15384 13960
rect 15436 13948 15442 14000
rect 15749 13991 15807 13997
rect 15749 13957 15761 13991
rect 15795 13988 15807 13991
rect 15838 13988 15844 14000
rect 15795 13960 15844 13988
rect 15795 13957 15807 13960
rect 15749 13951 15807 13957
rect 15838 13948 15844 13960
rect 15896 13988 15902 14000
rect 17218 13988 17224 14000
rect 15896 13960 17224 13988
rect 15896 13948 15902 13960
rect 17218 13948 17224 13960
rect 17276 13948 17282 14000
rect 19242 13948 19248 14000
rect 19300 13988 19306 14000
rect 19300 13960 20208 13988
rect 19300 13948 19306 13960
rect 11882 13920 11888 13932
rect 7760 13892 7880 13920
rect 10152 13892 11888 13920
rect 5169 13855 5227 13861
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5258 13852 5264 13864
rect 5215 13824 5264 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 7852 13852 7880 13892
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 12434 13920 12440 13932
rect 12347 13892 12440 13920
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15194 13920 15200 13932
rect 14875 13892 15200 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15194 13880 15200 13892
rect 15252 13920 15258 13932
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 15252 13892 16129 13920
rect 15252 13880 15258 13892
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20070 13920 20076 13932
rect 19935 13892 20076 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20180 13929 20208 13960
rect 20165 13923 20223 13929
rect 20165 13889 20177 13923
rect 20211 13920 20223 13923
rect 21453 13923 21511 13929
rect 21453 13920 21465 13923
rect 20211 13892 21465 13920
rect 20211 13889 20223 13892
rect 20165 13883 20223 13889
rect 21453 13889 21465 13892
rect 21499 13920 21511 13923
rect 21542 13920 21548 13932
rect 21499 13892 21548 13920
rect 21499 13889 21511 13892
rect 21453 13883 21511 13889
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 21634 13880 21640 13932
rect 21692 13920 21698 13932
rect 21729 13923 21787 13929
rect 21729 13920 21741 13923
rect 21692 13892 21741 13920
rect 21692 13880 21698 13892
rect 21729 13889 21741 13892
rect 21775 13889 21787 13923
rect 21729 13883 21787 13889
rect 22370 13880 22376 13932
rect 22428 13920 22434 13932
rect 24762 13920 24768 13932
rect 22428 13892 24768 13920
rect 22428 13880 22434 13892
rect 24762 13880 24768 13892
rect 24820 13880 24826 13932
rect 8700 13855 8758 13861
rect 8700 13852 8712 13855
rect 7852 13824 8712 13852
rect 8700 13821 8712 13824
rect 8746 13852 8758 13855
rect 9214 13852 9220 13864
rect 8746 13824 9220 13852
rect 8746 13821 8758 13824
rect 8700 13815 8758 13821
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 11698 13852 11704 13864
rect 11480 13824 11704 13852
rect 11480 13812 11486 13824
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 16298 13812 16304 13864
rect 16356 13852 16362 13864
rect 16980 13855 17038 13861
rect 16980 13852 16992 13855
rect 16356 13824 16992 13852
rect 16356 13812 16362 13824
rect 16980 13821 16992 13824
rect 17026 13852 17038 13855
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 17026 13824 17417 13852
rect 17026 13821 17038 13824
rect 16980 13815 17038 13821
rect 17405 13821 17417 13824
rect 17451 13821 17463 13855
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 18971 13824 19073 13852
rect 17405 13815 17463 13821
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 2409 13787 2467 13793
rect 2409 13753 2421 13787
rect 2455 13784 2467 13787
rect 3231 13787 3289 13793
rect 3231 13784 3243 13787
rect 2455 13756 3243 13784
rect 2455 13753 2467 13756
rect 2409 13747 2467 13753
rect 3231 13753 3243 13756
rect 3277 13784 3289 13787
rect 4338 13784 4344 13796
rect 3277 13756 4344 13784
rect 3277 13753 3289 13756
rect 3231 13747 3289 13753
rect 4338 13744 4344 13756
rect 4396 13744 4402 13796
rect 6086 13784 6092 13796
rect 6047 13756 6092 13784
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 7193 13787 7251 13793
rect 7193 13753 7205 13787
rect 7239 13753 7251 13787
rect 7193 13747 7251 13753
rect 2038 13716 2044 13728
rect 1999 13688 2044 13716
rect 2038 13676 2044 13688
rect 2096 13676 2102 13728
rect 3786 13716 3792 13728
rect 3747 13688 3792 13716
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 7208 13716 7236 13747
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 7340 13756 7385 13784
rect 7340 13744 7346 13756
rect 9858 13744 9864 13796
rect 9916 13784 9922 13796
rect 10045 13787 10103 13793
rect 10045 13784 10057 13787
rect 9916 13756 10057 13784
rect 9916 13744 9922 13756
rect 10045 13753 10057 13756
rect 10091 13753 10103 13787
rect 10045 13747 10103 13753
rect 10134 13744 10140 13796
rect 10192 13784 10198 13796
rect 10686 13784 10692 13796
rect 10192 13756 10237 13784
rect 10647 13756 10692 13784
rect 10192 13744 10198 13756
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 11238 13784 11244 13796
rect 11199 13756 11244 13784
rect 11238 13744 11244 13756
rect 11296 13744 11302 13796
rect 12758 13787 12816 13793
rect 12758 13753 12770 13787
rect 12804 13753 12816 13787
rect 12758 13747 12816 13753
rect 14645 13787 14703 13793
rect 14645 13753 14657 13787
rect 14691 13784 14703 13787
rect 15194 13784 15200 13796
rect 14691 13756 15200 13784
rect 14691 13753 14703 13756
rect 14645 13747 14703 13753
rect 7742 13716 7748 13728
rect 7208 13688 7748 13716
rect 7742 13676 7748 13688
rect 7800 13676 7806 13728
rect 9214 13716 9220 13728
rect 9175 13688 9220 13716
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 9490 13676 9496 13728
rect 9548 13716 9554 13728
rect 9950 13716 9956 13728
rect 9548 13688 9956 13716
rect 9548 13676 9554 13688
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 12158 13716 12164 13728
rect 12119 13688 12164 13716
rect 12158 13676 12164 13688
rect 12216 13716 12222 13728
rect 12773 13716 12801 13747
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 17083 13787 17141 13793
rect 15344 13756 15389 13784
rect 15344 13744 15350 13756
rect 17083 13753 17095 13787
rect 17129 13784 17141 13787
rect 18138 13784 18144 13796
rect 17129 13756 18144 13784
rect 17129 13753 17141 13756
rect 17083 13747 17141 13753
rect 18138 13744 18144 13756
rect 18196 13744 18202 13796
rect 18230 13744 18236 13796
rect 18288 13784 18294 13796
rect 18785 13787 18843 13793
rect 18288 13756 18333 13784
rect 18288 13744 18294 13756
rect 18785 13753 18797 13787
rect 18831 13784 18843 13787
rect 18966 13784 18972 13796
rect 18831 13756 18972 13784
rect 18831 13753 18843 13756
rect 18785 13747 18843 13753
rect 18966 13744 18972 13756
rect 19024 13744 19030 13796
rect 19076 13784 19104 13815
rect 22738 13812 22744 13864
rect 22796 13852 22802 13864
rect 23658 13852 23664 13864
rect 22796 13824 23664 13852
rect 22796 13812 22802 13824
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 24075 13855 24133 13861
rect 24075 13852 24087 13855
rect 23768 13824 24087 13852
rect 19518 13784 19524 13796
rect 19076 13756 19524 13784
rect 19518 13744 19524 13756
rect 19576 13744 19582 13796
rect 19705 13787 19763 13793
rect 19705 13753 19717 13787
rect 19751 13784 19763 13787
rect 19978 13784 19984 13796
rect 19751 13756 19984 13784
rect 19751 13753 19763 13756
rect 19705 13747 19763 13753
rect 19978 13744 19984 13756
rect 20036 13744 20042 13796
rect 21545 13787 21603 13793
rect 21545 13753 21557 13787
rect 21591 13784 21603 13787
rect 21818 13784 21824 13796
rect 21591 13756 21824 13784
rect 21591 13753 21603 13756
rect 21545 13747 21603 13753
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 23768 13784 23796 13824
rect 24075 13821 24087 13824
rect 24121 13821 24133 13855
rect 24075 13815 24133 13821
rect 24670 13812 24676 13864
rect 24728 13852 24734 13864
rect 24854 13852 24860 13864
rect 24728 13824 24860 13852
rect 24728 13812 24734 13824
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 25292 13855 25350 13861
rect 25292 13821 25304 13855
rect 25338 13852 25350 13855
rect 25682 13852 25688 13864
rect 25338 13824 25688 13852
rect 25338 13821 25350 13824
rect 25292 13815 25350 13821
rect 25682 13812 25688 13824
rect 25740 13812 25746 13864
rect 23492 13756 23796 13784
rect 12986 13716 12992 13728
rect 12216 13688 12992 13716
rect 12216 13676 12222 13688
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 17865 13719 17923 13725
rect 17865 13685 17877 13719
rect 17911 13716 17923 13719
rect 18248 13716 18276 13744
rect 23492 13728 23520 13756
rect 17911 13688 18276 13716
rect 17911 13685 17923 13688
rect 17865 13679 17923 13685
rect 19058 13676 19064 13728
rect 19116 13716 19122 13728
rect 20346 13716 20352 13728
rect 19116 13688 20352 13716
rect 19116 13676 19122 13688
rect 20346 13676 20352 13688
rect 20404 13676 20410 13728
rect 22925 13719 22983 13725
rect 22925 13685 22937 13719
rect 22971 13716 22983 13719
rect 23014 13716 23020 13728
rect 22971 13688 23020 13716
rect 22971 13685 22983 13688
rect 22925 13679 22983 13685
rect 23014 13676 23020 13688
rect 23072 13716 23078 13728
rect 23474 13716 23480 13728
rect 23072 13688 23480 13716
rect 23072 13676 23078 13688
rect 23474 13676 23480 13688
rect 23532 13676 23538 13728
rect 23750 13716 23756 13728
rect 23711 13688 23756 13716
rect 23750 13676 23756 13688
rect 23808 13676 23814 13728
rect 24118 13676 24124 13728
rect 24176 13716 24182 13728
rect 25363 13719 25421 13725
rect 25363 13716 25375 13719
rect 24176 13688 25375 13716
rect 24176 13676 24182 13688
rect 25363 13685 25375 13688
rect 25409 13685 25421 13719
rect 25363 13679 25421 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2038 13472 2044 13524
rect 2096 13512 2102 13524
rect 3881 13515 3939 13521
rect 3881 13512 3893 13515
rect 2096 13484 3893 13512
rect 2096 13472 2102 13484
rect 3881 13481 3893 13484
rect 3927 13481 3939 13515
rect 3881 13475 3939 13481
rect 2409 13447 2467 13453
rect 2409 13413 2421 13447
rect 2455 13444 2467 13447
rect 2682 13444 2688 13456
rect 2455 13416 2688 13444
rect 2455 13413 2467 13416
rect 2409 13407 2467 13413
rect 2682 13404 2688 13416
rect 2740 13444 2746 13456
rect 3786 13444 3792 13456
rect 2740 13416 3792 13444
rect 2740 13404 2746 13416
rect 3786 13404 3792 13416
rect 3844 13404 3850 13456
rect 3896 13376 3924 13475
rect 3970 13472 3976 13524
rect 4028 13512 4034 13524
rect 4154 13512 4160 13524
rect 4028 13484 4160 13512
rect 4028 13472 4034 13484
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4433 13515 4491 13521
rect 4433 13512 4445 13515
rect 4396 13484 4445 13512
rect 4396 13472 4402 13484
rect 4433 13481 4445 13484
rect 4479 13512 4491 13515
rect 4798 13512 4804 13524
rect 4479 13484 4804 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 6181 13515 6239 13521
rect 6181 13481 6193 13515
rect 6227 13512 6239 13515
rect 6362 13512 6368 13524
rect 6227 13484 6368 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 4522 13376 4528 13388
rect 3160 13348 3832 13376
rect 3896 13348 4528 13376
rect 1670 13268 1676 13320
rect 1728 13308 1734 13320
rect 2317 13311 2375 13317
rect 2317 13308 2329 13311
rect 1728 13280 2329 13308
rect 1728 13268 1734 13280
rect 2317 13277 2329 13280
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 2498 13268 2504 13320
rect 2556 13308 2562 13320
rect 2593 13311 2651 13317
rect 2593 13308 2605 13311
rect 2556 13280 2605 13308
rect 2556 13268 2562 13280
rect 2593 13277 2605 13280
rect 2639 13308 2651 13311
rect 3160 13308 3188 13348
rect 3804 13320 3832 13348
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 6288 13385 6316 13484
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 6546 13472 6552 13524
rect 6604 13512 6610 13524
rect 6641 13515 6699 13521
rect 6641 13512 6653 13515
rect 6604 13484 6653 13512
rect 6604 13472 6610 13484
rect 6641 13481 6653 13484
rect 6687 13481 6699 13515
rect 6641 13475 6699 13481
rect 7193 13515 7251 13521
rect 7193 13481 7205 13515
rect 7239 13512 7251 13515
rect 7282 13512 7288 13524
rect 7239 13484 7288 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 9858 13512 9864 13524
rect 7524 13484 8800 13512
rect 7524 13472 7530 13484
rect 8202 13444 8208 13456
rect 8163 13416 8208 13444
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 8772 13453 8800 13484
rect 9048 13484 9864 13512
rect 8757 13447 8815 13453
rect 8757 13413 8769 13447
rect 8803 13413 8815 13447
rect 8757 13407 8815 13413
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13345 6331 13379
rect 6273 13339 6331 13345
rect 2639 13280 3188 13308
rect 2639 13277 2651 13280
rect 2593 13271 2651 13277
rect 3234 13268 3240 13320
rect 3292 13268 3298 13320
rect 3786 13268 3792 13320
rect 3844 13268 3850 13320
rect 4062 13308 4068 13320
rect 4023 13280 4068 13308
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 9048 13317 9076 13484
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 11606 13512 11612 13524
rect 11567 13484 11612 13512
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 12434 13512 12440 13524
rect 12395 13484 12440 13512
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 12986 13512 12992 13524
rect 12947 13484 12992 13512
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 14182 13512 14188 13524
rect 13587 13484 14188 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 17865 13515 17923 13521
rect 17865 13512 17877 13515
rect 17644 13484 17877 13512
rect 17644 13472 17650 13484
rect 17865 13481 17877 13484
rect 17911 13481 17923 13515
rect 17865 13475 17923 13481
rect 18138 13472 18144 13524
rect 18196 13512 18202 13524
rect 18233 13515 18291 13521
rect 18233 13512 18245 13515
rect 18196 13484 18245 13512
rect 18196 13472 18202 13484
rect 18233 13481 18245 13484
rect 18279 13481 18291 13515
rect 18233 13475 18291 13481
rect 19058 13472 19064 13524
rect 19116 13512 19122 13524
rect 19889 13515 19947 13521
rect 19116 13484 19564 13512
rect 19116 13472 19122 13484
rect 9582 13404 9588 13456
rect 9640 13444 9646 13456
rect 9998 13447 10056 13453
rect 9998 13444 10010 13447
rect 9640 13416 10010 13444
rect 9640 13404 9646 13416
rect 9998 13413 10010 13416
rect 10044 13413 10056 13447
rect 9998 13407 10056 13413
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 15473 13447 15531 13453
rect 15473 13444 15485 13447
rect 15436 13416 15485 13444
rect 15436 13404 15442 13416
rect 15473 13413 15485 13416
rect 15519 13413 15531 13447
rect 17034 13444 17040 13456
rect 16995 13416 17040 13444
rect 15473 13407 15531 13413
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 18601 13447 18659 13453
rect 18601 13444 18613 13447
rect 18564 13416 18613 13444
rect 18564 13404 18570 13416
rect 18601 13413 18613 13416
rect 18647 13413 18659 13447
rect 18601 13407 18659 13413
rect 19153 13447 19211 13453
rect 19153 13413 19165 13447
rect 19199 13444 19211 13447
rect 19242 13444 19248 13456
rect 19199 13416 19248 13444
rect 19199 13413 19211 13416
rect 19153 13407 19211 13413
rect 19242 13404 19248 13416
rect 19300 13404 19306 13456
rect 19536 13453 19564 13484
rect 19889 13481 19901 13515
rect 19935 13512 19947 13515
rect 20070 13512 20076 13524
rect 19935 13484 20076 13512
rect 19935 13481 19947 13484
rect 19889 13475 19947 13481
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 20717 13515 20775 13521
rect 20717 13481 20729 13515
rect 20763 13512 20775 13515
rect 20990 13512 20996 13524
rect 20763 13484 20996 13512
rect 20763 13481 20775 13484
rect 20717 13475 20775 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 23750 13512 23756 13524
rect 21094 13484 23756 13512
rect 19521 13447 19579 13453
rect 19521 13413 19533 13447
rect 19567 13444 19579 13447
rect 21094 13444 21122 13484
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 21542 13444 21548 13456
rect 19567 13416 21122 13444
rect 21503 13416 21548 13444
rect 19567 13413 19579 13416
rect 19521 13407 19579 13413
rect 21542 13404 21548 13416
rect 21600 13404 21606 13456
rect 22830 13404 22836 13456
rect 22888 13444 22894 13456
rect 23109 13447 23167 13453
rect 23109 13444 23121 13447
rect 22888 13416 23121 13444
rect 22888 13404 22894 13416
rect 23109 13413 23121 13416
rect 23155 13413 23167 13447
rect 23109 13407 23167 13413
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 9858 13376 9864 13388
rect 9456 13348 9864 13376
rect 9456 13336 9462 13348
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13345 10655 13379
rect 10597 13339 10655 13345
rect 11425 13379 11483 13385
rect 11425 13345 11437 13379
rect 11471 13376 11483 13379
rect 12066 13376 12072 13388
rect 11471 13348 12072 13376
rect 11471 13345 11483 13348
rect 11425 13339 11483 13345
rect 9033 13311 9091 13317
rect 9033 13308 9045 13311
rect 8220 13280 9045 13308
rect 3252 13240 3280 13268
rect 8220 13240 8248 13280
rect 9033 13277 9045 13280
rect 9079 13277 9091 13311
rect 9674 13308 9680 13320
rect 9635 13280 9680 13308
rect 9033 13271 9091 13277
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 9950 13268 9956 13320
rect 10008 13308 10014 13320
rect 10134 13308 10140 13320
rect 10008 13280 10140 13308
rect 10008 13268 10014 13280
rect 10134 13268 10140 13280
rect 10192 13308 10198 13320
rect 10612 13308 10640 13339
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 24540 13379 24598 13385
rect 24540 13345 24552 13379
rect 24586 13376 24598 13379
rect 24762 13376 24768 13388
rect 24586 13348 24768 13376
rect 24586 13345 24598 13348
rect 24540 13339 24598 13345
rect 24762 13336 24768 13348
rect 24820 13336 24826 13388
rect 10192 13280 10640 13308
rect 10192 13268 10198 13280
rect 12434 13268 12440 13320
rect 12492 13308 12498 13320
rect 12621 13311 12679 13317
rect 12621 13308 12633 13311
rect 12492 13280 12633 13308
rect 12492 13268 12498 13280
rect 12621 13277 12633 13280
rect 12667 13277 12679 13311
rect 12621 13271 12679 13277
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 14608 13280 15393 13308
rect 14608 13268 14614 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 16942 13308 16948 13320
rect 16903 13280 16948 13308
rect 15381 13271 15439 13277
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 17218 13308 17224 13320
rect 17179 13280 17224 13308
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 18506 13308 18512 13320
rect 18467 13280 18512 13308
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18966 13268 18972 13320
rect 19024 13308 19030 13320
rect 21450 13308 21456 13320
rect 19024 13280 21456 13308
rect 19024 13268 19030 13280
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 21634 13268 21640 13320
rect 21692 13308 21698 13320
rect 21729 13311 21787 13317
rect 21729 13308 21741 13311
rect 21692 13280 21741 13308
rect 21692 13268 21698 13280
rect 21729 13277 21741 13280
rect 21775 13277 21787 13311
rect 23014 13308 23020 13320
rect 22975 13280 23020 13308
rect 21729 13271 21787 13277
rect 23014 13268 23020 13280
rect 23072 13308 23078 13320
rect 24627 13311 24685 13317
rect 24627 13308 24639 13311
rect 23072 13280 24639 13308
rect 23072 13268 23078 13280
rect 24627 13277 24639 13280
rect 24673 13277 24685 13311
rect 24627 13271 24685 13277
rect 3252 13212 8248 13240
rect 8570 13200 8576 13252
rect 8628 13240 8634 13252
rect 9493 13243 9551 13249
rect 9493 13240 9505 13243
rect 8628 13212 9505 13240
rect 8628 13200 8634 13212
rect 9493 13209 9505 13212
rect 9539 13240 9551 13243
rect 10042 13240 10048 13252
rect 9539 13212 10048 13240
rect 9539 13209 9551 13212
rect 9493 13203 9551 13209
rect 10042 13200 10048 13212
rect 10100 13200 10106 13252
rect 15105 13243 15163 13249
rect 15105 13209 15117 13243
rect 15151 13240 15163 13243
rect 15470 13240 15476 13252
rect 15151 13212 15476 13240
rect 15151 13209 15163 13212
rect 15105 13203 15163 13209
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 15933 13243 15991 13249
rect 15933 13240 15945 13243
rect 15620 13212 15945 13240
rect 15620 13200 15626 13212
rect 15933 13209 15945 13212
rect 15979 13240 15991 13243
rect 16022 13240 16028 13252
rect 15979 13212 16028 13240
rect 15979 13209 15991 13212
rect 15933 13203 15991 13209
rect 16022 13200 16028 13212
rect 16080 13200 16086 13252
rect 21468 13240 21496 13268
rect 22094 13240 22100 13252
rect 21468 13212 22100 13240
rect 22094 13200 22100 13212
rect 22152 13240 22158 13252
rect 23569 13243 23627 13249
rect 23569 13240 23581 13243
rect 22152 13212 23581 13240
rect 22152 13200 22158 13212
rect 23569 13209 23581 13212
rect 23615 13209 23627 13243
rect 23569 13203 23627 13209
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 3237 13175 3295 13181
rect 3237 13172 3249 13175
rect 2832 13144 3249 13172
rect 2832 13132 2838 13144
rect 3237 13141 3249 13144
rect 3283 13172 3295 13175
rect 3970 13172 3976 13184
rect 3283 13144 3976 13172
rect 3283 13141 3295 13144
rect 3237 13135 3295 13141
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 4338 13132 4344 13184
rect 4396 13172 4402 13184
rect 4985 13175 5043 13181
rect 4985 13172 4997 13175
rect 4396 13144 4997 13172
rect 4396 13132 4402 13144
rect 4985 13141 4997 13144
rect 5031 13141 5043 13175
rect 4985 13135 5043 13141
rect 7561 13175 7619 13181
rect 7561 13141 7573 13175
rect 7607 13172 7619 13175
rect 7742 13172 7748 13184
rect 7607 13144 7748 13172
rect 7607 13141 7619 13144
rect 7561 13135 7619 13141
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 7926 13172 7932 13184
rect 7839 13144 7932 13172
rect 7926 13132 7932 13144
rect 7984 13172 7990 13184
rect 8294 13172 8300 13184
rect 7984 13144 8300 13172
rect 7984 13132 7990 13144
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 12802 13172 12808 13184
rect 8812 13144 12808 13172
rect 8812 13132 8818 13144
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 13817 13175 13875 13181
rect 13817 13172 13829 13175
rect 13688 13144 13829 13172
rect 13688 13132 13694 13144
rect 13817 13141 13829 13144
rect 13863 13141 13875 13175
rect 13817 13135 13875 13141
rect 20990 13132 20996 13184
rect 21048 13172 21054 13184
rect 21085 13175 21143 13181
rect 21085 13172 21097 13175
rect 21048 13144 21097 13172
rect 21048 13132 21054 13144
rect 21085 13141 21097 13144
rect 21131 13141 21143 13175
rect 21085 13135 21143 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1670 12968 1676 12980
rect 1631 12940 1676 12968
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12968 2007 12971
rect 2314 12968 2320 12980
rect 1995 12940 2320 12968
rect 1995 12937 2007 12940
rect 1949 12931 2007 12937
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 2682 12968 2688 12980
rect 2643 12940 2688 12968
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 3694 12968 3700 12980
rect 3655 12940 3700 12968
rect 3694 12928 3700 12940
rect 3752 12928 3758 12980
rect 4798 12968 4804 12980
rect 4759 12940 4804 12968
rect 4798 12928 4804 12940
rect 4856 12968 4862 12980
rect 5445 12971 5503 12977
rect 5445 12968 5457 12971
rect 4856 12940 5457 12968
rect 4856 12928 4862 12940
rect 5445 12937 5457 12940
rect 5491 12937 5503 12971
rect 5445 12931 5503 12937
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 7745 12971 7803 12977
rect 6144 12940 7696 12968
rect 6144 12928 6150 12940
rect 2961 12903 3019 12909
rect 2961 12869 2973 12903
rect 3007 12900 3019 12903
rect 3007 12872 3648 12900
rect 3007 12869 3019 12872
rect 2961 12863 3019 12869
rect 2406 12792 2412 12844
rect 2464 12832 2470 12844
rect 3050 12832 3056 12844
rect 2464 12804 3056 12832
rect 2464 12792 2470 12804
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12764 1823 12767
rect 2317 12767 2375 12773
rect 2317 12764 2329 12767
rect 1811 12736 2329 12764
rect 1811 12733 1823 12736
rect 1765 12727 1823 12733
rect 2317 12733 2329 12736
rect 2363 12764 2375 12767
rect 2777 12767 2835 12773
rect 2777 12764 2789 12767
rect 2363 12736 2789 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 2777 12733 2789 12736
rect 2823 12764 2835 12767
rect 3620 12764 3648 12872
rect 3712 12832 3740 12928
rect 3786 12860 3792 12912
rect 3844 12900 3850 12912
rect 4433 12903 4491 12909
rect 4433 12900 4445 12903
rect 3844 12872 4445 12900
rect 3844 12860 3850 12872
rect 4433 12869 4445 12872
rect 4479 12900 4491 12903
rect 7466 12900 7472 12912
rect 4479 12872 7472 12900
rect 4479 12869 4491 12872
rect 4433 12863 4491 12869
rect 7466 12860 7472 12872
rect 7524 12860 7530 12912
rect 7668 12900 7696 12940
rect 7745 12937 7757 12971
rect 7791 12968 7803 12971
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 7791 12940 8125 12968
rect 7791 12937 7803 12940
rect 7745 12931 7803 12937
rect 8113 12937 8125 12940
rect 8159 12968 8171 12971
rect 8202 12968 8208 12980
rect 8159 12940 8208 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 11471 12971 11529 12977
rect 11471 12968 11483 12971
rect 8352 12940 11483 12968
rect 8352 12928 8358 12940
rect 11471 12937 11483 12940
rect 11517 12937 11529 12971
rect 11471 12931 11529 12937
rect 12986 12928 12992 12980
rect 13044 12968 13050 12980
rect 13265 12971 13323 12977
rect 13265 12968 13277 12971
rect 13044 12940 13277 12968
rect 13044 12928 13050 12940
rect 13265 12937 13277 12940
rect 13311 12968 13323 12971
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 13311 12940 13369 12968
rect 13311 12937 13323 12940
rect 13265 12931 13323 12937
rect 13357 12937 13369 12940
rect 13403 12937 13415 12971
rect 13357 12931 13415 12937
rect 13722 12928 13728 12980
rect 13780 12968 13786 12980
rect 14921 12971 14979 12977
rect 14921 12968 14933 12971
rect 13780 12940 14933 12968
rect 13780 12928 13786 12940
rect 14921 12937 14933 12940
rect 14967 12968 14979 12971
rect 15197 12971 15255 12977
rect 15197 12968 15209 12971
rect 14967 12940 15209 12968
rect 14967 12937 14979 12940
rect 14921 12931 14979 12937
rect 15197 12937 15209 12940
rect 15243 12937 15255 12971
rect 15378 12968 15384 12980
rect 15339 12940 15384 12968
rect 15197 12931 15255 12937
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 21542 12928 21548 12980
rect 21600 12968 21606 12980
rect 22005 12971 22063 12977
rect 22005 12968 22017 12971
rect 21600 12940 22017 12968
rect 21600 12928 21606 12940
rect 22005 12937 22017 12940
rect 22051 12937 22063 12971
rect 22005 12931 22063 12937
rect 22465 12971 22523 12977
rect 22465 12937 22477 12971
rect 22511 12968 22523 12971
rect 23014 12968 23020 12980
rect 22511 12940 23020 12968
rect 22511 12937 22523 12940
rect 22465 12931 22523 12937
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 24946 12968 24952 12980
rect 24907 12940 24952 12968
rect 24946 12928 24952 12940
rect 25004 12928 25010 12980
rect 8754 12900 8760 12912
rect 7668 12872 8760 12900
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 10962 12860 10968 12912
rect 11020 12900 11026 12912
rect 12667 12903 12725 12909
rect 11020 12872 11443 12900
rect 11020 12860 11026 12872
rect 3881 12835 3939 12841
rect 3881 12832 3893 12835
rect 3712 12804 3893 12832
rect 3881 12801 3893 12804
rect 3927 12801 3939 12835
rect 3881 12795 3939 12801
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 4120 12804 5181 12832
rect 4120 12792 4126 12804
rect 5169 12801 5181 12804
rect 5215 12801 5227 12835
rect 5169 12795 5227 12801
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 6273 12835 6331 12841
rect 6273 12832 6285 12835
rect 5491 12804 6285 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 6273 12801 6285 12804
rect 6319 12832 6331 12835
rect 6546 12832 6552 12844
rect 6319 12804 6552 12832
rect 6319 12801 6331 12804
rect 6273 12795 6331 12801
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9180 12804 9873 12832
rect 9180 12792 9186 12804
rect 9861 12801 9873 12804
rect 9907 12832 9919 12835
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 9907 12804 11161 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 11149 12801 11161 12804
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 3694 12764 3700 12776
rect 2823 12736 3372 12764
rect 3620 12736 3700 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 3344 12640 3372 12736
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 5721 12727 5779 12733
rect 3973 12699 4031 12705
rect 3973 12665 3985 12699
rect 4019 12696 4031 12699
rect 4338 12696 4344 12708
rect 4019 12668 4344 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 5629 12699 5687 12705
rect 5629 12665 5641 12699
rect 5675 12696 5687 12699
rect 5736 12696 5764 12727
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 11415 12773 11443 12872
rect 12667 12869 12679 12903
rect 12713 12900 12725 12903
rect 14826 12900 14832 12912
rect 12713 12872 14832 12900
rect 12713 12869 12725 12872
rect 12667 12863 12725 12869
rect 14826 12860 14832 12872
rect 14884 12860 14890 12912
rect 16390 12900 16396 12912
rect 15856 12872 16396 12900
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 13630 12832 13636 12844
rect 13044 12804 13636 12832
rect 13044 12792 13050 12804
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 15856 12841 15884 12872
rect 16390 12860 16396 12872
rect 16448 12900 16454 12912
rect 25179 12903 25237 12909
rect 25179 12900 25191 12903
rect 16448 12872 25191 12900
rect 16448 12860 16454 12872
rect 25179 12869 25191 12872
rect 25225 12869 25237 12903
rect 25590 12900 25596 12912
rect 25551 12872 25596 12900
rect 25179 12863 25237 12869
rect 25590 12860 25596 12872
rect 25648 12860 25654 12912
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 16022 12792 16028 12844
rect 16080 12832 16086 12844
rect 16117 12835 16175 12841
rect 16117 12832 16129 12835
rect 16080 12804 16129 12832
rect 16080 12792 16086 12804
rect 16117 12801 16129 12804
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 17368 12804 18337 12832
rect 17368 12792 17374 12804
rect 18325 12801 18337 12804
rect 18371 12832 18383 12835
rect 18782 12832 18788 12844
rect 18371 12804 18788 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 18966 12832 18972 12844
rect 18927 12804 18972 12832
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 20349 12835 20407 12841
rect 20349 12832 20361 12835
rect 19879 12804 20361 12832
rect 19879 12773 19907 12804
rect 20349 12801 20361 12804
rect 20395 12832 20407 12835
rect 21174 12832 21180 12844
rect 20395 12804 21180 12832
rect 20395 12801 20407 12804
rect 20349 12795 20407 12801
rect 21174 12792 21180 12804
rect 21232 12792 21238 12844
rect 23109 12835 23167 12841
rect 23109 12832 23121 12835
rect 22639 12804 23121 12832
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 6972 12736 8585 12764
rect 6972 12724 6978 12736
rect 8573 12733 8585 12736
rect 8619 12764 8631 12767
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8619 12736 9045 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 11400 12767 11458 12773
rect 11400 12733 11412 12767
rect 11446 12764 11458 12767
rect 12596 12767 12654 12773
rect 11446 12736 11928 12764
rect 11446 12733 11458 12736
rect 11400 12727 11458 12733
rect 5994 12696 6000 12708
rect 5675 12668 6000 12696
rect 5675 12665 5687 12668
rect 5629 12659 5687 12665
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 6546 12656 6552 12708
rect 6604 12696 6610 12708
rect 7146 12699 7204 12705
rect 7146 12696 7158 12699
rect 6604 12668 7158 12696
rect 6604 12656 6610 12668
rect 7146 12665 7158 12668
rect 7192 12665 7204 12699
rect 9950 12696 9956 12708
rect 9911 12668 9956 12696
rect 7146 12659 7204 12665
rect 9950 12656 9956 12668
rect 10008 12656 10014 12708
rect 10505 12699 10563 12705
rect 10505 12665 10517 12699
rect 10551 12696 10563 12699
rect 10962 12696 10968 12708
rect 10551 12668 10968 12696
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 3326 12628 3332 12640
rect 3287 12600 3332 12628
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 5902 12628 5908 12640
rect 5863 12600 5908 12628
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 8110 12588 8116 12640
rect 8168 12628 8174 12640
rect 8478 12628 8484 12640
rect 8168 12600 8484 12628
rect 8168 12588 8174 12600
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 9582 12628 9588 12640
rect 9456 12600 9588 12628
rect 9456 12588 9462 12600
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 11900 12637 11928 12736
rect 12596 12733 12608 12767
rect 12642 12764 12654 12767
rect 19864 12767 19922 12773
rect 12642 12736 12940 12764
rect 12642 12733 12654 12736
rect 12596 12727 12654 12733
rect 12912 12640 12940 12736
rect 19864 12733 19876 12767
rect 19910 12733 19922 12767
rect 19864 12727 19922 12733
rect 13722 12696 13728 12708
rect 13683 12668 13728 12696
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 15933 12699 15991 12705
rect 15933 12665 15945 12699
rect 15979 12665 15991 12699
rect 15933 12659 15991 12665
rect 10781 12631 10839 12637
rect 10781 12628 10793 12631
rect 9732 12600 10793 12628
rect 9732 12588 9738 12600
rect 10781 12597 10793 12600
rect 10827 12597 10839 12631
rect 10781 12591 10839 12597
rect 11885 12631 11943 12637
rect 11885 12597 11897 12631
rect 11931 12628 11943 12631
rect 11974 12628 11980 12640
rect 11931 12600 11980 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 12066 12588 12072 12640
rect 12124 12628 12130 12640
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 12124 12600 12173 12628
rect 12124 12588 12130 12600
rect 12161 12597 12173 12600
rect 12207 12597 12219 12631
rect 12161 12591 12219 12597
rect 12894 12588 12900 12640
rect 12952 12628 12958 12640
rect 12989 12631 13047 12637
rect 12989 12628 13001 12631
rect 12952 12600 13001 12628
rect 12952 12588 12958 12600
rect 12989 12597 13001 12600
rect 13035 12597 13047 12631
rect 12989 12591 13047 12597
rect 13265 12631 13323 12637
rect 13265 12597 13277 12631
rect 13311 12628 13323 12631
rect 13906 12628 13912 12640
rect 13311 12600 13912 12628
rect 13311 12597 13323 12600
rect 13265 12591 13323 12597
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 14550 12628 14556 12640
rect 14511 12600 14556 12628
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 15197 12631 15255 12637
rect 15197 12597 15209 12631
rect 15243 12628 15255 12631
rect 15948 12628 15976 12659
rect 16942 12656 16948 12708
rect 17000 12696 17006 12708
rect 17000 12668 17264 12696
rect 17000 12656 17006 12668
rect 17236 12640 17264 12668
rect 18414 12656 18420 12708
rect 18472 12696 18478 12708
rect 18472 12668 18517 12696
rect 18472 12656 18478 12668
rect 18690 12656 18696 12708
rect 18748 12696 18754 12708
rect 19879 12696 19907 12727
rect 19978 12724 19984 12776
rect 20036 12764 20042 12776
rect 20809 12767 20867 12773
rect 20809 12764 20821 12767
rect 20036 12736 20821 12764
rect 20036 12724 20042 12736
rect 20809 12733 20821 12736
rect 20855 12764 20867 12767
rect 20990 12764 20996 12776
rect 20855 12736 20996 12764
rect 20855 12733 20867 12736
rect 20809 12727 20867 12733
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 21450 12724 21456 12776
rect 21508 12764 21514 12776
rect 22278 12764 22284 12776
rect 21508 12736 22284 12764
rect 21508 12724 21514 12736
rect 22278 12724 22284 12736
rect 22336 12724 22342 12776
rect 22639 12773 22667 12804
rect 23109 12801 23121 12804
rect 23155 12832 23167 12835
rect 23155 12804 25151 12832
rect 23155 12801 23167 12804
rect 23109 12795 23167 12801
rect 22624 12767 22682 12773
rect 22624 12733 22636 12767
rect 22670 12733 22682 12767
rect 22624 12727 22682 12733
rect 24096 12767 24154 12773
rect 24096 12733 24108 12767
rect 24142 12764 24154 12767
rect 24946 12764 24952 12776
rect 24142 12736 24952 12764
rect 24142 12733 24154 12736
rect 24096 12727 24154 12733
rect 24946 12724 24952 12736
rect 25004 12724 25010 12776
rect 25123 12773 25151 12804
rect 25108 12767 25166 12773
rect 25108 12733 25120 12767
rect 25154 12764 25166 12767
rect 25608 12764 25636 12860
rect 25154 12736 25636 12764
rect 25154 12733 25166 12736
rect 25108 12727 25166 12733
rect 18748 12668 19907 12696
rect 21171 12699 21229 12705
rect 18748 12656 18754 12668
rect 21171 12665 21183 12699
rect 21217 12665 21229 12699
rect 22830 12696 22836 12708
rect 21171 12659 21229 12665
rect 22296 12668 22836 12696
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 15243 12600 16865 12628
rect 15243 12597 15255 12600
rect 15197 12591 15255 12597
rect 16853 12597 16865 12600
rect 16899 12628 16911 12631
rect 17034 12628 17040 12640
rect 16899 12600 17040 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 17218 12628 17224 12640
rect 17179 12600 17224 12628
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17865 12631 17923 12637
rect 17865 12597 17877 12631
rect 17911 12628 17923 12631
rect 18432 12628 18460 12656
rect 19245 12631 19303 12637
rect 19245 12628 19257 12631
rect 17911 12600 19257 12628
rect 17911 12597 17923 12600
rect 17865 12591 17923 12597
rect 19245 12597 19257 12600
rect 19291 12597 19303 12631
rect 19245 12591 19303 12597
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 19935 12631 19993 12637
rect 19935 12628 19947 12631
rect 19392 12600 19947 12628
rect 19392 12588 19398 12600
rect 19935 12597 19947 12600
rect 19981 12597 19993 12631
rect 19935 12591 19993 12597
rect 20717 12631 20775 12637
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 21186 12628 21214 12659
rect 22296 12640 22324 12668
rect 22830 12656 22836 12668
rect 22888 12696 22894 12708
rect 23385 12699 23443 12705
rect 23385 12696 23397 12699
rect 22888 12668 23397 12696
rect 22888 12656 22894 12668
rect 23385 12665 23397 12668
rect 23431 12665 23443 12699
rect 23385 12659 23443 12665
rect 21266 12628 21272 12640
rect 20763 12600 21272 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 21729 12631 21787 12637
rect 21729 12597 21741 12631
rect 21775 12628 21787 12631
rect 22278 12628 22284 12640
rect 21775 12600 22284 12628
rect 21775 12597 21787 12600
rect 21729 12591 21787 12597
rect 22278 12588 22284 12600
rect 22336 12588 22342 12640
rect 22554 12588 22560 12640
rect 22612 12628 22618 12640
rect 22695 12631 22753 12637
rect 22695 12628 22707 12631
rect 22612 12600 22707 12628
rect 22612 12588 22618 12600
rect 22695 12597 22707 12600
rect 22741 12597 22753 12631
rect 22695 12591 22753 12597
rect 23658 12588 23664 12640
rect 23716 12628 23722 12640
rect 24167 12631 24225 12637
rect 24167 12628 24179 12631
rect 23716 12600 24179 12628
rect 23716 12588 23722 12600
rect 24167 12597 24179 12600
rect 24213 12597 24225 12631
rect 24167 12591 24225 12597
rect 24581 12631 24639 12637
rect 24581 12597 24593 12631
rect 24627 12628 24639 12631
rect 24762 12628 24768 12640
rect 24627 12600 24768 12628
rect 24627 12597 24639 12600
rect 24581 12591 24639 12597
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 3970 12424 3976 12436
rect 2004 12396 3976 12424
rect 2004 12384 2010 12396
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 4157 12427 4215 12433
rect 4157 12424 4169 12427
rect 4120 12396 4169 12424
rect 4120 12384 4126 12396
rect 4157 12393 4169 12396
rect 4203 12393 4215 12427
rect 4157 12387 4215 12393
rect 6546 12384 6552 12436
rect 6604 12424 6610 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6604 12396 6929 12424
rect 6604 12384 6610 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 9858 12424 9864 12436
rect 9819 12396 9864 12424
rect 6917 12387 6975 12393
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10008 12396 10241 12424
rect 10008 12384 10014 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 12434 12424 12440 12436
rect 12395 12396 12440 12424
rect 10229 12387 10287 12393
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 13449 12427 13507 12433
rect 13449 12393 13461 12427
rect 13495 12424 13507 12427
rect 13722 12424 13728 12436
rect 13495 12396 13728 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 16390 12424 16396 12436
rect 16351 12396 16396 12424
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 18141 12427 18199 12433
rect 18141 12393 18153 12427
rect 18187 12424 18199 12427
rect 18230 12424 18236 12436
rect 18187 12396 18236 12424
rect 18187 12393 18199 12396
rect 18141 12387 18199 12393
rect 18230 12384 18236 12396
rect 18288 12384 18294 12436
rect 18506 12424 18512 12436
rect 18419 12396 18512 12424
rect 18506 12384 18512 12396
rect 18564 12424 18570 12436
rect 19334 12424 19340 12436
rect 18564 12396 19340 12424
rect 18564 12384 18570 12396
rect 19334 12384 19340 12396
rect 19392 12384 19398 12436
rect 20806 12384 20812 12436
rect 20864 12424 20870 12436
rect 21082 12424 21088 12436
rect 20864 12396 21088 12424
rect 20864 12384 20870 12396
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 21266 12424 21272 12436
rect 21227 12396 21272 12424
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 21818 12424 21824 12436
rect 21779 12396 21824 12424
rect 21818 12384 21824 12396
rect 21876 12384 21882 12436
rect 22094 12424 22100 12436
rect 22055 12396 22100 12424
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 22278 12384 22284 12436
rect 22336 12424 22342 12436
rect 22336 12396 22876 12424
rect 22336 12384 22342 12396
rect 2700 12328 4200 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1486 12288 1492 12300
rect 1443 12260 1492 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1486 12248 1492 12260
rect 1544 12248 1550 12300
rect 2314 12248 2320 12300
rect 2372 12288 2378 12300
rect 2700 12297 2728 12328
rect 2685 12291 2743 12297
rect 2685 12288 2697 12291
rect 2372 12260 2697 12288
rect 2372 12248 2378 12260
rect 2685 12257 2697 12260
rect 2731 12257 2743 12291
rect 2866 12288 2872 12300
rect 2827 12260 2872 12288
rect 2685 12251 2743 12257
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 4062 12288 4068 12300
rect 4023 12260 4068 12288
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4172 12288 4200 12328
rect 4246 12316 4252 12368
rect 4304 12356 4310 12368
rect 4522 12356 4528 12368
rect 4304 12328 4528 12356
rect 4304 12316 4310 12328
rect 4522 12316 4528 12328
rect 4580 12356 4586 12368
rect 6365 12359 6423 12365
rect 4580 12328 6132 12356
rect 4580 12316 4586 12328
rect 4430 12288 4436 12300
rect 4172 12260 4436 12288
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 4632 12297 4660 12328
rect 6104 12300 6132 12328
rect 6365 12325 6377 12359
rect 6411 12356 6423 12359
rect 6822 12356 6828 12368
rect 6411 12328 6828 12356
rect 6411 12325 6423 12328
rect 6365 12319 6423 12325
rect 6822 12316 6828 12328
rect 6880 12356 6886 12368
rect 7193 12359 7251 12365
rect 7193 12356 7205 12359
rect 6880 12328 7205 12356
rect 6880 12316 6886 12328
rect 7193 12325 7205 12328
rect 7239 12325 7251 12359
rect 7193 12319 7251 12325
rect 8757 12359 8815 12365
rect 8757 12325 8769 12359
rect 8803 12356 8815 12359
rect 9674 12356 9680 12368
rect 8803 12328 9680 12356
rect 8803 12325 8815 12328
rect 8757 12319 8815 12325
rect 9674 12316 9680 12328
rect 9732 12316 9738 12368
rect 10689 12359 10747 12365
rect 10689 12325 10701 12359
rect 10735 12356 10747 12359
rect 10870 12356 10876 12368
rect 10735 12328 10876 12356
rect 10735 12325 10747 12328
rect 10689 12319 10747 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 12158 12316 12164 12368
rect 12216 12356 12222 12368
rect 12850 12359 12908 12365
rect 12850 12356 12862 12359
rect 12216 12328 12862 12356
rect 12216 12316 12222 12328
rect 12850 12325 12862 12328
rect 12896 12325 12908 12359
rect 12850 12319 12908 12325
rect 15378 12316 15384 12368
rect 15436 12356 15442 12368
rect 15473 12359 15531 12365
rect 15473 12356 15485 12359
rect 15436 12328 15485 12356
rect 15436 12316 15442 12328
rect 15473 12325 15485 12328
rect 15519 12325 15531 12359
rect 15473 12319 15531 12325
rect 16025 12359 16083 12365
rect 16025 12325 16037 12359
rect 16071 12356 16083 12359
rect 16114 12356 16120 12368
rect 16071 12328 16120 12356
rect 16071 12325 16083 12328
rect 16025 12319 16083 12325
rect 16114 12316 16120 12328
rect 16172 12316 16178 12368
rect 16942 12316 16948 12368
rect 17000 12356 17006 12368
rect 17542 12359 17600 12365
rect 17542 12356 17554 12359
rect 17000 12328 17554 12356
rect 17000 12316 17006 12328
rect 17542 12325 17554 12328
rect 17588 12325 17600 12359
rect 18782 12356 18788 12368
rect 18743 12328 18788 12356
rect 17542 12319 17600 12325
rect 18782 12316 18788 12328
rect 18840 12316 18846 12368
rect 19426 12356 19432 12368
rect 19387 12328 19432 12356
rect 19426 12316 19432 12328
rect 19484 12316 19490 12368
rect 20530 12316 20536 12368
rect 20588 12356 20594 12368
rect 20990 12356 20996 12368
rect 20588 12328 20996 12356
rect 20588 12316 20594 12328
rect 20990 12316 20996 12328
rect 21048 12316 21054 12368
rect 22554 12316 22560 12368
rect 22612 12356 22618 12368
rect 22848 12365 22876 12396
rect 23198 12384 23204 12436
rect 23256 12424 23262 12436
rect 23842 12424 23848 12436
rect 23256 12396 23848 12424
rect 23256 12384 23262 12396
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 22741 12359 22799 12365
rect 22741 12356 22753 12359
rect 22612 12328 22753 12356
rect 22612 12316 22618 12328
rect 22741 12325 22753 12328
rect 22787 12325 22799 12359
rect 22741 12319 22799 12325
rect 22833 12359 22891 12365
rect 22833 12325 22845 12359
rect 22879 12325 22891 12359
rect 22833 12319 22891 12325
rect 4617 12291 4675 12297
rect 4617 12257 4629 12291
rect 4663 12257 4675 12291
rect 4617 12251 4675 12257
rect 5442 12248 5448 12300
rect 5500 12288 5506 12300
rect 5629 12291 5687 12297
rect 5629 12288 5641 12291
rect 5500 12260 5641 12288
rect 5500 12248 5506 12260
rect 5629 12257 5641 12260
rect 5675 12257 5687 12291
rect 6086 12288 6092 12300
rect 6047 12260 6092 12288
rect 5629 12251 5687 12257
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 8294 12288 8300 12300
rect 8076 12260 8300 12288
rect 8076 12248 8082 12260
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 8570 12288 8576 12300
rect 8531 12260 8576 12288
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 19981 12291 20039 12297
rect 19981 12257 19993 12291
rect 20027 12288 20039 12291
rect 21634 12288 21640 12300
rect 20027 12260 21640 12288
rect 20027 12257 20039 12260
rect 19981 12251 20039 12257
rect 21634 12248 21640 12260
rect 21692 12248 21698 12300
rect 24489 12291 24547 12297
rect 24489 12257 24501 12291
rect 24535 12288 24547 12291
rect 24578 12288 24584 12300
rect 24535 12260 24584 12288
rect 24535 12257 24547 12260
rect 24489 12251 24547 12257
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 24673 12291 24731 12297
rect 24673 12257 24685 12291
rect 24719 12288 24731 12291
rect 25406 12288 25412 12300
rect 24719 12260 25412 12288
rect 24719 12257 24731 12260
rect 24673 12251 24731 12257
rect 25406 12248 25412 12260
rect 25464 12248 25470 12300
rect 3142 12220 3148 12232
rect 3103 12192 3148 12220
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12220 3939 12223
rect 4338 12220 4344 12232
rect 3927 12192 4344 12220
rect 3927 12189 3939 12192
rect 3881 12183 3939 12189
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6822 12220 6828 12232
rect 5960 12192 6828 12220
rect 5960 12180 5966 12192
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 10778 12220 10784 12232
rect 10643 12192 10784 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 10962 12220 10968 12232
rect 10923 12192 10968 12220
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12220 12587 12223
rect 13078 12220 13084 12232
rect 12575 12192 13084 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 13078 12180 13084 12192
rect 13136 12180 13142 12232
rect 14090 12180 14096 12232
rect 14148 12220 14154 12232
rect 14826 12220 14832 12232
rect 14148 12192 14832 12220
rect 14148 12180 14154 12192
rect 14826 12180 14832 12192
rect 14884 12220 14890 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 14884 12192 15393 12220
rect 14884 12180 14890 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 17221 12223 17279 12229
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 17770 12220 17776 12232
rect 17267 12192 17776 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 19337 12223 19395 12229
rect 19337 12189 19349 12223
rect 19383 12220 19395 12223
rect 20070 12220 20076 12232
rect 19383 12192 20076 12220
rect 19383 12189 19395 12192
rect 19337 12183 19395 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 20898 12220 20904 12232
rect 20859 12192 20904 12220
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 22922 12180 22928 12232
rect 22980 12220 22986 12232
rect 23017 12223 23075 12229
rect 23017 12220 23029 12223
rect 22980 12192 23029 12220
rect 22980 12180 22986 12192
rect 23017 12189 23029 12192
rect 23063 12189 23075 12223
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 23017 12183 23075 12189
rect 23446 12192 24777 12220
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 4154 12152 4160 12164
rect 1627 12124 4160 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 4154 12112 4160 12124
rect 4212 12152 4218 12164
rect 4522 12152 4528 12164
rect 4212 12124 4528 12152
rect 4212 12112 4218 12124
rect 4522 12112 4528 12124
rect 4580 12152 4586 12164
rect 4890 12152 4896 12164
rect 4580 12124 4896 12152
rect 4580 12112 4586 12124
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 6730 12112 6736 12164
rect 6788 12152 6794 12164
rect 13722 12152 13728 12164
rect 6788 12124 13728 12152
rect 6788 12112 6794 12124
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 22370 12112 22376 12164
rect 22428 12152 22434 12164
rect 23446 12152 23474 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 22428 12124 23474 12152
rect 22428 12112 22434 12124
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2225 12087 2283 12093
rect 2225 12084 2237 12087
rect 2096 12056 2237 12084
rect 2096 12044 2102 12056
rect 2225 12053 2237 12056
rect 2271 12053 2283 12087
rect 2225 12047 2283 12053
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4672 12056 5089 12084
rect 4672 12044 4678 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5077 12047 5135 12053
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 8018 12084 8024 12096
rect 7975 12056 8024 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 13170 12084 13176 12096
rect 12952 12056 13176 12084
rect 12952 12044 12958 12056
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 14182 12084 14188 12096
rect 14143 12056 14188 12084
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 20714 12084 20720 12096
rect 20675 12056 20720 12084
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 23661 12087 23719 12093
rect 23661 12084 23673 12087
rect 23624 12056 23673 12084
rect 23624 12044 23630 12056
rect 23661 12053 23673 12056
rect 23707 12053 23719 12087
rect 23661 12047 23719 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2225 11883 2283 11889
rect 2225 11849 2237 11883
rect 2271 11880 2283 11883
rect 2314 11880 2320 11892
rect 2271 11852 2320 11880
rect 2271 11849 2283 11852
rect 2225 11843 2283 11849
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11880 3295 11883
rect 3418 11880 3424 11892
rect 3283 11852 3424 11880
rect 3283 11849 3295 11852
rect 3237 11843 3295 11849
rect 3418 11840 3424 11852
rect 3476 11840 3482 11892
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 5500 11852 5641 11880
rect 5500 11840 5506 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 7009 11883 7067 11889
rect 7009 11849 7021 11883
rect 7055 11880 7067 11883
rect 7098 11880 7104 11892
rect 7055 11852 7104 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 8941 11883 8999 11889
rect 8941 11880 8953 11883
rect 8352 11852 8953 11880
rect 8352 11840 8358 11852
rect 8941 11849 8953 11852
rect 8987 11880 8999 11883
rect 10597 11883 10655 11889
rect 10597 11880 10609 11883
rect 8987 11852 10609 11880
rect 8987 11849 8999 11852
rect 8941 11843 8999 11849
rect 10597 11849 10609 11852
rect 10643 11849 10655 11883
rect 10597 11843 10655 11849
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 10836 11852 11161 11880
rect 10836 11840 10842 11852
rect 11149 11849 11161 11852
rect 11195 11849 11207 11883
rect 11149 11843 11207 11849
rect 16945 11883 17003 11889
rect 16945 11849 16957 11883
rect 16991 11880 17003 11883
rect 17310 11880 17316 11892
rect 16991 11852 17316 11880
rect 16991 11849 17003 11852
rect 16945 11843 17003 11849
rect 7742 11772 7748 11824
rect 7800 11812 7806 11824
rect 8481 11815 8539 11821
rect 8481 11812 8493 11815
rect 7800 11784 8493 11812
rect 7800 11772 7806 11784
rect 8481 11781 8493 11784
rect 8527 11812 8539 11815
rect 10686 11812 10692 11824
rect 8527 11784 10692 11812
rect 8527 11781 8539 11784
rect 8481 11775 8539 11781
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 11517 11815 11575 11821
rect 11517 11781 11529 11815
rect 11563 11812 11575 11815
rect 12342 11812 12348 11824
rect 11563 11784 12348 11812
rect 11563 11781 11575 11784
rect 11517 11775 11575 11781
rect 2869 11747 2927 11753
rect 2869 11744 2881 11747
rect 2332 11716 2881 11744
rect 2332 11685 2360 11716
rect 2869 11713 2881 11716
rect 2915 11744 2927 11747
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 2915 11716 4813 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 4801 11713 4813 11716
rect 4847 11744 4859 11747
rect 9585 11747 9643 11753
rect 4847 11716 8616 11744
rect 4847 11713 4859 11716
rect 4801 11707 4859 11713
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11645 2375 11679
rect 2317 11639 2375 11645
rect 2406 11636 2412 11688
rect 2464 11676 2470 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 2464 11648 3341 11676
rect 2464 11636 2470 11648
rect 3329 11645 3341 11648
rect 3375 11676 3387 11679
rect 3418 11676 3424 11688
rect 3375 11648 3424 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 4338 11676 4344 11688
rect 4299 11648 4344 11676
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 4433 11679 4491 11685
rect 4433 11645 4445 11679
rect 4479 11645 4491 11679
rect 4614 11676 4620 11688
rect 4575 11648 4620 11676
rect 4433 11639 4491 11645
rect 3789 11611 3847 11617
rect 3789 11608 3801 11611
rect 1596 11580 3801 11608
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 1596 11549 1624 11580
rect 3789 11577 3801 11580
rect 3835 11608 3847 11611
rect 4062 11608 4068 11620
rect 3835 11580 4068 11608
rect 3835 11577 3847 11580
rect 3789 11571 3847 11577
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 1544 11512 1593 11540
rect 1544 11500 1550 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 1581 11503 1639 11509
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 2590 11540 2596 11552
rect 2547 11512 2596 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3476 11512 3525 11540
rect 3476 11500 3482 11512
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 3513 11503 3571 11509
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 4448 11540 4476 11639
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 5592 11648 6837 11676
rect 5592 11636 5598 11648
rect 6825 11645 6837 11648
rect 6871 11676 6883 11679
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 6871 11648 7297 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 8588 11676 8616 11716
rect 9585 11713 9597 11747
rect 9631 11744 9643 11747
rect 9858 11744 9864 11756
rect 9631 11716 9864 11744
rect 9631 11713 9643 11716
rect 9585 11707 9643 11713
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11744 10655 11747
rect 11532 11744 11560 11775
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 16960 11812 16988 11843
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 21542 11840 21548 11892
rect 21600 11880 21606 11892
rect 21637 11883 21695 11889
rect 21637 11880 21649 11883
rect 21600 11852 21649 11880
rect 21600 11840 21606 11852
rect 21637 11849 21649 11852
rect 21683 11849 21695 11883
rect 22278 11880 22284 11892
rect 22239 11852 22284 11880
rect 21637 11843 21695 11849
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 24670 11880 24676 11892
rect 23446 11852 24676 11880
rect 15948 11784 16988 11812
rect 18417 11815 18475 11821
rect 10643 11716 11560 11744
rect 10643 11713 10655 11716
rect 10597 11707 10655 11713
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11882 11744 11888 11756
rect 11664 11716 11888 11744
rect 11664 11704 11670 11716
rect 11882 11704 11888 11716
rect 11940 11744 11946 11756
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 11940 11716 13553 11744
rect 11940 11704 11946 11716
rect 11333 11679 11391 11685
rect 11333 11676 11345 11679
rect 8588 11648 11345 11676
rect 7285 11639 7343 11645
rect 11333 11645 11345 11648
rect 11379 11676 11391 11679
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11379 11648 11805 11676
rect 11379 11645 11391 11648
rect 11333 11639 11391 11645
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 12802 11676 12808 11688
rect 12763 11648 12808 11676
rect 11793 11639 11851 11645
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 13004 11685 13032 11716
rect 13541 11713 13553 11716
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11744 14151 11747
rect 14182 11744 14188 11756
rect 14139 11716 14188 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11645 13047 11679
rect 13556 11676 13584 11707
rect 14182 11704 14188 11716
rect 14240 11744 14246 11756
rect 15746 11744 15752 11756
rect 14240 11716 15752 11744
rect 14240 11704 14246 11716
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 15948 11753 15976 11784
rect 18417 11781 18429 11815
rect 18463 11812 18475 11815
rect 19426 11812 19432 11824
rect 18463 11784 19432 11812
rect 18463 11781 18475 11784
rect 18417 11775 18475 11781
rect 19426 11772 19432 11784
rect 19484 11812 19490 11824
rect 19797 11815 19855 11821
rect 19797 11812 19809 11815
rect 19484 11784 19809 11812
rect 19484 11772 19490 11784
rect 19797 11781 19809 11784
rect 19843 11781 19855 11815
rect 19797 11775 19855 11781
rect 20070 11772 20076 11824
rect 20128 11812 20134 11824
rect 22603 11815 22661 11821
rect 22603 11812 22615 11815
rect 20128 11784 22615 11812
rect 20128 11772 20134 11784
rect 22603 11781 22615 11784
rect 22649 11781 22661 11815
rect 22603 11775 22661 11781
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 16172 11716 16221 11744
rect 16172 11704 16178 11716
rect 16209 11713 16221 11716
rect 16255 11713 16267 11747
rect 20714 11744 20720 11756
rect 20627 11716 20720 11744
rect 16209 11707 16267 11713
rect 20714 11704 20720 11716
rect 20772 11744 20778 11756
rect 22094 11744 22100 11756
rect 20772 11716 22100 11744
rect 20772 11704 20778 11716
rect 22094 11704 22100 11716
rect 22152 11704 22158 11756
rect 22922 11744 22928 11756
rect 22883 11716 22928 11744
rect 22922 11704 22928 11716
rect 22980 11704 22986 11756
rect 14734 11676 14740 11688
rect 13556 11648 14740 11676
rect 12989 11639 13047 11645
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15013 11679 15071 11685
rect 15013 11645 15025 11679
rect 15059 11676 15071 11679
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 15059 11648 15669 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 15657 11645 15669 11648
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 18966 11676 18972 11688
rect 18923 11648 18972 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 6086 11608 6092 11620
rect 5999 11580 6092 11608
rect 6086 11568 6092 11580
rect 6144 11608 6150 11620
rect 6144 11580 7696 11608
rect 6144 11568 6150 11580
rect 4522 11540 4528 11552
rect 4295 11512 4528 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 7668 11549 7696 11580
rect 7742 11568 7748 11620
rect 7800 11608 7806 11620
rect 7929 11611 7987 11617
rect 7929 11608 7941 11611
rect 7800 11580 7941 11608
rect 7800 11568 7806 11580
rect 7929 11577 7941 11580
rect 7975 11577 7987 11611
rect 7929 11571 7987 11577
rect 8018 11568 8024 11620
rect 8076 11608 8082 11620
rect 9906 11611 9964 11617
rect 9906 11608 9918 11611
rect 8076 11580 8121 11608
rect 9416 11580 9918 11608
rect 8076 11568 8082 11580
rect 9416 11552 9444 11580
rect 9906 11577 9918 11580
rect 9952 11608 9964 11611
rect 12158 11608 12164 11620
rect 9952 11580 12164 11608
rect 9952 11577 9964 11580
rect 9906 11571 9964 11577
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 13262 11608 13268 11620
rect 13223 11580 13268 11608
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 14414 11611 14472 11617
rect 14414 11608 14426 11611
rect 14200 11580 14426 11608
rect 14200 11552 14228 11580
rect 14414 11577 14426 11580
rect 14460 11577 14472 11611
rect 14414 11571 14472 11577
rect 7653 11543 7711 11549
rect 7653 11509 7665 11543
rect 7699 11540 7711 11543
rect 8570 11540 8576 11552
rect 7699 11512 8576 11540
rect 7699 11509 7711 11512
rect 7653 11503 7711 11509
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 9398 11540 9404 11552
rect 9359 11512 9404 11540
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 10870 11540 10876 11552
rect 10551 11512 10876 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 13906 11500 13912 11552
rect 13964 11540 13970 11552
rect 14001 11543 14059 11549
rect 14001 11540 14013 11543
rect 13964 11512 14013 11540
rect 13964 11500 13970 11512
rect 14001 11509 14013 11512
rect 14047 11540 14059 11543
rect 14182 11540 14188 11552
rect 14047 11512 14188 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 15286 11540 15292 11552
rect 15247 11512 15292 11540
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 15672 11540 15700 11639
rect 18966 11636 18972 11648
rect 19024 11636 19030 11688
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 21913 11679 21971 11685
rect 21913 11676 21925 11679
rect 20956 11648 21925 11676
rect 20956 11636 20962 11648
rect 21913 11645 21925 11648
rect 21959 11645 21971 11679
rect 21913 11639 21971 11645
rect 22532 11679 22590 11685
rect 22532 11645 22544 11679
rect 22578 11676 22590 11679
rect 22940 11676 22968 11704
rect 22578 11648 22968 11676
rect 22578 11645 22590 11648
rect 22532 11639 22590 11645
rect 23014 11636 23020 11688
rect 23072 11676 23078 11688
rect 23446 11676 23474 11852
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 23934 11772 23940 11824
rect 23992 11812 23998 11824
rect 25409 11815 25467 11821
rect 25409 11812 25421 11815
rect 23992 11784 25421 11812
rect 23992 11772 23998 11784
rect 25409 11781 25421 11784
rect 25455 11781 25467 11815
rect 25409 11775 25467 11781
rect 23072 11648 23474 11676
rect 23072 11636 23078 11648
rect 23566 11636 23572 11688
rect 23624 11676 23630 11688
rect 23661 11679 23719 11685
rect 23661 11676 23673 11679
rect 23624 11648 23673 11676
rect 23624 11636 23630 11648
rect 23661 11645 23673 11648
rect 23707 11645 23719 11679
rect 23661 11639 23719 11645
rect 24121 11679 24179 11685
rect 24121 11645 24133 11679
rect 24167 11645 24179 11679
rect 24121 11639 24179 11645
rect 25225 11679 25283 11685
rect 25225 11645 25237 11679
rect 25271 11676 25283 11679
rect 25498 11676 25504 11688
rect 25271 11648 25504 11676
rect 25271 11645 25283 11648
rect 25225 11639 25283 11645
rect 16025 11611 16083 11617
rect 16025 11577 16037 11611
rect 16071 11577 16083 11611
rect 18693 11611 18751 11617
rect 18693 11608 18705 11611
rect 16025 11571 16083 11577
rect 17236 11580 18705 11608
rect 16040 11540 16068 11571
rect 15672 11512 16068 11540
rect 16942 11500 16948 11552
rect 17000 11540 17006 11552
rect 17236 11549 17264 11580
rect 18693 11577 18705 11580
rect 18739 11608 18751 11611
rect 19198 11611 19256 11617
rect 19198 11608 19210 11611
rect 18739 11580 19210 11608
rect 18739 11577 18751 11580
rect 18693 11571 18751 11577
rect 19198 11577 19210 11580
rect 19244 11608 19256 11611
rect 19518 11608 19524 11620
rect 19244 11580 19524 11608
rect 19244 11577 19256 11580
rect 19198 11571 19256 11577
rect 19518 11568 19524 11580
rect 19576 11608 19582 11620
rect 20165 11611 20223 11617
rect 20165 11608 20177 11611
rect 19576 11580 20177 11608
rect 19576 11568 19582 11580
rect 20165 11577 20177 11580
rect 20211 11608 20223 11611
rect 20533 11611 20591 11617
rect 20533 11608 20545 11611
rect 20211 11580 20545 11608
rect 20211 11577 20223 11580
rect 20165 11571 20223 11577
rect 20533 11577 20545 11580
rect 20579 11608 20591 11611
rect 21038 11611 21096 11617
rect 21038 11608 21050 11611
rect 20579 11580 21050 11608
rect 20579 11577 20591 11580
rect 20533 11571 20591 11577
rect 21038 11577 21050 11580
rect 21084 11608 21096 11611
rect 21266 11608 21272 11620
rect 21084 11580 21272 11608
rect 21084 11577 21096 11580
rect 21038 11571 21096 11577
rect 21266 11568 21272 11580
rect 21324 11568 21330 11620
rect 23106 11568 23112 11620
rect 23164 11608 23170 11620
rect 23385 11611 23443 11617
rect 23385 11608 23397 11611
rect 23164 11580 23397 11608
rect 23164 11568 23170 11580
rect 23385 11577 23397 11580
rect 23431 11577 23443 11611
rect 23385 11571 23443 11577
rect 23474 11568 23480 11620
rect 23532 11608 23538 11620
rect 24136 11608 24164 11639
rect 25498 11636 25504 11648
rect 25556 11676 25562 11688
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 25556 11648 25789 11676
rect 25556 11636 25562 11648
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 23532 11580 24164 11608
rect 23532 11568 23538 11580
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 17000 11512 17233 11540
rect 17000 11500 17006 11512
rect 17221 11509 17233 11512
rect 17267 11509 17279 11543
rect 17221 11503 17279 11509
rect 17681 11543 17739 11549
rect 17681 11509 17693 11543
rect 17727 11540 17739 11543
rect 17770 11540 17776 11552
rect 17727 11512 17776 11540
rect 17727 11509 17739 11512
rect 17681 11503 17739 11509
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 21174 11500 21180 11552
rect 21232 11540 21238 11552
rect 21818 11540 21824 11552
rect 21232 11512 21824 11540
rect 21232 11500 21238 11512
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 23750 11540 23756 11552
rect 23711 11512 23756 11540
rect 23750 11500 23756 11512
rect 23808 11500 23814 11552
rect 25133 11543 25191 11549
rect 25133 11509 25145 11543
rect 25179 11540 25191 11543
rect 25406 11540 25412 11552
rect 25179 11512 25412 11540
rect 25179 11509 25191 11512
rect 25133 11503 25191 11509
rect 25406 11500 25412 11512
rect 25464 11500 25470 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 2406 11336 2412 11348
rect 1627 11308 2412 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 3326 11296 3332 11348
rect 3384 11336 3390 11348
rect 4893 11339 4951 11345
rect 4893 11336 4905 11339
rect 3384 11308 4905 11336
rect 3384 11296 3390 11308
rect 4893 11305 4905 11308
rect 4939 11305 4951 11339
rect 4893 11299 4951 11305
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 7650 11336 7656 11348
rect 6604 11308 7656 11336
rect 6604 11296 6610 11308
rect 7650 11296 7656 11308
rect 7708 11336 7714 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 7708 11308 7941 11336
rect 7708 11296 7714 11308
rect 7929 11305 7941 11308
rect 7975 11305 7987 11339
rect 7929 11299 7987 11305
rect 8018 11296 8024 11348
rect 8076 11336 8082 11348
rect 8481 11339 8539 11345
rect 8481 11336 8493 11339
rect 8076 11308 8493 11336
rect 8076 11296 8082 11308
rect 8481 11305 8493 11308
rect 8527 11305 8539 11339
rect 12802 11336 12808 11348
rect 12763 11308 12808 11336
rect 8481 11299 8539 11305
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13078 11336 13084 11348
rect 13039 11308 13084 11336
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11305 13783 11339
rect 13725 11299 13783 11305
rect 14277 11339 14335 11345
rect 14277 11305 14289 11339
rect 14323 11336 14335 11339
rect 15286 11336 15292 11348
rect 14323 11308 15292 11336
rect 14323 11305 14335 11308
rect 14277 11299 14335 11305
rect 2038 11228 2044 11280
rect 2096 11268 2102 11280
rect 3789 11271 3847 11277
rect 3789 11268 3801 11271
rect 2096 11240 3801 11268
rect 2096 11228 2102 11240
rect 3789 11237 3801 11240
rect 3835 11268 3847 11271
rect 4338 11268 4344 11280
rect 3835 11240 4344 11268
rect 3835 11237 3847 11240
rect 3789 11231 3847 11237
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 4798 11228 4804 11280
rect 4856 11268 4862 11280
rect 7377 11271 7435 11277
rect 7377 11268 7389 11271
rect 4856 11240 7389 11268
rect 4856 11228 4862 11240
rect 7377 11237 7389 11240
rect 7423 11268 7435 11271
rect 7742 11268 7748 11280
rect 7423 11240 7748 11268
rect 7423 11237 7435 11240
rect 7377 11231 7435 11237
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 10870 11268 10876 11280
rect 10831 11240 10876 11268
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 13740 11268 13768 11299
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 18233 11339 18291 11345
rect 18233 11305 18245 11339
rect 18279 11336 18291 11339
rect 18414 11336 18420 11348
rect 18279 11308 18420 11336
rect 18279 11305 18291 11308
rect 18233 11299 18291 11305
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 18601 11339 18659 11345
rect 18601 11305 18613 11339
rect 18647 11336 18659 11339
rect 20070 11336 20076 11348
rect 18647 11308 20076 11336
rect 18647 11305 18659 11308
rect 18601 11299 18659 11305
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 20441 11339 20499 11345
rect 20441 11336 20453 11339
rect 20404 11308 20453 11336
rect 20404 11296 20410 11308
rect 20441 11305 20453 11308
rect 20487 11305 20499 11339
rect 20441 11299 20499 11305
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20956 11308 21005 11336
rect 20956 11296 20962 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 22554 11296 22560 11348
rect 22612 11336 22618 11348
rect 22649 11339 22707 11345
rect 22649 11336 22661 11339
rect 22612 11308 22661 11336
rect 22612 11296 22618 11308
rect 22649 11305 22661 11308
rect 22695 11305 22707 11339
rect 24946 11336 24952 11348
rect 24907 11308 24952 11336
rect 22649 11299 22707 11305
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 14182 11268 14188 11280
rect 13740 11240 14188 11268
rect 14182 11228 14188 11240
rect 14240 11228 14246 11280
rect 14826 11228 14832 11280
rect 14884 11268 14890 11280
rect 15013 11271 15071 11277
rect 15013 11268 15025 11271
rect 14884 11240 15025 11268
rect 14884 11228 14890 11240
rect 15013 11237 15025 11240
rect 15059 11237 15071 11271
rect 15654 11268 15660 11280
rect 15615 11240 15660 11268
rect 15013 11231 15071 11237
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 16942 11228 16948 11280
rect 17000 11268 17006 11280
rect 17634 11271 17692 11277
rect 17634 11268 17646 11271
rect 17000 11240 17646 11268
rect 17000 11228 17006 11240
rect 17634 11237 17646 11240
rect 17680 11237 17692 11271
rect 19978 11268 19984 11280
rect 19939 11240 19984 11268
rect 17634 11231 17692 11237
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 23532 11240 23577 11268
rect 23532 11228 23538 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11169 1455 11203
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 1397 11163 1455 11169
rect 1412 11132 1440 11163
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2682 11200 2688 11212
rect 2643 11172 2688 11200
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 4246 11200 4252 11212
rect 4207 11172 4252 11200
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4430 11200 4436 11212
rect 4391 11172 4436 11200
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 4614 11160 4620 11212
rect 4672 11200 4678 11212
rect 4709 11203 4767 11209
rect 4709 11200 4721 11203
rect 4672 11172 4721 11200
rect 4672 11160 4678 11172
rect 4709 11169 4721 11172
rect 4755 11169 4767 11203
rect 4709 11163 4767 11169
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5224 11172 6009 11200
rect 5224 11160 5230 11172
rect 5997 11169 6009 11172
rect 6043 11200 6055 11203
rect 6362 11200 6368 11212
rect 6043 11172 6368 11200
rect 6043 11169 6055 11172
rect 5997 11163 6055 11169
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 8386 11200 8392 11212
rect 6503 11172 8392 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 1670 11132 1676 11144
rect 1412 11104 1676 11132
rect 1670 11092 1676 11104
rect 1728 11132 1734 11144
rect 2869 11135 2927 11141
rect 2869 11132 2881 11135
rect 1728 11104 2881 11132
rect 1728 11092 1734 11104
rect 2869 11101 2881 11104
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 5442 11092 5448 11144
rect 5500 11132 5506 11144
rect 6472 11132 6500 11163
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 8720 11172 9689 11200
rect 8720 11160 8726 11172
rect 9677 11169 9689 11172
rect 9723 11200 9735 11203
rect 10502 11200 10508 11212
rect 9723 11172 10508 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 12158 11160 12164 11212
rect 12216 11200 12222 11212
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 12216 11172 12265 11200
rect 12216 11160 12222 11172
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 13320 11172 13369 11200
rect 13320 11160 13326 11172
rect 13357 11169 13369 11172
rect 13403 11169 13415 11203
rect 19426 11200 19432 11212
rect 19387 11172 19432 11200
rect 13357 11163 13415 11169
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 19705 11203 19763 11209
rect 19705 11200 19717 11203
rect 19576 11172 19717 11200
rect 19576 11160 19582 11172
rect 19705 11169 19717 11172
rect 19751 11169 19763 11203
rect 20898 11200 20904 11212
rect 20859 11172 20904 11200
rect 19705 11163 19763 11169
rect 5500 11104 6500 11132
rect 6733 11135 6791 11141
rect 5500 11092 5506 11104
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 7190 11132 7196 11144
rect 6779 11104 7196 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 7190 11092 7196 11104
rect 7248 11132 7254 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7248 11104 7573 11132
rect 7248 11092 7254 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 11054 11132 11060 11144
rect 10827 11104 11060 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 15562 11132 15568 11144
rect 15523 11104 15568 11132
rect 15562 11092 15568 11104
rect 15620 11132 15626 11144
rect 16022 11132 16028 11144
rect 15620 11104 16028 11132
rect 15620 11092 15626 11104
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 19720 11132 19748 11163
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 21361 11203 21419 11209
rect 21361 11169 21373 11203
rect 21407 11169 21419 11203
rect 25130 11200 25136 11212
rect 25091 11172 25136 11200
rect 21361 11163 21419 11169
rect 21376 11132 21404 11163
rect 25130 11160 25136 11172
rect 25188 11160 25194 11212
rect 25317 11203 25375 11209
rect 25317 11169 25329 11203
rect 25363 11169 25375 11203
rect 25317 11163 25375 11169
rect 21542 11132 21548 11144
rect 19720 11104 21548 11132
rect 21542 11092 21548 11104
rect 21600 11092 21606 11144
rect 22002 11092 22008 11144
rect 22060 11092 22066 11144
rect 23385 11135 23443 11141
rect 23385 11101 23397 11135
rect 23431 11132 23443 11135
rect 23658 11132 23664 11144
rect 23431 11104 23664 11132
rect 23431 11101 23443 11104
rect 23385 11095 23443 11101
rect 23658 11092 23664 11104
rect 23716 11092 23722 11144
rect 23768 11104 24583 11132
rect 2498 11064 2504 11076
rect 2411 11036 2504 11064
rect 2498 11024 2504 11036
rect 2556 11064 2562 11076
rect 3513 11067 3571 11073
rect 3513 11064 3525 11067
rect 2556 11036 3525 11064
rect 2556 11024 2562 11036
rect 3513 11033 3525 11036
rect 3559 11064 3571 11067
rect 4062 11064 4068 11076
rect 3559 11036 4068 11064
rect 3559 11033 3571 11036
rect 3513 11027 3571 11033
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 4522 11064 4528 11076
rect 4483 11036 4528 11064
rect 4522 11024 4528 11036
rect 4580 11024 4586 11076
rect 10686 11024 10692 11076
rect 10744 11064 10750 11076
rect 11333 11067 11391 11073
rect 11333 11064 11345 11067
rect 10744 11036 11345 11064
rect 10744 11024 10750 11036
rect 11333 11033 11345 11036
rect 11379 11033 11391 11067
rect 11333 11027 11391 11033
rect 12161 11067 12219 11073
rect 12161 11033 12173 11067
rect 12207 11064 12219 11067
rect 12526 11064 12532 11076
rect 12207 11036 12532 11064
rect 12207 11033 12219 11036
rect 12161 11027 12219 11033
rect 12526 11024 12532 11036
rect 12584 11024 12590 11076
rect 16114 11064 16120 11076
rect 16075 11036 16120 11064
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 22020 11064 22048 11092
rect 23768 11064 23796 11104
rect 23934 11064 23940 11076
rect 22020 11036 23796 11064
rect 23895 11036 23940 11064
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 24555 11064 24583 11104
rect 24946 11092 24952 11144
rect 25004 11132 25010 11144
rect 25332 11132 25360 11163
rect 25004 11104 25360 11132
rect 25004 11092 25010 11104
rect 25314 11064 25320 11076
rect 24555 11036 25320 11064
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 1854 10996 1860 11008
rect 1815 10968 1860 10996
rect 1854 10956 1860 10968
rect 1912 10956 1918 11008
rect 2314 10996 2320 11008
rect 2275 10968 2320 10996
rect 2314 10956 2320 10968
rect 2372 10956 2378 11008
rect 9858 10996 9864 11008
rect 9819 10968 9864 10996
rect 9858 10956 9864 10968
rect 9916 10956 9922 11008
rect 12434 10996 12440 11008
rect 12395 10968 12440 10996
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 13630 10956 13636 11008
rect 13688 10996 13694 11008
rect 16666 10996 16672 11008
rect 13688 10968 16672 10996
rect 13688 10956 13694 10968
rect 16666 10956 16672 10968
rect 16724 10956 16730 11008
rect 18966 10996 18972 11008
rect 18927 10968 18972 10996
rect 18966 10956 18972 10968
rect 19024 10956 19030 11008
rect 22097 10999 22155 11005
rect 22097 10965 22109 10999
rect 22143 10996 22155 10999
rect 22186 10996 22192 11008
rect 22143 10968 22192 10996
rect 22143 10965 22155 10968
rect 22097 10959 22155 10965
rect 22186 10956 22192 10968
rect 22244 10956 22250 11008
rect 23842 10956 23848 11008
rect 23900 10996 23906 11008
rect 24305 10999 24363 11005
rect 24305 10996 24317 10999
rect 23900 10968 24317 10996
rect 23900 10956 23906 10968
rect 24305 10965 24317 10968
rect 24351 10965 24363 10999
rect 24305 10959 24363 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1670 10792 1676 10804
rect 1631 10764 1676 10792
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 2464 10764 3249 10792
rect 2464 10752 2470 10764
rect 3237 10761 3249 10764
rect 3283 10792 3295 10795
rect 3421 10795 3479 10801
rect 3421 10792 3433 10795
rect 3283 10764 3433 10792
rect 3283 10761 3295 10764
rect 3237 10755 3295 10761
rect 3421 10761 3433 10764
rect 3467 10761 3479 10795
rect 3421 10755 3479 10761
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 5537 10795 5595 10801
rect 5537 10792 5549 10795
rect 5500 10764 5549 10792
rect 5500 10752 5506 10764
rect 5537 10761 5549 10764
rect 5583 10761 5595 10795
rect 5537 10755 5595 10761
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6420 10764 6561 10792
rect 6420 10752 6426 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 7190 10792 7196 10804
rect 7151 10764 7196 10792
rect 6549 10755 6607 10761
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 7650 10792 7656 10804
rect 7611 10764 7656 10792
rect 7650 10752 7656 10764
rect 7708 10792 7714 10804
rect 9125 10795 9183 10801
rect 9125 10792 9137 10795
rect 7708 10764 9137 10792
rect 7708 10752 7714 10764
rect 9125 10761 9137 10764
rect 9171 10792 9183 10795
rect 9398 10792 9404 10804
rect 9171 10764 9404 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 10502 10792 10508 10804
rect 10463 10764 10508 10792
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 10870 10792 10876 10804
rect 10831 10764 10876 10792
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11241 10795 11299 10801
rect 11241 10761 11253 10795
rect 11287 10792 11299 10795
rect 11698 10792 11704 10804
rect 11287 10764 11704 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 12158 10792 12164 10804
rect 12119 10764 12164 10792
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 12492 10764 15945 10792
rect 12492 10752 12498 10764
rect 15933 10761 15945 10764
rect 15979 10792 15991 10795
rect 16758 10792 16764 10804
rect 15979 10764 16764 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 2317 10727 2375 10733
rect 2317 10693 2329 10727
rect 2363 10724 2375 10727
rect 2498 10724 2504 10736
rect 2363 10696 2504 10724
rect 2363 10693 2375 10696
rect 2317 10687 2375 10693
rect 2498 10684 2504 10696
rect 2556 10684 2562 10736
rect 6273 10727 6331 10733
rect 2976 10696 5764 10724
rect 2976 10665 3004 10696
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10625 3019 10659
rect 5074 10656 5080 10668
rect 2961 10619 3019 10625
rect 3068 10628 5080 10656
rect 2038 10548 2044 10600
rect 2096 10588 2102 10600
rect 2225 10591 2283 10597
rect 2225 10588 2237 10591
rect 2096 10560 2237 10588
rect 2096 10548 2102 10560
rect 2225 10557 2237 10560
rect 2271 10588 2283 10591
rect 2314 10588 2320 10600
rect 2271 10560 2320 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 3068 10588 3096 10628
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 2547 10560 3096 10588
rect 3697 10591 3755 10597
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 3743 10560 4353 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 4341 10557 4353 10560
rect 4387 10588 4399 10591
rect 4522 10588 4528 10600
rect 4387 10560 4528 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 2133 10523 2191 10529
rect 2133 10489 2145 10523
rect 2179 10520 2191 10523
rect 2516 10520 2544 10551
rect 4522 10548 4528 10560
rect 4580 10588 4586 10600
rect 5736 10597 5764 10696
rect 6273 10693 6285 10727
rect 6319 10724 6331 10727
rect 6914 10724 6920 10736
rect 6319 10696 6920 10724
rect 6319 10693 6331 10696
rect 6273 10687 6331 10693
rect 5721 10591 5779 10597
rect 4580 10560 4936 10588
rect 4580 10548 4586 10560
rect 2179 10492 2544 10520
rect 3421 10523 3479 10529
rect 2179 10489 2191 10492
rect 2133 10483 2191 10489
rect 3421 10489 3433 10523
rect 3467 10520 3479 10523
rect 4430 10520 4436 10532
rect 3467 10492 4436 10520
rect 3467 10489 3479 10492
rect 3421 10483 3479 10489
rect 4430 10480 4436 10492
rect 4488 10520 4494 10532
rect 4488 10492 4752 10520
rect 4488 10480 4494 10492
rect 4724 10464 4752 10492
rect 4908 10464 4936 10560
rect 5721 10557 5733 10591
rect 5767 10588 5779 10591
rect 6288 10588 6316 10687
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 8389 10727 8447 10733
rect 8389 10693 8401 10727
rect 8435 10724 8447 10727
rect 8478 10724 8484 10736
rect 8435 10696 8484 10724
rect 8435 10693 8447 10696
rect 8389 10687 8447 10693
rect 8478 10684 8484 10696
rect 8536 10724 8542 10736
rect 10962 10724 10968 10736
rect 8536 10696 10968 10724
rect 8536 10684 8542 10696
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7616 10628 7849 10656
rect 7616 10616 7622 10628
rect 7837 10625 7849 10628
rect 7883 10656 7895 10659
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 7883 10628 8769 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 8757 10625 8769 10628
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 12176 10656 12204 10752
rect 12342 10684 12348 10736
rect 12400 10724 12406 10736
rect 13814 10724 13820 10736
rect 12400 10696 13820 10724
rect 12400 10684 12406 10696
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 15378 10724 15384 10736
rect 14792 10696 15384 10724
rect 14792 10684 14798 10696
rect 15378 10684 15384 10696
rect 15436 10724 15442 10736
rect 15473 10727 15531 10733
rect 15473 10724 15485 10727
rect 15436 10696 15485 10724
rect 15436 10684 15442 10696
rect 15473 10693 15485 10696
rect 15519 10693 15531 10727
rect 15473 10687 15531 10693
rect 9088 10628 12204 10656
rect 13173 10659 13231 10665
rect 9088 10616 9094 10628
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 13538 10656 13544 10668
rect 13219 10628 13544 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 9306 10588 9312 10600
rect 5767 10560 6316 10588
rect 9267 10560 9312 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 10502 10548 10508 10600
rect 10560 10588 10566 10600
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 10560 10560 11069 10588
rect 10560 10548 10566 10560
rect 11057 10557 11069 10560
rect 11103 10588 11115 10591
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11103 10560 11529 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10588 14335 10591
rect 14366 10588 14372 10600
rect 14323 10560 14372 10588
rect 14323 10557 14335 10560
rect 14277 10551 14335 10557
rect 14366 10548 14372 10560
rect 14424 10588 14430 10600
rect 16316 10597 16344 10764
rect 16758 10752 16764 10764
rect 16816 10752 16822 10804
rect 21542 10792 21548 10804
rect 21503 10764 21548 10792
rect 21542 10752 21548 10764
rect 21600 10792 21606 10804
rect 21821 10795 21879 10801
rect 21821 10792 21833 10795
rect 21600 10764 21833 10792
rect 21600 10752 21606 10764
rect 21821 10761 21833 10764
rect 21867 10761 21879 10795
rect 25498 10792 25504 10804
rect 25459 10764 25504 10792
rect 21821 10755 21879 10761
rect 17586 10684 17592 10736
rect 17644 10724 17650 10736
rect 20257 10727 20315 10733
rect 20257 10724 20269 10727
rect 17644 10696 20269 10724
rect 17644 10684 17650 10696
rect 20257 10693 20269 10696
rect 20303 10724 20315 10727
rect 20898 10724 20904 10736
rect 20303 10696 20904 10724
rect 20303 10693 20315 10696
rect 20257 10687 20315 10693
rect 20898 10684 20904 10696
rect 20956 10684 20962 10736
rect 18414 10656 18420 10668
rect 16500 10628 18420 10656
rect 16301 10591 16359 10597
rect 14424 10560 15700 10588
rect 14424 10548 14430 10560
rect 7929 10523 7987 10529
rect 7929 10489 7941 10523
rect 7975 10520 7987 10523
rect 8018 10520 8024 10532
rect 7975 10492 8024 10520
rect 7975 10489 7987 10492
rect 7929 10483 7987 10489
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 9398 10480 9404 10532
rect 9456 10520 9462 10532
rect 9630 10523 9688 10529
rect 9630 10520 9642 10523
rect 9456 10492 9642 10520
rect 9456 10480 9462 10492
rect 9630 10489 9642 10492
rect 9676 10489 9688 10523
rect 12526 10520 12532 10532
rect 12487 10492 12532 10520
rect 9630 10483 9688 10489
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 13541 10523 13599 10529
rect 12676 10492 12721 10520
rect 12676 10480 12682 10492
rect 13541 10489 13553 10523
rect 13587 10520 13599 10523
rect 14598 10523 14656 10529
rect 14598 10520 14610 10523
rect 13587 10492 14610 10520
rect 13587 10489 13599 10492
rect 13541 10483 13599 10489
rect 14200 10464 14228 10492
rect 14598 10489 14610 10492
rect 14644 10489 14656 10523
rect 14598 10483 14656 10489
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4706 10412 4712 10464
rect 4764 10452 4770 10464
rect 4801 10455 4859 10461
rect 4801 10452 4813 10455
rect 4764 10424 4813 10452
rect 4764 10412 4770 10424
rect 4801 10421 4813 10424
rect 4847 10421 4859 10455
rect 4801 10415 4859 10421
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 5169 10455 5227 10461
rect 5169 10452 5181 10455
rect 4948 10424 5181 10452
rect 4948 10412 4954 10424
rect 5169 10421 5181 10424
rect 5215 10421 5227 10455
rect 5169 10415 5227 10421
rect 5905 10455 5963 10461
rect 5905 10421 5917 10455
rect 5951 10452 5963 10455
rect 6086 10452 6092 10464
rect 5951 10424 6092 10452
rect 5951 10421 5963 10424
rect 5905 10415 5963 10421
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 10192 10424 10241 10452
rect 10192 10412 10198 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 14182 10452 14188 10464
rect 14143 10424 14188 10452
rect 10229 10415 10287 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 15194 10452 15200 10464
rect 15155 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15672 10452 15700 10560
rect 16301 10557 16313 10591
rect 16347 10557 16359 10591
rect 16301 10551 16359 10557
rect 16390 10548 16396 10600
rect 16448 10588 16454 10600
rect 16500 10597 16528 10628
rect 18414 10616 18420 10628
rect 18472 10656 18478 10668
rect 18472 10628 18552 10656
rect 18472 10616 18478 10628
rect 16485 10591 16543 10597
rect 16485 10588 16497 10591
rect 16448 10560 16497 10588
rect 16448 10548 16454 10560
rect 16485 10557 16497 10560
rect 16531 10557 16543 10591
rect 17862 10588 17868 10600
rect 17775 10560 17868 10588
rect 16485 10551 16543 10557
rect 17862 10548 17868 10560
rect 17920 10588 17926 10600
rect 18524 10597 18552 10628
rect 20346 10616 20352 10668
rect 20404 10656 20410 10668
rect 21836 10656 21864 10755
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 23382 10684 23388 10736
rect 23440 10724 23446 10736
rect 25590 10724 25596 10736
rect 23440 10696 25596 10724
rect 23440 10684 23446 10696
rect 25590 10684 25596 10696
rect 25648 10684 25654 10736
rect 20404 10628 20944 10656
rect 21836 10628 22508 10656
rect 20404 10616 20410 10628
rect 20916 10597 20944 10628
rect 18325 10591 18383 10597
rect 18325 10588 18337 10591
rect 17920 10560 18337 10588
rect 17920 10548 17926 10560
rect 18325 10557 18337 10560
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 20441 10591 20499 10597
rect 20441 10557 20453 10591
rect 20487 10557 20499 10591
rect 20441 10551 20499 10557
rect 20901 10591 20959 10597
rect 20901 10557 20913 10591
rect 20947 10557 20959 10591
rect 22186 10588 22192 10600
rect 22147 10560 22192 10588
rect 20901 10551 20959 10557
rect 15746 10480 15752 10532
rect 15804 10520 15810 10532
rect 18340 10520 18368 10551
rect 18598 10520 18604 10532
rect 15804 10492 18184 10520
rect 18340 10492 18604 10520
rect 15804 10480 15810 10492
rect 16117 10455 16175 10461
rect 16117 10452 16129 10455
rect 15672 10424 16129 10452
rect 16117 10421 16129 10424
rect 16163 10421 16175 10455
rect 16117 10415 16175 10421
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 18156 10461 18184 10492
rect 18598 10480 18604 10492
rect 18656 10480 18662 10532
rect 19426 10480 19432 10532
rect 19484 10520 19490 10532
rect 19484 10492 19748 10520
rect 19484 10480 19490 10492
rect 17313 10455 17371 10461
rect 17313 10452 17325 10455
rect 17000 10424 17325 10452
rect 17000 10412 17006 10424
rect 17313 10421 17325 10424
rect 17359 10421 17371 10455
rect 17313 10415 17371 10421
rect 18141 10455 18199 10461
rect 18141 10421 18153 10455
rect 18187 10421 18199 10455
rect 18141 10415 18199 10421
rect 18230 10412 18236 10464
rect 18288 10452 18294 10464
rect 19245 10455 19303 10461
rect 19245 10452 19257 10455
rect 18288 10424 19257 10452
rect 18288 10412 18294 10424
rect 19245 10421 19257 10424
rect 19291 10452 19303 10455
rect 19518 10452 19524 10464
rect 19291 10424 19524 10452
rect 19291 10421 19303 10424
rect 19245 10415 19303 10421
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 19720 10461 19748 10492
rect 19705 10455 19763 10461
rect 19705 10421 19717 10455
rect 19751 10452 19763 10455
rect 20456 10452 20484 10551
rect 22186 10548 22192 10560
rect 22244 10548 22250 10600
rect 22480 10597 22508 10628
rect 22830 10616 22836 10668
rect 22888 10656 22894 10668
rect 24029 10659 24087 10665
rect 24029 10656 24041 10659
rect 22888 10628 24041 10656
rect 22888 10616 22894 10628
rect 24029 10625 24041 10628
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 25130 10616 25136 10668
rect 25188 10656 25194 10668
rect 25685 10659 25743 10665
rect 25685 10656 25697 10659
rect 25188 10628 25697 10656
rect 25188 10616 25194 10628
rect 25685 10625 25697 10628
rect 25731 10625 25743 10659
rect 25685 10619 25743 10625
rect 22465 10591 22523 10597
rect 22465 10557 22477 10591
rect 22511 10588 22523 10591
rect 23106 10588 23112 10600
rect 22511 10560 23112 10588
rect 22511 10557 22523 10560
rect 22465 10551 22523 10557
rect 23106 10548 23112 10560
rect 23164 10548 23170 10600
rect 24394 10548 24400 10600
rect 24452 10588 24458 10600
rect 25292 10591 25350 10597
rect 25292 10588 25304 10591
rect 24452 10560 25304 10588
rect 24452 10548 24458 10560
rect 25292 10557 25304 10560
rect 25338 10588 25350 10591
rect 26053 10591 26111 10597
rect 26053 10588 26065 10591
rect 25338 10560 26065 10588
rect 25338 10557 25350 10560
rect 25292 10551 25350 10557
rect 26053 10557 26065 10560
rect 26099 10557 26111 10591
rect 26053 10551 26111 10557
rect 21174 10520 21180 10532
rect 21135 10492 21180 10520
rect 21174 10480 21180 10492
rect 21232 10480 21238 10532
rect 21266 10480 21272 10532
rect 21324 10520 21330 10532
rect 23750 10520 23756 10532
rect 21324 10492 23756 10520
rect 21324 10480 21330 10492
rect 23750 10480 23756 10492
rect 23808 10480 23814 10532
rect 23845 10523 23903 10529
rect 23845 10489 23857 10523
rect 23891 10489 23903 10523
rect 23845 10483 23903 10489
rect 20714 10452 20720 10464
rect 19751 10424 20720 10452
rect 19751 10421 19763 10424
rect 19705 10415 19763 10421
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 22094 10452 22100 10464
rect 22055 10424 22100 10452
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 23014 10452 23020 10464
rect 22975 10424 23020 10452
rect 23014 10412 23020 10424
rect 23072 10452 23078 10464
rect 23385 10455 23443 10461
rect 23385 10452 23397 10455
rect 23072 10424 23397 10452
rect 23072 10412 23078 10424
rect 23385 10421 23397 10424
rect 23431 10452 23443 10455
rect 23474 10452 23480 10464
rect 23431 10424 23480 10452
rect 23431 10421 23443 10424
rect 23385 10415 23443 10421
rect 23474 10412 23480 10424
rect 23532 10452 23538 10464
rect 23860 10452 23888 10483
rect 24946 10452 24952 10464
rect 23532 10424 23888 10452
rect 24907 10424 24952 10452
rect 23532 10412 23538 10424
rect 24946 10412 24952 10424
rect 25004 10412 25010 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 4126 10220 4353 10248
rect 937 10183 995 10189
rect 937 10149 949 10183
rect 983 10180 995 10183
rect 2866 10180 2872 10192
rect 983 10152 2872 10180
rect 983 10149 995 10152
rect 937 10143 995 10149
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 2130 10112 2136 10124
rect 1443 10084 2136 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 2130 10072 2136 10084
rect 2188 10072 2194 10124
rect 2314 10072 2320 10124
rect 2372 10112 2378 10124
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 2372 10084 2421 10112
rect 2372 10072 2378 10084
rect 2409 10081 2421 10084
rect 2455 10081 2467 10115
rect 2682 10112 2688 10124
rect 2643 10084 2688 10112
rect 2409 10075 2467 10081
rect 2682 10072 2688 10084
rect 2740 10112 2746 10124
rect 3421 10115 3479 10121
rect 3421 10112 3433 10115
rect 2740 10084 3433 10112
rect 2740 10072 2746 10084
rect 3421 10081 3433 10084
rect 3467 10112 3479 10115
rect 3786 10112 3792 10124
rect 3467 10084 3792 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 3786 10072 3792 10084
rect 3844 10112 3850 10124
rect 4126 10112 4154 10220
rect 4341 10217 4353 10220
rect 4387 10248 4399 10251
rect 4614 10248 4620 10260
rect 4387 10220 4620 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 8018 10248 8024 10260
rect 7883 10220 8024 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 11241 10251 11299 10257
rect 11241 10248 11253 10251
rect 11112 10220 11253 10248
rect 11112 10208 11118 10220
rect 11241 10217 11253 10220
rect 11287 10217 11299 10251
rect 11241 10211 11299 10217
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12618 10248 12624 10260
rect 12575 10220 12624 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12897 10251 12955 10257
rect 12897 10217 12909 10251
rect 12943 10248 12955 10251
rect 13262 10248 13268 10260
rect 12943 10220 13268 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 15194 10208 15200 10260
rect 15252 10248 15258 10260
rect 15654 10248 15660 10260
rect 15252 10220 15660 10248
rect 15252 10208 15258 10220
rect 15654 10208 15660 10220
rect 15712 10248 15718 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 15712 10220 16313 10248
rect 15712 10208 15718 10220
rect 16301 10217 16313 10220
rect 16347 10217 16359 10251
rect 16301 10211 16359 10217
rect 17221 10251 17279 10257
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 17310 10248 17316 10260
rect 17267 10220 17316 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18414 10248 18420 10260
rect 18375 10220 18420 10248
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 18969 10251 19027 10257
rect 18969 10248 18981 10251
rect 18656 10220 18981 10248
rect 18656 10208 18662 10220
rect 18969 10217 18981 10220
rect 19015 10217 19027 10251
rect 18969 10211 19027 10217
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 21729 10251 21787 10257
rect 21729 10248 21741 10251
rect 21232 10220 21741 10248
rect 21232 10208 21238 10220
rect 21729 10217 21741 10220
rect 21775 10248 21787 10251
rect 21818 10248 21824 10260
rect 21775 10220 21824 10248
rect 21775 10217 21787 10220
rect 21729 10211 21787 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 22278 10248 22284 10260
rect 22239 10220 22284 10248
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 22833 10251 22891 10257
rect 22833 10217 22845 10251
rect 22879 10248 22891 10251
rect 22879 10220 23888 10248
rect 22879 10217 22891 10220
rect 22833 10211 22891 10217
rect 23860 10192 23888 10220
rect 5537 10183 5595 10189
rect 4816 10152 5212 10180
rect 3844 10084 4154 10112
rect 3844 10072 3850 10084
rect 4706 10072 4712 10124
rect 4764 10112 4770 10124
rect 4816 10121 4844 10152
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 4764 10084 4813 10112
rect 4764 10072 4770 10084
rect 4801 10081 4813 10084
rect 4847 10081 4859 10115
rect 5074 10112 5080 10124
rect 5035 10084 5080 10112
rect 4801 10075 4859 10081
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 5184 10112 5212 10152
rect 5537 10149 5549 10183
rect 5583 10180 5595 10183
rect 8662 10180 8668 10192
rect 5583 10152 8668 10180
rect 5583 10149 5595 10152
rect 5537 10143 5595 10149
rect 8662 10140 8668 10152
rect 8720 10140 8726 10192
rect 8757 10183 8815 10189
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 9306 10180 9312 10192
rect 8803 10152 9312 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 10134 10140 10140 10192
rect 10192 10180 10198 10192
rect 10413 10183 10471 10189
rect 10413 10180 10425 10183
rect 10192 10152 10425 10180
rect 10192 10140 10198 10152
rect 10413 10149 10425 10152
rect 10459 10149 10471 10183
rect 10413 10143 10471 10149
rect 10686 10140 10692 10192
rect 10744 10180 10750 10192
rect 10965 10183 11023 10189
rect 10965 10180 10977 10183
rect 10744 10152 10977 10180
rect 10744 10140 10750 10152
rect 10965 10149 10977 10152
rect 11011 10149 11023 10183
rect 13170 10180 13176 10192
rect 13131 10152 13176 10180
rect 10965 10143 11023 10149
rect 13170 10140 13176 10152
rect 13228 10140 13234 10192
rect 15105 10183 15163 10189
rect 15105 10149 15117 10183
rect 15151 10180 15163 10183
rect 15562 10180 15568 10192
rect 15151 10152 15568 10180
rect 15151 10149 15163 10152
rect 15105 10143 15163 10149
rect 15562 10140 15568 10152
rect 15620 10140 15626 10192
rect 17494 10180 17500 10192
rect 17455 10152 17500 10180
rect 17494 10140 17500 10152
rect 17552 10140 17558 10192
rect 19334 10180 19340 10192
rect 19168 10152 19340 10180
rect 6362 10112 6368 10124
rect 5184 10084 6368 10112
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 6546 10072 6552 10124
rect 6604 10112 6610 10124
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 6604 10084 6653 10112
rect 6604 10072 6610 10084
rect 6641 10081 6653 10084
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 8018 10112 8024 10124
rect 7248 10084 8024 10112
rect 7248 10072 7254 10084
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8481 10115 8539 10121
rect 8481 10112 8493 10115
rect 8444 10084 8493 10112
rect 8444 10072 8450 10084
rect 8481 10081 8493 10084
rect 8527 10081 8539 10115
rect 11974 10112 11980 10124
rect 11935 10084 11980 10112
rect 8481 10075 8539 10081
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10081 15347 10115
rect 15289 10075 15347 10081
rect 1946 10004 1952 10056
rect 2004 10044 2010 10056
rect 2869 10047 2927 10053
rect 2869 10044 2881 10047
rect 2004 10016 2881 10044
rect 2004 10004 2010 10016
rect 2869 10013 2881 10016
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4120 10016 5212 10044
rect 4120 10004 4154 10016
rect 2501 9979 2559 9985
rect 2501 9945 2513 9979
rect 2547 9945 2559 9979
rect 2501 9939 2559 9945
rect 1394 9868 1400 9920
rect 1452 9908 1458 9920
rect 1581 9911 1639 9917
rect 1581 9908 1593 9911
rect 1452 9880 1593 9908
rect 1452 9868 1458 9880
rect 1581 9877 1593 9880
rect 1627 9877 1639 9911
rect 1581 9871 1639 9877
rect 1670 9868 1676 9920
rect 1728 9908 1734 9920
rect 1857 9911 1915 9917
rect 1857 9908 1869 9911
rect 1728 9880 1869 9908
rect 1728 9868 1734 9880
rect 1857 9877 1869 9880
rect 1903 9877 1915 9911
rect 1857 9871 1915 9877
rect 2317 9911 2375 9917
rect 2317 9877 2329 9911
rect 2363 9908 2375 9911
rect 2406 9908 2412 9920
rect 2363 9880 2412 9908
rect 2363 9877 2375 9880
rect 2317 9871 2375 9877
rect 2406 9868 2412 9880
rect 2464 9868 2470 9920
rect 2516 9908 2544 9939
rect 3142 9908 3148 9920
rect 2516 9880 3148 9908
rect 3142 9868 3148 9880
rect 3200 9908 3206 9920
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3200 9880 3801 9908
rect 3200 9868 3206 9880
rect 3789 9877 3801 9880
rect 3835 9908 3847 9911
rect 4126 9908 4154 10004
rect 4709 9979 4767 9985
rect 4709 9945 4721 9979
rect 4755 9976 4767 9979
rect 4890 9976 4896 9988
rect 4755 9948 4896 9976
rect 4755 9945 4767 9948
rect 4709 9939 4767 9945
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 5184 9976 5212 10016
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 6052 10016 7113 10044
rect 6052 10004 6058 10016
rect 7101 10013 7113 10016
rect 7147 10044 7159 10047
rect 9030 10044 9036 10056
rect 7147 10016 9036 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 13446 10044 13452 10056
rect 13127 10016 13452 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 6273 9979 6331 9985
rect 6273 9976 6285 9979
rect 5184 9948 6285 9976
rect 6273 9945 6285 9948
rect 6319 9976 6331 9979
rect 6457 9979 6515 9985
rect 6457 9976 6469 9979
rect 6319 9948 6469 9976
rect 6319 9945 6331 9948
rect 6273 9939 6331 9945
rect 6457 9945 6469 9948
rect 6503 9945 6515 9979
rect 6457 9939 6515 9945
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 10336 9976 10364 10007
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 15304 10044 15332 10075
rect 15378 10072 15384 10124
rect 15436 10112 15442 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15436 10084 15761 10112
rect 15436 10072 15442 10084
rect 15749 10081 15761 10084
rect 15795 10112 15807 10115
rect 16206 10112 16212 10124
rect 15795 10084 16212 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 19168 10121 19196 10152
rect 19334 10140 19340 10152
rect 19392 10180 19398 10192
rect 21039 10183 21097 10189
rect 19392 10152 20944 10180
rect 19392 10140 19398 10152
rect 19153 10115 19211 10121
rect 19153 10081 19165 10115
rect 19199 10081 19211 10115
rect 19153 10075 19211 10081
rect 19429 10115 19487 10121
rect 19429 10081 19441 10115
rect 19475 10112 19487 10115
rect 19978 10112 19984 10124
rect 19475 10084 19984 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19978 10072 19984 10084
rect 20036 10112 20042 10124
rect 20346 10112 20352 10124
rect 20036 10084 20352 10112
rect 20036 10072 20042 10084
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 20806 10112 20812 10124
rect 20767 10084 20812 10112
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 20916 10112 20944 10152
rect 21039 10149 21051 10183
rect 21085 10180 21097 10183
rect 21266 10180 21272 10192
rect 21085 10152 21272 10180
rect 21085 10149 21097 10152
rect 21039 10143 21097 10149
rect 21266 10140 21272 10152
rect 21324 10140 21330 10192
rect 23385 10183 23443 10189
rect 23385 10149 23397 10183
rect 23431 10180 23443 10183
rect 23566 10180 23572 10192
rect 23431 10152 23572 10180
rect 23431 10149 23443 10152
rect 23385 10143 23443 10149
rect 23566 10140 23572 10152
rect 23624 10140 23630 10192
rect 23842 10180 23848 10192
rect 23803 10152 23848 10180
rect 23842 10140 23848 10152
rect 23900 10140 23906 10192
rect 24394 10180 24400 10192
rect 24355 10152 24400 10180
rect 24394 10140 24400 10152
rect 24452 10140 24458 10192
rect 22738 10112 22744 10124
rect 20916 10084 22744 10112
rect 21284 10056 21312 10084
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 24854 10072 24860 10124
rect 24912 10112 24918 10124
rect 25225 10115 25283 10121
rect 25225 10112 25237 10115
rect 24912 10084 25237 10112
rect 24912 10072 24918 10084
rect 25225 10081 25237 10084
rect 25271 10112 25283 10115
rect 26050 10112 26056 10124
rect 25271 10084 26056 10112
rect 25271 10081 25283 10084
rect 25225 10075 25283 10081
rect 26050 10072 26056 10084
rect 26108 10072 26114 10124
rect 15838 10044 15844 10056
rect 13596 10016 13641 10044
rect 15304 10016 15516 10044
rect 15799 10016 15844 10044
rect 13596 10004 13602 10016
rect 10686 9976 10692 9988
rect 7064 9948 10692 9976
rect 7064 9936 7070 9948
rect 10686 9936 10692 9948
rect 10744 9936 10750 9988
rect 12115 9979 12173 9985
rect 12115 9945 12127 9979
rect 12161 9976 12173 9979
rect 15488 9976 15516 10016
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10044 17463 10047
rect 17678 10044 17684 10056
rect 17451 10016 17684 10044
rect 17451 10013 17463 10016
rect 17405 10007 17463 10013
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 18966 10004 18972 10056
rect 19024 10044 19030 10056
rect 20438 10044 20444 10056
rect 19024 10016 20444 10044
rect 19024 10004 19030 10016
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 21266 10004 21272 10056
rect 21324 10004 21330 10056
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10044 21971 10047
rect 22094 10044 22100 10056
rect 21959 10016 22100 10044
rect 21959 10013 21971 10016
rect 21913 10007 21971 10013
rect 22094 10004 22100 10016
rect 22152 10004 22158 10056
rect 23106 10004 23112 10056
rect 23164 10044 23170 10056
rect 23753 10047 23811 10053
rect 23753 10044 23765 10047
rect 23164 10016 23765 10044
rect 23164 10004 23170 10016
rect 23753 10013 23765 10016
rect 23799 10044 23811 10047
rect 23934 10044 23940 10056
rect 23799 10016 23940 10044
rect 23799 10013 23811 10016
rect 23753 10007 23811 10013
rect 23934 10004 23940 10016
rect 23992 10004 23998 10056
rect 15930 9976 15936 9988
rect 12161 9948 13584 9976
rect 15488 9948 15936 9976
rect 12161 9945 12173 9948
rect 12115 9939 12173 9945
rect 3835 9880 4154 9908
rect 13556 9908 13584 9948
rect 15930 9936 15936 9948
rect 15988 9936 15994 9988
rect 16850 9936 16856 9988
rect 16908 9976 16914 9988
rect 17957 9979 18015 9985
rect 17957 9976 17969 9979
rect 16908 9948 17969 9976
rect 16908 9936 16914 9948
rect 17957 9945 17969 9948
rect 18003 9976 18015 9979
rect 19518 9976 19524 9988
rect 18003 9948 19524 9976
rect 18003 9945 18015 9948
rect 17957 9939 18015 9945
rect 19518 9936 19524 9948
rect 19576 9936 19582 9988
rect 14550 9908 14556 9920
rect 13556 9880 14556 9908
rect 3835 9877 3847 9880
rect 3789 9871 3847 9877
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 16114 9868 16120 9920
rect 16172 9908 16178 9920
rect 16669 9911 16727 9917
rect 16669 9908 16681 9911
rect 16172 9880 16681 9908
rect 16172 9868 16178 9880
rect 16669 9877 16681 9880
rect 16715 9877 16727 9911
rect 16669 9871 16727 9877
rect 19242 9868 19248 9920
rect 19300 9908 19306 9920
rect 19889 9911 19947 9917
rect 19889 9908 19901 9911
rect 19300 9880 19901 9908
rect 19300 9868 19306 9880
rect 19889 9877 19901 9880
rect 19935 9877 19947 9911
rect 19889 9871 19947 9877
rect 20533 9911 20591 9917
rect 20533 9877 20545 9911
rect 20579 9908 20591 9911
rect 20714 9908 20720 9920
rect 20579 9880 20720 9908
rect 20579 9877 20591 9880
rect 20533 9871 20591 9877
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 25409 9911 25467 9917
rect 25409 9877 25421 9911
rect 25455 9908 25467 9911
rect 27522 9908 27528 9920
rect 25455 9880 27528 9908
rect 25455 9877 25467 9880
rect 25409 9871 25467 9877
rect 27522 9868 27528 9880
rect 27580 9868 27586 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 937 9707 995 9713
rect 937 9673 949 9707
rect 983 9704 995 9707
rect 1857 9707 1915 9713
rect 1857 9704 1869 9707
rect 983 9676 1869 9704
rect 983 9673 995 9676
rect 937 9667 995 9673
rect 1857 9673 1869 9676
rect 1903 9673 1915 9707
rect 1857 9667 1915 9673
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 2685 9707 2743 9713
rect 2280 9676 2325 9704
rect 2280 9664 2286 9676
rect 2685 9673 2697 9707
rect 2731 9704 2743 9707
rect 2866 9704 2872 9716
rect 2731 9676 2872 9704
rect 2731 9673 2743 9676
rect 2685 9667 2743 9673
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 4706 9704 4712 9716
rect 4667 9676 4712 9704
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 6362 9704 6368 9716
rect 6323 9676 6368 9704
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 8018 9704 8024 9716
rect 7979 9676 8024 9704
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 8386 9704 8392 9716
rect 8347 9676 8392 9704
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 10045 9707 10103 9713
rect 10045 9704 10057 9707
rect 9723 9676 10057 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 10045 9673 10057 9676
rect 10091 9704 10103 9707
rect 10134 9704 10140 9716
rect 10091 9676 10140 9704
rect 10091 9673 10103 9676
rect 10045 9667 10103 9673
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 12897 9707 12955 9713
rect 10704 9676 11468 9704
rect 1670 9596 1676 9648
rect 1728 9596 1734 9648
rect 2130 9596 2136 9648
rect 2188 9636 2194 9648
rect 10704 9636 10732 9676
rect 2188 9608 5580 9636
rect 2188 9596 2194 9608
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 1688 9568 1716 9596
rect 5552 9580 5580 9608
rect 9508 9608 10732 9636
rect 10781 9639 10839 9645
rect 9508 9580 9536 9608
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 10962 9636 10968 9648
rect 10827 9608 10968 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 1949 9571 2007 9577
rect 1949 9568 1961 9571
rect 1360 9540 1961 9568
rect 1360 9528 1366 9540
rect 1949 9537 1961 9540
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2314 9528 2320 9580
rect 2372 9568 2378 9580
rect 4890 9568 4896 9580
rect 2372 9540 4154 9568
rect 4803 9540 4896 9568
rect 2372 9528 2378 9540
rect 1728 9503 1786 9509
rect 1728 9469 1740 9503
rect 1774 9500 1786 9503
rect 2498 9500 2504 9512
rect 1774 9472 2504 9500
rect 1774 9469 1786 9472
rect 1728 9463 1786 9469
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9469 3663 9503
rect 4126 9500 4154 9540
rect 4890 9528 4896 9540
rect 4948 9568 4954 9580
rect 5258 9568 5264 9580
rect 4948 9540 5264 9568
rect 4948 9528 4954 9540
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 9490 9568 9496 9580
rect 8711 9540 9496 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 10226 9568 10232 9580
rect 10187 9540 10232 9568
rect 10226 9528 10232 9540
rect 10284 9568 10290 9580
rect 11149 9571 11207 9577
rect 11149 9568 11161 9571
rect 10284 9540 11161 9568
rect 10284 9528 10290 9540
rect 11149 9537 11161 9540
rect 11195 9537 11207 9571
rect 11440 9568 11468 9676
rect 12897 9673 12909 9707
rect 12943 9704 12955 9707
rect 13170 9704 13176 9716
rect 12943 9676 13176 9704
rect 12943 9673 12955 9676
rect 12897 9667 12955 9673
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 15197 9707 15255 9713
rect 15197 9673 15209 9707
rect 15243 9704 15255 9707
rect 17221 9707 17279 9713
rect 17221 9704 17233 9707
rect 15243 9676 17233 9704
rect 15243 9673 15255 9676
rect 15197 9667 15255 9673
rect 17221 9673 17233 9676
rect 17267 9673 17279 9707
rect 17221 9667 17279 9673
rect 17405 9707 17463 9713
rect 17405 9673 17417 9707
rect 17451 9704 17463 9707
rect 17494 9704 17500 9716
rect 17451 9676 17500 9704
rect 17451 9673 17463 9676
rect 17405 9667 17463 9673
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 18230 9704 18236 9716
rect 18191 9676 18236 9704
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 18690 9664 18696 9716
rect 18748 9704 18754 9716
rect 18969 9707 19027 9713
rect 18969 9704 18981 9707
rect 18748 9676 18981 9704
rect 18748 9664 18754 9676
rect 18969 9673 18981 9676
rect 19015 9704 19027 9707
rect 19334 9704 19340 9716
rect 19015 9676 19340 9704
rect 19015 9673 19027 9676
rect 18969 9667 19027 9673
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 20806 9704 20812 9716
rect 20220 9676 20812 9704
rect 20220 9664 20226 9676
rect 20806 9664 20812 9676
rect 20864 9704 20870 9716
rect 21177 9707 21235 9713
rect 21177 9704 21189 9707
rect 20864 9676 21189 9704
rect 20864 9664 20870 9676
rect 21177 9673 21189 9676
rect 21223 9673 21235 9707
rect 21177 9667 21235 9673
rect 22741 9707 22799 9713
rect 22741 9673 22753 9707
rect 22787 9704 22799 9707
rect 23014 9704 23020 9716
rect 22787 9676 23020 9704
rect 22787 9673 22799 9676
rect 22741 9667 22799 9673
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 23842 9664 23848 9716
rect 23900 9704 23906 9716
rect 24673 9707 24731 9713
rect 24673 9704 24685 9707
rect 23900 9676 24685 9704
rect 23900 9664 23906 9676
rect 24673 9673 24685 9676
rect 24719 9673 24731 9707
rect 24673 9667 24731 9673
rect 24854 9664 24860 9716
rect 24912 9704 24918 9716
rect 25222 9704 25228 9716
rect 24912 9676 25228 9704
rect 24912 9664 24918 9676
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 26050 9704 26056 9716
rect 26011 9676 26056 9704
rect 26050 9664 26056 9676
rect 26108 9664 26114 9716
rect 11974 9636 11980 9648
rect 11935 9608 11980 9636
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 14093 9639 14151 9645
rect 14093 9636 14105 9639
rect 13786 9608 14105 9636
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 11440 9540 13369 9568
rect 11149 9531 11207 9537
rect 13357 9537 13369 9540
rect 13403 9568 13415 9571
rect 13538 9568 13544 9580
rect 13403 9540 13544 9568
rect 13403 9537 13415 9540
rect 13357 9531 13415 9537
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 4798 9500 4804 9512
rect 4126 9472 4804 9500
rect 3605 9463 3663 9469
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 1854 9432 1860 9444
rect 1627 9404 1860 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 1854 9392 1860 9404
rect 1912 9392 1918 9444
rect 2961 9435 3019 9441
rect 2961 9432 2973 9435
rect 2424 9404 2973 9432
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1670 9364 1676 9376
rect 1544 9336 1676 9364
rect 1544 9324 1550 9336
rect 1670 9324 1676 9336
rect 1728 9364 1734 9376
rect 2424 9364 2452 9404
rect 2961 9401 2973 9404
rect 3007 9432 3019 9435
rect 3160 9432 3188 9463
rect 3007 9404 3188 9432
rect 3007 9401 3019 9404
rect 2961 9395 3019 9401
rect 3620 9376 3648 9463
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 5074 9500 5080 9512
rect 4987 9472 5080 9500
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 6914 9500 6920 9512
rect 6875 9472 6920 9500
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 5092 9432 5120 9460
rect 5997 9435 6055 9441
rect 5997 9432 6009 9435
rect 4448 9404 6009 9432
rect 4448 9376 4476 9404
rect 5997 9401 6009 9404
rect 6043 9432 6055 9435
rect 6546 9432 6552 9444
rect 6043 9404 6552 9432
rect 6043 9401 6055 9404
rect 5997 9395 6055 9401
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 8754 9392 8760 9444
rect 8812 9432 8818 9444
rect 9306 9432 9312 9444
rect 8812 9404 8857 9432
rect 9267 9404 9312 9432
rect 8812 9392 8818 9404
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 10321 9435 10379 9441
rect 10321 9401 10333 9435
rect 10367 9401 10379 9435
rect 13078 9432 13084 9444
rect 13039 9404 13084 9432
rect 10321 9395 10379 9401
rect 3234 9364 3240 9376
rect 1728 9336 2452 9364
rect 3195 9336 3240 9364
rect 1728 9324 1734 9336
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3602 9324 3608 9376
rect 3660 9324 3666 9376
rect 4341 9367 4399 9373
rect 4341 9333 4353 9367
rect 4387 9364 4399 9367
rect 4430 9364 4436 9376
rect 4387 9336 4436 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 7006 9364 7012 9376
rect 6967 9336 7012 9364
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10336 9364 10364 9395
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 13170 9392 13176 9444
rect 13228 9432 13234 9444
rect 13228 9404 13273 9432
rect 13228 9392 13234 9404
rect 10192 9336 10364 9364
rect 10192 9324 10198 9336
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 13786 9364 13814 9608
rect 14093 9605 14105 9608
rect 14139 9636 14151 9639
rect 20346 9636 20352 9648
rect 14139 9608 20352 9636
rect 14139 9605 14151 9608
rect 14093 9599 14151 9605
rect 20346 9596 20352 9608
rect 20404 9596 20410 9648
rect 20898 9596 20904 9648
rect 20956 9636 20962 9648
rect 23382 9636 23388 9648
rect 20956 9608 23388 9636
rect 20956 9596 20962 9608
rect 23382 9596 23388 9608
rect 23440 9596 23446 9648
rect 25038 9636 25044 9648
rect 23492 9608 25044 9636
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9568 14979 9571
rect 15378 9568 15384 9580
rect 14967 9540 15384 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 19242 9568 19248 9580
rect 19203 9540 19248 9568
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 20254 9568 20260 9580
rect 19484 9540 20260 9568
rect 19484 9528 19490 9540
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 21818 9568 21824 9580
rect 21779 9540 21824 9568
rect 21818 9528 21824 9540
rect 21876 9528 21882 9580
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14884 9472 15025 9500
rect 14884 9460 14890 9472
rect 15013 9469 15025 9472
rect 15059 9500 15071 9503
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15059 9472 15485 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9500 17279 9503
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17267 9472 18061 9500
rect 17267 9469 17279 9472
rect 17221 9463 17279 9469
rect 18049 9469 18061 9472
rect 18095 9500 18107 9503
rect 18506 9500 18512 9512
rect 18095 9472 18512 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 18506 9460 18512 9472
rect 18564 9460 18570 9512
rect 19978 9460 19984 9512
rect 20036 9500 20042 9512
rect 20165 9503 20223 9509
rect 20165 9500 20177 9503
rect 20036 9472 20177 9500
rect 20036 9460 20042 9472
rect 20165 9469 20177 9472
rect 20211 9500 20223 9503
rect 20622 9500 20628 9512
rect 20211 9472 20628 9500
rect 20211 9469 20223 9472
rect 20165 9463 20223 9469
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 20784 9503 20842 9509
rect 20784 9469 20796 9503
rect 20830 9500 20842 9503
rect 21542 9500 21548 9512
rect 20830 9472 21548 9500
rect 20830 9469 20842 9472
rect 20784 9463 20842 9469
rect 21542 9460 21548 9472
rect 21600 9500 21606 9512
rect 23492 9500 23520 9608
rect 25038 9596 25044 9608
rect 25096 9596 25102 9648
rect 24210 9568 24216 9580
rect 24171 9540 24216 9568
rect 24210 9528 24216 9540
rect 24268 9528 24274 9580
rect 21600 9472 23520 9500
rect 25292 9503 25350 9509
rect 21600 9460 21606 9472
rect 25292 9469 25304 9503
rect 25338 9500 25350 9503
rect 25682 9500 25688 9512
rect 25338 9472 25688 9500
rect 25338 9469 25350 9472
rect 25292 9463 25350 9469
rect 25682 9460 25688 9472
rect 25740 9460 25746 9512
rect 15746 9392 15752 9444
rect 15804 9432 15810 9444
rect 16114 9432 16120 9444
rect 15804 9404 16120 9432
rect 15804 9392 15810 9404
rect 16114 9392 16120 9404
rect 16172 9392 16178 9444
rect 16206 9392 16212 9444
rect 16264 9432 16270 9444
rect 16761 9435 16819 9441
rect 16264 9404 16309 9432
rect 16264 9392 16270 9404
rect 16761 9401 16773 9435
rect 16807 9432 16819 9435
rect 17310 9432 17316 9444
rect 16807 9404 17316 9432
rect 16807 9401 16819 9404
rect 16761 9395 16819 9401
rect 17310 9392 17316 9404
rect 17368 9432 17374 9444
rect 17368 9404 19288 9432
rect 17368 9392 17374 9404
rect 15930 9364 15936 9376
rect 13504 9336 13814 9364
rect 15891 9336 15936 9364
rect 13504 9324 13510 9336
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 17678 9364 17684 9376
rect 17639 9336 17684 9364
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 19260 9364 19288 9404
rect 19334 9392 19340 9444
rect 19392 9432 19398 9444
rect 19889 9435 19947 9441
rect 19392 9404 19437 9432
rect 19392 9392 19398 9404
rect 19889 9401 19901 9435
rect 19935 9432 19947 9435
rect 22002 9432 22008 9444
rect 19935 9404 22008 9432
rect 19935 9401 19947 9404
rect 19889 9395 19947 9401
rect 19904 9364 19932 9395
rect 22002 9392 22008 9404
rect 22060 9392 22066 9444
rect 22142 9435 22200 9441
rect 22142 9401 22154 9435
rect 22188 9401 22200 9435
rect 22142 9395 22200 9401
rect 19260 9336 19932 9364
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 20855 9367 20913 9373
rect 20855 9364 20867 9367
rect 20312 9336 20867 9364
rect 20312 9324 20318 9336
rect 20855 9333 20867 9336
rect 20901 9333 20913 9367
rect 20855 9327 20913 9333
rect 21818 9324 21824 9376
rect 21876 9364 21882 9376
rect 22157 9364 22185 9395
rect 22830 9392 22836 9444
rect 22888 9432 22894 9444
rect 23753 9435 23811 9441
rect 23753 9432 23765 9435
rect 22888 9404 23765 9432
rect 22888 9392 22894 9404
rect 23753 9401 23765 9404
rect 23799 9401 23811 9435
rect 23753 9395 23811 9401
rect 23845 9435 23903 9441
rect 23845 9401 23857 9435
rect 23891 9401 23903 9435
rect 25041 9435 25099 9441
rect 25041 9432 25053 9435
rect 23845 9395 23903 9401
rect 24555 9404 25053 9432
rect 22278 9364 22284 9376
rect 21876 9336 22284 9364
rect 21876 9324 21882 9336
rect 22278 9324 22284 9336
rect 22336 9364 22342 9376
rect 23017 9367 23075 9373
rect 23017 9364 23029 9367
rect 22336 9336 23029 9364
rect 22336 9324 22342 9336
rect 23017 9333 23029 9336
rect 23063 9364 23075 9367
rect 23385 9367 23443 9373
rect 23385 9364 23397 9367
rect 23063 9336 23397 9364
rect 23063 9333 23075 9336
rect 23017 9327 23075 9333
rect 23385 9333 23397 9336
rect 23431 9333 23443 9367
rect 23385 9327 23443 9333
rect 23566 9324 23572 9376
rect 23624 9364 23630 9376
rect 23860 9364 23888 9395
rect 24555 9364 24583 9404
rect 25041 9401 25053 9404
rect 25087 9401 25099 9435
rect 25041 9395 25099 9401
rect 23624 9336 24583 9364
rect 23624 9324 23630 9336
rect 24670 9324 24676 9376
rect 24728 9364 24734 9376
rect 25363 9367 25421 9373
rect 25363 9364 25375 9367
rect 24728 9336 25375 9364
rect 24728 9324 24734 9336
rect 25363 9333 25375 9336
rect 25409 9333 25421 9367
rect 25363 9327 25421 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 1670 9160 1676 9172
rect 1627 9132 1676 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 2225 9163 2283 9169
rect 2225 9160 2237 9163
rect 2188 9132 2237 9160
rect 2188 9120 2194 9132
rect 2225 9129 2237 9132
rect 2271 9129 2283 9163
rect 2225 9123 2283 9129
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 3602 9160 3608 9172
rect 3559 9132 3608 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 3786 9160 3792 9172
rect 3747 9132 3792 9160
rect 3786 9120 3792 9132
rect 3844 9160 3850 9172
rect 3844 9132 4108 9160
rect 3844 9120 3850 9132
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1964 9024 1992 9120
rect 3620 9092 3648 9120
rect 3970 9092 3976 9104
rect 3620 9064 3976 9092
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 4080 9101 4108 9132
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 4856 9132 5825 9160
rect 4856 9120 4862 9132
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 7926 9160 7932 9172
rect 7887 9132 7932 9160
rect 5813 9123 5871 9129
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 10686 9160 10692 9172
rect 10647 9132 10692 9160
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 12437 9163 12495 9169
rect 12437 9160 12449 9163
rect 12400 9132 12449 9160
rect 12400 9120 12406 9132
rect 12437 9129 12449 9132
rect 12483 9129 12495 9163
rect 12437 9123 12495 9129
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 13136 9132 13553 9160
rect 13136 9120 13142 9132
rect 13541 9129 13553 9132
rect 13587 9160 13599 9163
rect 13633 9163 13691 9169
rect 13633 9160 13645 9163
rect 13587 9132 13645 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13633 9129 13645 9132
rect 13679 9129 13691 9163
rect 13633 9123 13691 9129
rect 16022 9120 16028 9172
rect 16080 9160 16086 9172
rect 16482 9160 16488 9172
rect 16080 9132 16488 9160
rect 16080 9120 16086 9132
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 21545 9163 21603 9169
rect 21545 9129 21557 9163
rect 21591 9160 21603 9163
rect 22094 9160 22100 9172
rect 21591 9132 22100 9160
rect 21591 9129 21603 9132
rect 21545 9123 21603 9129
rect 22094 9120 22100 9132
rect 22152 9160 22158 9172
rect 22557 9163 22615 9169
rect 22152 9132 22318 9160
rect 22152 9120 22158 9132
rect 4065 9095 4123 9101
rect 4065 9061 4077 9095
rect 4111 9061 4123 9095
rect 4065 9055 4123 9061
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 9861 9095 9919 9101
rect 4212 9064 6592 9092
rect 4212 9052 4218 9064
rect 6564 9036 6592 9064
rect 9861 9061 9873 9095
rect 9907 9092 9919 9095
rect 10042 9092 10048 9104
rect 9907 9064 10048 9092
rect 9907 9061 9919 9064
rect 9861 9055 9919 9061
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 15565 9095 15623 9101
rect 15565 9061 15577 9095
rect 15611 9092 15623 9095
rect 16206 9092 16212 9104
rect 15611 9064 16212 9092
rect 15611 9061 15623 9064
rect 15565 9055 15623 9061
rect 16206 9052 16212 9064
rect 16264 9052 16270 9104
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 17129 9095 17187 9101
rect 17129 9092 17141 9095
rect 17092 9064 17141 9092
rect 17092 9052 17098 9064
rect 17129 9061 17141 9064
rect 17175 9092 17187 9095
rect 17494 9092 17500 9104
rect 17175 9064 17500 9092
rect 17175 9061 17187 9064
rect 17129 9055 17187 9061
rect 17494 9052 17500 9064
rect 17552 9052 17558 9104
rect 18782 9052 18788 9104
rect 18840 9092 18846 9104
rect 18922 9095 18980 9101
rect 18922 9092 18934 9095
rect 18840 9064 18934 9092
rect 18840 9052 18846 9064
rect 18922 9061 18934 9064
rect 18968 9061 18980 9095
rect 18922 9055 18980 9061
rect 21818 9052 21824 9104
rect 21876 9092 21882 9104
rect 21958 9095 22016 9101
rect 21958 9092 21970 9095
rect 21876 9064 21970 9092
rect 21876 9052 21882 9064
rect 21958 9061 21970 9064
rect 22004 9061 22016 9095
rect 22290 9092 22318 9132
rect 22557 9129 22569 9163
rect 22603 9160 22615 9163
rect 23566 9160 23572 9172
rect 22603 9132 23572 9160
rect 22603 9129 22615 9132
rect 22557 9123 22615 9129
rect 23566 9120 23572 9132
rect 23624 9120 23630 9172
rect 23661 9163 23719 9169
rect 23661 9129 23673 9163
rect 23707 9129 23719 9163
rect 23661 9123 23719 9129
rect 23676 9092 23704 9123
rect 24026 9120 24032 9172
rect 24084 9160 24090 9172
rect 24397 9163 24455 9169
rect 24397 9160 24409 9163
rect 24084 9132 24409 9160
rect 24084 9120 24090 9132
rect 24397 9129 24409 9132
rect 24443 9129 24455 9163
rect 24397 9123 24455 9129
rect 22290 9064 23704 9092
rect 21958 9055 22016 9061
rect 2682 9024 2688 9036
rect 1443 8996 1992 9024
rect 2643 8996 2688 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2682 8984 2688 8996
rect 2740 9024 2746 9036
rect 4430 9024 4436 9036
rect 2740 8996 4154 9024
rect 4391 8996 4436 9024
rect 2740 8984 2746 8996
rect 2406 8956 2412 8968
rect 2367 8928 2412 8956
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 4126 8956 4154 8996
rect 4430 8984 4436 8996
rect 4488 9024 4494 9036
rect 5077 9027 5135 9033
rect 5077 9024 5089 9027
rect 4488 8996 5089 9024
rect 4488 8984 4494 8996
rect 5077 8993 5089 8996
rect 5123 8993 5135 9027
rect 6086 9024 6092 9036
rect 6047 8996 6092 9024
rect 5077 8987 5135 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6546 9024 6552 9036
rect 6459 8996 6552 9024
rect 6546 8984 6552 8996
rect 6604 9024 6610 9036
rect 7466 9024 7472 9036
rect 6604 8996 7472 9024
rect 6604 8984 6610 8996
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 13906 9024 13912 9036
rect 13412 8996 13912 9024
rect 13412 8984 13418 8996
rect 13906 8984 13912 8996
rect 13964 9024 13970 9036
rect 14220 9027 14278 9033
rect 14220 9024 14232 9027
rect 13964 8996 14232 9024
rect 13964 8984 13970 8996
rect 14220 8993 14232 8996
rect 14266 8993 14278 9027
rect 14220 8987 14278 8993
rect 16117 9027 16175 9033
rect 16117 8993 16129 9027
rect 16163 9024 16175 9027
rect 16850 9024 16856 9036
rect 16163 8996 16856 9024
rect 16163 8993 16175 8996
rect 16117 8987 16175 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 18598 9024 18604 9036
rect 18559 8996 18604 9024
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 19518 8984 19524 9036
rect 19576 9024 19582 9036
rect 23106 9024 23112 9036
rect 19576 8996 23112 9024
rect 19576 8984 19582 8996
rect 23106 8984 23112 8996
rect 23164 9024 23170 9036
rect 23201 9027 23259 9033
rect 23201 9024 23213 9027
rect 23164 8996 23213 9024
rect 23164 8984 23170 8996
rect 23201 8993 23213 8996
rect 23247 8993 23259 9027
rect 23382 9024 23388 9036
rect 23343 8996 23388 9024
rect 23201 8987 23259 8993
rect 23382 8984 23388 8996
rect 23440 8984 23446 9036
rect 23842 9024 23848 9036
rect 23803 8996 23848 9024
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 25016 9027 25074 9033
rect 25016 8993 25028 9027
rect 25062 9024 25074 9027
rect 25314 9024 25320 9036
rect 25062 8996 25320 9024
rect 25062 8993 25074 8996
rect 25016 8987 25074 8993
rect 25314 8984 25320 8996
rect 25372 8984 25378 9036
rect 4706 8956 4712 8968
rect 4126 8928 4712 8956
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 6779 8928 7573 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 7561 8925 7573 8928
rect 7607 8956 7619 8959
rect 8846 8956 8852 8968
rect 7607 8928 8852 8956
rect 7607 8925 7619 8928
rect 7561 8919 7619 8925
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 9214 8916 9220 8968
rect 9272 8956 9278 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 9272 8928 9781 8956
rect 9272 8916 9278 8928
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 3050 8848 3056 8900
rect 3108 8888 3114 8900
rect 5350 8888 5356 8900
rect 3108 8860 5356 8888
rect 3108 8848 3114 8860
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 8481 8891 8539 8897
rect 8481 8857 8493 8891
rect 8527 8888 8539 8891
rect 9030 8888 9036 8900
rect 8527 8860 9036 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 9030 8848 9036 8860
rect 9088 8848 9094 8900
rect 9398 8848 9404 8900
rect 9456 8888 9462 8900
rect 10060 8888 10088 8919
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 11388 8928 12081 8956
rect 11388 8916 11394 8928
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 15473 8959 15531 8965
rect 15473 8925 15485 8959
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 15948 8928 16528 8956
rect 9456 8860 10088 8888
rect 12989 8891 13047 8897
rect 9456 8848 9462 8860
rect 12989 8857 13001 8891
rect 13035 8888 13047 8891
rect 13170 8888 13176 8900
rect 13035 8860 13176 8888
rect 13035 8857 13047 8860
rect 12989 8851 13047 8857
rect 13170 8848 13176 8860
rect 13228 8888 13234 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 13228 8860 13369 8888
rect 13228 8848 13234 8860
rect 13357 8857 13369 8860
rect 13403 8888 13415 8891
rect 13814 8888 13820 8900
rect 13403 8860 13820 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 14323 8891 14381 8897
rect 14323 8857 14335 8891
rect 14369 8888 14381 8891
rect 15013 8891 15071 8897
rect 15013 8888 15025 8891
rect 14369 8860 15025 8888
rect 14369 8857 14381 8860
rect 14323 8851 14381 8857
rect 15013 8857 15025 8860
rect 15059 8888 15071 8891
rect 15488 8888 15516 8919
rect 15059 8860 15516 8888
rect 15059 8857 15071 8860
rect 15013 8851 15071 8857
rect 5258 8780 5264 8832
rect 5316 8820 5322 8832
rect 5445 8823 5503 8829
rect 5445 8820 5457 8823
rect 5316 8792 5457 8820
rect 5316 8780 5322 8792
rect 5445 8789 5457 8792
rect 5491 8789 5503 8823
rect 5445 8783 5503 8789
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7009 8823 7067 8829
rect 7009 8820 7021 8823
rect 6972 8792 7021 8820
rect 6972 8780 6978 8792
rect 7009 8789 7021 8792
rect 7055 8789 7067 8823
rect 7466 8820 7472 8832
rect 7379 8792 7472 8820
rect 7009 8783 7067 8789
rect 7466 8780 7472 8792
rect 7524 8820 7530 8832
rect 8386 8820 8392 8832
rect 7524 8792 8392 8820
rect 7524 8780 7530 8792
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8754 8820 8760 8832
rect 8715 8792 8760 8820
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9217 8823 9275 8829
rect 9217 8789 9229 8823
rect 9263 8820 9275 8823
rect 9490 8820 9496 8832
rect 9263 8792 9496 8820
rect 9263 8789 9275 8792
rect 9217 8783 9275 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 13541 8823 13599 8829
rect 13541 8789 13553 8823
rect 13587 8820 13599 8823
rect 15948 8820 15976 8928
rect 13587 8792 15976 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 16172 8792 16405 8820
rect 16172 8780 16178 8792
rect 16393 8789 16405 8792
rect 16439 8789 16451 8823
rect 16500 8820 16528 8928
rect 16758 8916 16764 8968
rect 16816 8956 16822 8968
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 16816 8928 17049 8956
rect 16816 8916 16822 8928
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 17310 8956 17316 8968
rect 17271 8928 17316 8956
rect 17037 8919 17095 8925
rect 17310 8916 17316 8928
rect 17368 8916 17374 8968
rect 20438 8916 20444 8968
rect 20496 8956 20502 8968
rect 21358 8956 21364 8968
rect 20496 8928 21364 8956
rect 20496 8916 20502 8928
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 21637 8959 21695 8965
rect 21637 8925 21649 8959
rect 21683 8956 21695 8959
rect 21726 8956 21732 8968
rect 21683 8928 21732 8956
rect 21683 8925 21695 8928
rect 21637 8919 21695 8925
rect 21726 8916 21732 8928
rect 21784 8916 21790 8968
rect 22002 8916 22008 8968
rect 22060 8956 22066 8968
rect 22830 8956 22836 8968
rect 22060 8928 22836 8956
rect 22060 8916 22066 8928
rect 22830 8916 22836 8928
rect 22888 8916 22894 8968
rect 23290 8916 23296 8968
rect 23348 8956 23354 8968
rect 23566 8956 23572 8968
rect 23348 8928 23572 8956
rect 23348 8916 23354 8928
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 23658 8916 23664 8968
rect 23716 8956 23722 8968
rect 24118 8956 24124 8968
rect 23716 8928 24124 8956
rect 23716 8916 23722 8928
rect 24118 8916 24124 8928
rect 24176 8916 24182 8968
rect 16850 8848 16856 8900
rect 16908 8888 16914 8900
rect 17402 8888 17408 8900
rect 16908 8860 17408 8888
rect 16908 8848 16914 8860
rect 17402 8848 17408 8860
rect 17460 8848 17466 8900
rect 25087 8891 25145 8897
rect 25087 8888 25099 8891
rect 18616 8860 25099 8888
rect 18616 8820 18644 8860
rect 25087 8857 25099 8860
rect 25133 8857 25145 8891
rect 25087 8851 25145 8857
rect 16500 8792 18644 8820
rect 16393 8783 16451 8789
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 19521 8823 19579 8829
rect 19521 8820 19533 8823
rect 19392 8792 19533 8820
rect 19392 8780 19398 8792
rect 19521 8789 19533 8792
rect 19567 8820 19579 8823
rect 19797 8823 19855 8829
rect 19797 8820 19809 8823
rect 19567 8792 19809 8820
rect 19567 8789 19579 8792
rect 19521 8783 19579 8789
rect 19797 8789 19809 8792
rect 19843 8789 19855 8823
rect 21174 8820 21180 8832
rect 21135 8792 21180 8820
rect 19797 8783 19855 8789
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4801 8619 4859 8625
rect 4801 8616 4813 8619
rect 4120 8588 4813 8616
rect 4120 8576 4126 8588
rect 4801 8585 4813 8588
rect 4847 8585 4859 8619
rect 6086 8616 6092 8628
rect 6047 8588 6092 8616
rect 4801 8579 4859 8585
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 3234 8480 3240 8492
rect 3191 8452 3240 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 1670 8412 1676 8424
rect 1631 8384 1676 8412
rect 1670 8372 1676 8384
rect 1728 8372 1734 8424
rect 4522 8412 4528 8424
rect 3481 8384 4528 8412
rect 3050 8344 3056 8356
rect 2963 8316 3056 8344
rect 3050 8304 3056 8316
rect 3108 8344 3114 8356
rect 3481 8353 3509 8384
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 4816 8412 4844 8579
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 6457 8619 6515 8625
rect 6457 8585 6469 8619
rect 6503 8616 6515 8619
rect 6546 8616 6552 8628
rect 6503 8588 6552 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 8481 8619 8539 8625
rect 8481 8585 8493 8619
rect 8527 8616 8539 8619
rect 8754 8616 8760 8628
rect 8527 8588 8760 8616
rect 8527 8585 8539 8588
rect 8481 8579 8539 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 8904 8588 8949 8616
rect 8904 8576 8910 8588
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 9125 8619 9183 8625
rect 9125 8616 9137 8619
rect 9088 8588 9137 8616
rect 9088 8576 9094 8588
rect 9125 8585 9137 8588
rect 9171 8585 9183 8619
rect 9125 8579 9183 8585
rect 11471 8619 11529 8625
rect 11471 8585 11483 8619
rect 11517 8616 11529 8619
rect 12986 8616 12992 8628
rect 11517 8588 12992 8616
rect 11517 8585 11529 8588
rect 11471 8579 11529 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 13320 8588 13369 8616
rect 13320 8576 13326 8588
rect 13357 8585 13369 8588
rect 13403 8585 13415 8619
rect 14366 8616 14372 8628
rect 13357 8579 13415 8585
rect 13786 8588 14372 8616
rect 5534 8480 5540 8492
rect 5495 8452 5540 8480
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 7024 8480 7052 8576
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 9306 8548 9312 8560
rect 8260 8520 9312 8548
rect 8260 8508 8266 8520
rect 9306 8508 9312 8520
rect 9364 8548 9370 8560
rect 9953 8551 10011 8557
rect 9953 8548 9965 8551
rect 9364 8520 9965 8548
rect 9364 8508 9370 8520
rect 9953 8517 9965 8520
rect 9999 8517 10011 8551
rect 11790 8548 11796 8560
rect 11751 8520 11796 8548
rect 9953 8511 10011 8517
rect 11790 8508 11796 8520
rect 11848 8508 11854 8560
rect 13078 8508 13084 8560
rect 13136 8548 13142 8560
rect 13786 8548 13814 8588
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 14599 8619 14657 8625
rect 14599 8585 14611 8619
rect 14645 8616 14657 8619
rect 15746 8616 15752 8628
rect 14645 8588 15752 8616
rect 14645 8585 14657 8588
rect 14599 8579 14657 8585
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 17034 8616 17040 8628
rect 16995 8588 17040 8616
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 18279 8619 18337 8625
rect 18279 8585 18291 8619
rect 18325 8616 18337 8619
rect 19242 8616 19248 8628
rect 18325 8588 19248 8616
rect 18325 8585 18337 8588
rect 18279 8579 18337 8585
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 20254 8616 20260 8628
rect 20215 8588 20260 8616
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 20622 8576 20628 8628
rect 20680 8616 20686 8628
rect 22830 8616 22836 8628
rect 20680 8588 22836 8616
rect 20680 8576 20686 8588
rect 22830 8576 22836 8588
rect 22888 8616 22894 8628
rect 23017 8619 23075 8625
rect 23017 8616 23029 8619
rect 22888 8588 23029 8616
rect 22888 8576 22894 8588
rect 23017 8585 23029 8588
rect 23063 8616 23075 8619
rect 23842 8616 23848 8628
rect 23063 8588 23848 8616
rect 23063 8585 23075 8588
rect 23017 8579 23075 8585
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 13136 8520 13814 8548
rect 13136 8508 13142 8520
rect 13906 8508 13912 8560
rect 13964 8548 13970 8560
rect 14277 8551 14335 8557
rect 14277 8548 14289 8551
rect 13964 8520 14289 8548
rect 13964 8508 13970 8520
rect 14277 8517 14289 8520
rect 14323 8548 14335 8551
rect 17865 8551 17923 8557
rect 14323 8520 16849 8548
rect 14323 8517 14335 8520
rect 14277 8511 14335 8517
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7024 8452 7573 8480
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 7561 8443 7619 8449
rect 9232 8452 10701 8480
rect 9232 8424 9260 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 4816 8384 4997 8412
rect 4985 8381 4997 8384
rect 5031 8381 5043 8415
rect 5442 8412 5448 8424
rect 5403 8384 5448 8412
rect 4985 8375 5043 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 9214 8412 9220 8424
rect 7760 8384 9220 8412
rect 3466 8347 3524 8353
rect 3466 8344 3478 8347
rect 3108 8316 3478 8344
rect 3108 8304 3114 8316
rect 3466 8313 3478 8316
rect 3512 8313 3524 8347
rect 3466 8307 3524 8313
rect 3602 8304 3608 8356
rect 3660 8344 3666 8356
rect 7760 8344 7788 8384
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 11400 8415 11458 8421
rect 11400 8381 11412 8415
rect 11446 8412 11458 8415
rect 11808 8412 11836 8508
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 14090 8480 14096 8492
rect 12308 8452 14096 8480
rect 12308 8440 12314 8452
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15160 8452 15485 8480
rect 15160 8440 15166 8452
rect 15473 8449 15485 8452
rect 15519 8480 15531 8483
rect 15838 8480 15844 8492
rect 15519 8452 15844 8480
rect 15519 8449 15531 8452
rect 15473 8443 15531 8449
rect 15838 8440 15844 8452
rect 15896 8440 15902 8492
rect 16821 8480 16849 8520
rect 17865 8517 17877 8551
rect 17911 8548 17923 8551
rect 18598 8548 18604 8560
rect 17911 8520 18604 8548
rect 17911 8517 17923 8520
rect 17865 8511 17923 8517
rect 18598 8508 18604 8520
rect 18656 8508 18662 8560
rect 20073 8551 20131 8557
rect 20073 8548 20085 8551
rect 18892 8520 20085 8548
rect 18892 8480 18920 8520
rect 20073 8517 20085 8520
rect 20119 8517 20131 8551
rect 20073 8511 20131 8517
rect 16821 8452 18920 8480
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8480 19303 8483
rect 20272 8480 20300 8576
rect 20346 8508 20352 8560
rect 20404 8548 20410 8560
rect 25363 8551 25421 8557
rect 25363 8548 25375 8551
rect 20404 8520 25375 8548
rect 20404 8508 20410 8520
rect 25363 8517 25375 8520
rect 25409 8517 25421 8551
rect 25363 8511 25421 8517
rect 19291 8452 20300 8480
rect 19291 8449 19303 8452
rect 19245 8443 19303 8449
rect 21174 8440 21180 8492
rect 21232 8480 21238 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21232 8452 21833 8480
rect 21232 8440 21238 8452
rect 21821 8449 21833 8452
rect 21867 8480 21879 8483
rect 23750 8480 23756 8492
rect 21867 8452 23756 8480
rect 21867 8449 21879 8452
rect 21821 8443 21879 8449
rect 23750 8440 23756 8452
rect 23808 8440 23814 8492
rect 24210 8480 24216 8492
rect 24171 8452 24216 8480
rect 24210 8440 24216 8452
rect 24268 8440 24274 8492
rect 12434 8412 12440 8424
rect 11446 8384 11836 8412
rect 12395 8384 12440 8412
rect 11446 8381 11458 8384
rect 11400 8375 11458 8381
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 14108 8412 14136 8440
rect 14496 8415 14554 8421
rect 14496 8412 14508 8415
rect 14108 8384 14508 8412
rect 14496 8381 14508 8384
rect 14542 8412 14554 8415
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14542 8384 14933 8412
rect 14542 8381 14554 8384
rect 14496 8375 14554 8381
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 18176 8415 18234 8421
rect 18176 8412 18188 8415
rect 14921 8375 14979 8381
rect 15672 8384 18188 8412
rect 9398 8344 9404 8356
rect 3660 8316 7788 8344
rect 9359 8316 9404 8344
rect 3660 8304 3666 8316
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 9493 8347 9551 8353
rect 9493 8313 9505 8347
rect 9539 8313 9551 8347
rect 12799 8347 12857 8353
rect 12799 8344 12811 8347
rect 9493 8307 9551 8313
rect 12544 8316 12811 8344
rect 2041 8279 2099 8285
rect 2041 8245 2053 8279
rect 2087 8276 2099 8279
rect 2130 8276 2136 8288
rect 2087 8248 2136 8276
rect 2087 8245 2099 8248
rect 2041 8239 2099 8245
rect 2130 8236 2136 8248
rect 2188 8236 2194 8288
rect 2682 8276 2688 8288
rect 2643 8248 2688 8276
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 4065 8279 4123 8285
rect 4065 8245 4077 8279
rect 4111 8276 4123 8279
rect 4246 8276 4252 8288
rect 4111 8248 4252 8276
rect 4111 8245 4123 8248
rect 4065 8239 4123 8245
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4430 8276 4436 8288
rect 4391 8248 4436 8276
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 7466 8276 7472 8288
rect 7427 8248 7472 8276
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 7926 8236 7932 8288
rect 7984 8276 7990 8288
rect 7984 8248 8029 8276
rect 7984 8236 7990 8248
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9508 8276 9536 8307
rect 12544 8288 12572 8316
rect 12799 8313 12811 8316
rect 12845 8344 12857 8347
rect 12845 8316 13952 8344
rect 12845 8313 12857 8316
rect 12799 8307 12857 8313
rect 9088 8248 9536 8276
rect 9088 8236 9094 8248
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10321 8279 10379 8285
rect 10321 8276 10333 8279
rect 10192 8248 10333 8276
rect 10192 8236 10198 8248
rect 10321 8245 10333 8248
rect 10367 8245 10379 8279
rect 10321 8239 10379 8245
rect 11241 8279 11299 8285
rect 11241 8245 11253 8279
rect 11287 8276 11299 8279
rect 11330 8276 11336 8288
rect 11287 8248 11336 8276
rect 11287 8245 11299 8248
rect 11241 8239 11299 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 12253 8279 12311 8285
rect 12253 8245 12265 8279
rect 12299 8276 12311 8279
rect 12342 8276 12348 8288
rect 12299 8248 12348 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 12342 8236 12348 8248
rect 12400 8276 12406 8288
rect 12526 8276 12532 8288
rect 12400 8248 12532 8276
rect 12400 8236 12406 8248
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 13722 8276 13728 8288
rect 13683 8248 13728 8276
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 13924 8276 13952 8316
rect 13998 8304 14004 8356
rect 14056 8344 14062 8356
rect 15672 8344 15700 8384
rect 18176 8381 18188 8384
rect 18222 8412 18234 8415
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 18222 8384 18613 8412
rect 18222 8381 18234 8384
rect 18176 8375 18234 8381
rect 18601 8381 18613 8384
rect 18647 8381 18659 8415
rect 18601 8375 18659 8381
rect 20073 8415 20131 8421
rect 20073 8381 20085 8415
rect 20119 8412 20131 8415
rect 20768 8415 20826 8421
rect 20768 8412 20780 8415
rect 20119 8384 20780 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 20768 8381 20780 8384
rect 20814 8412 20826 8415
rect 21269 8415 21327 8421
rect 21269 8412 21281 8415
rect 20814 8384 21281 8412
rect 20814 8381 20826 8384
rect 20768 8375 20826 8381
rect 21269 8381 21281 8384
rect 21315 8381 21327 8415
rect 21269 8375 21327 8381
rect 25038 8372 25044 8424
rect 25096 8412 25102 8424
rect 25292 8415 25350 8421
rect 25292 8412 25304 8415
rect 25096 8384 25304 8412
rect 25096 8372 25102 8384
rect 25292 8381 25304 8384
rect 25338 8412 25350 8415
rect 25338 8384 25820 8412
rect 25338 8381 25350 8384
rect 25292 8375 25350 8381
rect 14056 8316 15700 8344
rect 14056 8304 14062 8316
rect 19334 8304 19340 8356
rect 19392 8344 19398 8356
rect 19392 8316 19437 8344
rect 19392 8304 19398 8316
rect 19518 8304 19524 8356
rect 19576 8344 19582 8356
rect 19889 8347 19947 8353
rect 19889 8344 19901 8347
rect 19576 8316 19901 8344
rect 19576 8304 19582 8316
rect 19889 8313 19901 8316
rect 19935 8313 19947 8347
rect 19889 8307 19947 8313
rect 19978 8304 19984 8356
rect 20036 8344 20042 8356
rect 20855 8347 20913 8353
rect 20855 8344 20867 8347
rect 20036 8316 20867 8344
rect 20036 8304 20042 8316
rect 20855 8313 20867 8316
rect 20901 8313 20913 8347
rect 20855 8307 20913 8313
rect 22142 8347 22200 8353
rect 22142 8313 22154 8347
rect 22188 8313 22200 8347
rect 23382 8344 23388 8356
rect 23343 8316 23388 8344
rect 22142 8307 22200 8313
rect 14182 8276 14188 8288
rect 13924 8248 14188 8276
rect 14182 8236 14188 8248
rect 14240 8276 14246 8288
rect 15381 8279 15439 8285
rect 15381 8276 15393 8279
rect 14240 8248 15393 8276
rect 14240 8236 14246 8248
rect 15381 8245 15393 8248
rect 15427 8276 15439 8279
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15427 8248 15853 8276
rect 15427 8245 15439 8248
rect 15381 8239 15439 8245
rect 15841 8245 15853 8248
rect 15887 8245 15899 8279
rect 15841 8239 15899 8245
rect 16114 8236 16120 8288
rect 16172 8276 16178 8288
rect 16393 8279 16451 8285
rect 16393 8276 16405 8279
rect 16172 8248 16405 8276
rect 16172 8236 16178 8248
rect 16393 8245 16405 8248
rect 16439 8245 16451 8279
rect 16393 8239 16451 8245
rect 16758 8236 16764 8288
rect 16816 8276 16822 8288
rect 17313 8279 17371 8285
rect 17313 8276 17325 8279
rect 16816 8248 17325 8276
rect 16816 8236 16822 8248
rect 17313 8245 17325 8248
rect 17359 8245 17371 8279
rect 17313 8239 17371 8245
rect 18138 8236 18144 8288
rect 18196 8276 18202 8288
rect 18782 8276 18788 8288
rect 18196 8248 18788 8276
rect 18196 8236 18202 8248
rect 18782 8236 18788 8248
rect 18840 8276 18846 8288
rect 18969 8279 19027 8285
rect 18969 8276 18981 8279
rect 18840 8248 18981 8276
rect 18840 8236 18846 8248
rect 18969 8245 18981 8248
rect 19015 8245 19027 8279
rect 18969 8239 19027 8245
rect 21542 8236 21548 8288
rect 21600 8276 21606 8288
rect 21637 8279 21695 8285
rect 21637 8276 21649 8279
rect 21600 8248 21649 8276
rect 21600 8236 21606 8248
rect 21637 8245 21649 8248
rect 21683 8276 21695 8279
rect 21818 8276 21824 8288
rect 21683 8248 21824 8276
rect 21683 8245 21695 8248
rect 21637 8239 21695 8245
rect 21818 8236 21824 8248
rect 21876 8276 21882 8288
rect 22157 8276 22185 8307
rect 23382 8304 23388 8316
rect 23440 8304 23446 8356
rect 23753 8347 23811 8353
rect 23753 8313 23765 8347
rect 23799 8313 23811 8347
rect 23753 8307 23811 8313
rect 22738 8276 22744 8288
rect 21876 8248 22185 8276
rect 22699 8248 22744 8276
rect 21876 8236 21882 8248
rect 22738 8236 22744 8248
rect 22796 8236 22802 8288
rect 23768 8276 23796 8307
rect 23842 8304 23848 8356
rect 23900 8344 23906 8356
rect 23900 8316 23945 8344
rect 23900 8304 23906 8316
rect 25792 8288 25820 8384
rect 24026 8276 24032 8288
rect 23768 8248 24032 8276
rect 24026 8236 24032 8248
rect 24084 8236 24090 8288
rect 25041 8279 25099 8285
rect 25041 8245 25053 8279
rect 25087 8276 25099 8279
rect 25314 8276 25320 8288
rect 25087 8248 25320 8276
rect 25087 8245 25099 8248
rect 25041 8239 25099 8245
rect 25314 8236 25320 8248
rect 25372 8236 25378 8288
rect 25774 8276 25780 8288
rect 25735 8248 25780 8276
rect 25774 8236 25780 8248
rect 25832 8236 25838 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2041 8075 2099 8081
rect 2041 8041 2053 8075
rect 2087 8072 2099 8075
rect 2406 8072 2412 8084
rect 2087 8044 2412 8072
rect 2087 8041 2099 8044
rect 2041 8035 2099 8041
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 3142 8072 3148 8084
rect 3103 8044 3148 8072
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 3292 8044 5825 8072
rect 3292 8032 3298 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 5813 8035 5871 8041
rect 11793 8075 11851 8081
rect 11793 8041 11805 8075
rect 11839 8041 11851 8075
rect 11793 8035 11851 8041
rect 12345 8075 12403 8081
rect 12345 8041 12357 8075
rect 12391 8072 12403 8075
rect 12618 8072 12624 8084
rect 12391 8044 12624 8072
rect 12391 8041 12403 8044
rect 12345 8035 12403 8041
rect 2314 8004 2320 8016
rect 2275 7976 2320 8004
rect 2314 7964 2320 7976
rect 2372 7964 2378 8016
rect 4246 8004 4252 8016
rect 4207 7976 4252 8004
rect 4246 7964 4252 7976
rect 4304 7964 4310 8016
rect 6638 8004 6644 8016
rect 6599 7976 6644 8004
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 7466 7964 7472 8016
rect 7524 8004 7530 8016
rect 7653 8007 7711 8013
rect 7653 8004 7665 8007
rect 7524 7976 7665 8004
rect 7524 7964 7530 7976
rect 7653 7973 7665 7976
rect 7699 8004 7711 8007
rect 7926 8004 7932 8016
rect 7699 7976 7932 8004
rect 7699 7973 7711 7976
rect 7653 7967 7711 7973
rect 7926 7964 7932 7976
rect 7984 8004 7990 8016
rect 10039 8007 10097 8013
rect 10039 8004 10051 8007
rect 7984 7976 10051 8004
rect 7984 7964 7990 7976
rect 10039 7973 10051 7976
rect 10085 8004 10097 8007
rect 10134 8004 10140 8016
rect 10085 7976 10140 8004
rect 10085 7973 10097 7976
rect 10039 7967 10097 7973
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 11808 8004 11836 8035
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 16114 8072 16120 8084
rect 16075 8044 16120 8072
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 17092 8044 17509 8072
rect 17092 8032 17098 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 18417 8075 18475 8081
rect 18417 8072 18429 8075
rect 17497 8035 17555 8041
rect 17880 8044 18429 8072
rect 12526 8004 12532 8016
rect 11808 7976 12532 8004
rect 12526 7964 12532 7976
rect 12584 7964 12590 8016
rect 13262 7964 13268 8016
rect 13320 8004 13326 8016
rect 13817 8007 13875 8013
rect 13817 8004 13829 8007
rect 13320 7976 13829 8004
rect 13320 7964 13326 7976
rect 13817 7973 13829 7976
rect 13863 7973 13875 8007
rect 13817 7967 13875 7973
rect 15703 8007 15761 8013
rect 15703 7973 15715 8007
rect 15749 8004 15761 8007
rect 16758 8004 16764 8016
rect 15749 7976 16764 8004
rect 15749 7973 15761 7976
rect 15703 7967 15761 7973
rect 16758 7964 16764 7976
rect 16816 7964 16822 8016
rect 16942 8013 16948 8016
rect 16939 7967 16948 8013
rect 17000 8004 17006 8016
rect 17310 8004 17316 8016
rect 17000 7976 17316 8004
rect 16942 7964 16948 7967
rect 17000 7964 17006 7976
rect 17310 7964 17316 7976
rect 17368 7964 17374 8016
rect 8297 7939 8355 7945
rect 8297 7905 8309 7939
rect 8343 7905 8355 7939
rect 8478 7936 8484 7948
rect 8439 7908 8484 7936
rect 8297 7899 8355 7905
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 2038 7760 2044 7812
rect 2096 7800 2102 7812
rect 2516 7800 2544 7831
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 3384 7840 4169 7868
rect 3384 7828 3390 7840
rect 4157 7837 4169 7840
rect 4203 7868 4215 7871
rect 4338 7868 4344 7880
rect 4203 7840 4344 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5442 7868 5448 7880
rect 5215 7840 5448 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 4448 7800 4476 7831
rect 5442 7828 5448 7840
rect 5500 7868 5506 7880
rect 6270 7868 6276 7880
rect 5500 7840 6276 7868
rect 5500 7828 5506 7840
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6411 7840 6561 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 6549 7837 6561 7840
rect 6595 7868 6607 7871
rect 6730 7868 6736 7880
rect 6595 7840 6736 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 8202 7868 8208 7880
rect 7024 7840 8208 7868
rect 7024 7800 7052 7840
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8312 7868 8340 7899
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 12434 7936 12440 7948
rect 8803 7908 12440 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 12434 7896 12440 7908
rect 12492 7936 12498 7948
rect 12989 7939 13047 7945
rect 12989 7936 13001 7939
rect 12492 7908 13001 7936
rect 12492 7896 12498 7908
rect 12989 7905 13001 7908
rect 13035 7905 13047 7939
rect 15600 7939 15658 7945
rect 15600 7936 15612 7939
rect 12989 7899 13047 7905
rect 15304 7908 15612 7936
rect 8386 7868 8392 7880
rect 8312 7840 8392 7868
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 9674 7868 9680 7880
rect 9635 7840 9680 7868
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11296 7840 11437 7868
rect 11296 7828 11302 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7868 13599 7871
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13587 7840 13737 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 13725 7837 13737 7840
rect 13771 7868 13783 7871
rect 14734 7868 14740 7880
rect 13771 7840 14740 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 2096 7772 7052 7800
rect 7101 7803 7159 7809
rect 2096 7760 2102 7772
rect 7101 7769 7113 7803
rect 7147 7800 7159 7803
rect 8018 7800 8024 7812
rect 7147 7772 8024 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 9398 7800 9404 7812
rect 9311 7772 9404 7800
rect 9398 7760 9404 7772
rect 9456 7800 9462 7812
rect 13170 7800 13176 7812
rect 9456 7772 13176 7800
rect 9456 7760 9462 7772
rect 13170 7760 13176 7772
rect 13228 7760 13234 7812
rect 14274 7800 14280 7812
rect 14235 7772 14280 7800
rect 14274 7760 14280 7772
rect 14332 7760 14338 7812
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 3786 7732 3792 7744
rect 3651 7704 3792 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 5442 7732 5448 7744
rect 5403 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 10100 7704 10609 7732
rect 10100 7692 10106 7704
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10597 7695 10655 7701
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 12621 7735 12679 7741
rect 12621 7732 12633 7735
rect 12584 7704 12633 7732
rect 12584 7692 12590 7704
rect 12621 7701 12633 7704
rect 12667 7701 12679 7735
rect 12621 7695 12679 7701
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 15304 7732 15332 7908
rect 15600 7905 15612 7908
rect 15646 7936 15658 7939
rect 16206 7936 16212 7948
rect 15646 7908 16212 7936
rect 15646 7905 15658 7908
rect 15600 7899 15658 7905
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 17402 7936 17408 7948
rect 16623 7908 17408 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 17402 7896 17408 7908
rect 17460 7936 17466 7948
rect 17880 7936 17908 8044
rect 18417 8041 18429 8044
rect 18463 8041 18475 8075
rect 19334 8072 19340 8084
rect 19295 8044 19340 8072
rect 18417 8035 18475 8041
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 23477 8075 23535 8081
rect 23477 8072 23489 8075
rect 22664 8044 23489 8072
rect 21818 7964 21824 8016
rect 21876 8004 21882 8016
rect 22142 8007 22200 8013
rect 22142 8004 22154 8007
rect 21876 7976 22154 8004
rect 21876 7964 21882 7976
rect 22142 7973 22154 7976
rect 22188 7973 22200 8007
rect 22142 7967 22200 7973
rect 17460 7908 17908 7936
rect 17460 7896 17466 7908
rect 18230 7896 18236 7948
rect 18288 7936 18294 7948
rect 18325 7939 18383 7945
rect 18325 7936 18337 7939
rect 18288 7908 18337 7936
rect 18288 7896 18294 7908
rect 18325 7905 18337 7908
rect 18371 7905 18383 7939
rect 18325 7899 18383 7905
rect 18414 7896 18420 7948
rect 18472 7936 18478 7948
rect 18785 7939 18843 7945
rect 18785 7936 18797 7939
rect 18472 7908 18797 7936
rect 18472 7896 18478 7908
rect 18785 7905 18797 7908
rect 18831 7905 18843 7939
rect 18785 7899 18843 7905
rect 21821 7871 21879 7877
rect 21821 7837 21833 7871
rect 21867 7868 21879 7871
rect 22554 7868 22560 7880
rect 21867 7840 22560 7868
rect 21867 7837 21879 7840
rect 21821 7831 21879 7837
rect 22554 7828 22560 7840
rect 22612 7828 22618 7880
rect 21361 7803 21419 7809
rect 21361 7769 21373 7803
rect 21407 7800 21419 7803
rect 21726 7800 21732 7812
rect 21407 7772 21732 7800
rect 21407 7769 21419 7772
rect 21361 7763 21419 7769
rect 21726 7760 21732 7772
rect 21784 7760 21790 7812
rect 22664 7800 22692 8044
rect 23477 8041 23489 8044
rect 23523 8072 23535 8075
rect 23842 8072 23848 8084
rect 23523 8044 23848 8072
rect 23523 8041 23535 8044
rect 23477 8035 23535 8041
rect 23842 8032 23848 8044
rect 23900 8032 23906 8084
rect 22738 7964 22744 8016
rect 22796 8004 22802 8016
rect 23753 8007 23811 8013
rect 23753 8004 23765 8007
rect 22796 7976 23765 8004
rect 22796 7964 22802 7976
rect 23753 7973 23765 7976
rect 23799 8004 23811 8007
rect 23934 8004 23940 8016
rect 23799 7976 23940 8004
rect 23799 7973 23811 7976
rect 23753 7967 23811 7973
rect 23934 7964 23940 7976
rect 23992 7964 23998 8016
rect 25184 7939 25242 7945
rect 25184 7905 25196 7939
rect 25230 7936 25242 7939
rect 25590 7936 25596 7948
rect 25230 7908 25596 7936
rect 25230 7905 25242 7908
rect 25184 7899 25242 7905
rect 25590 7896 25596 7908
rect 25648 7896 25654 7948
rect 23661 7871 23719 7877
rect 23661 7837 23673 7871
rect 23707 7868 23719 7871
rect 25038 7868 25044 7880
rect 23707 7840 25044 7868
rect 23707 7837 23719 7840
rect 23661 7831 23719 7837
rect 25038 7828 25044 7840
rect 25096 7868 25102 7880
rect 25271 7871 25329 7877
rect 25271 7868 25283 7871
rect 25096 7840 25283 7868
rect 25096 7828 25102 7840
rect 25271 7837 25283 7840
rect 25317 7837 25329 7871
rect 25271 7831 25329 7837
rect 22741 7803 22799 7809
rect 22741 7800 22753 7803
rect 22664 7772 22753 7800
rect 22741 7769 22753 7772
rect 22787 7769 22799 7803
rect 24210 7800 24216 7812
rect 24171 7772 24216 7800
rect 22741 7763 22799 7769
rect 24210 7760 24216 7772
rect 24268 7760 24274 7812
rect 13044 7704 15332 7732
rect 13044 7692 13050 7704
rect 21542 7692 21548 7744
rect 21600 7732 21606 7744
rect 21637 7735 21695 7741
rect 21637 7732 21649 7735
rect 21600 7704 21649 7732
rect 21600 7692 21606 7704
rect 21637 7701 21649 7704
rect 21683 7701 21695 7735
rect 21637 7695 21695 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 1719 7531 1777 7537
rect 1719 7528 1731 7531
rect 1636 7500 1731 7528
rect 1636 7488 1642 7500
rect 1719 7497 1731 7500
rect 1765 7497 1777 7531
rect 3970 7528 3976 7540
rect 3931 7500 3976 7528
rect 1719 7491 1777 7497
rect 3970 7488 3976 7500
rect 4028 7528 4034 7540
rect 4154 7528 4160 7540
rect 4028 7500 4160 7528
rect 4028 7488 4034 7500
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4338 7528 4344 7540
rect 4299 7500 4344 7528
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 6273 7531 6331 7537
rect 6273 7528 6285 7531
rect 5951 7500 6285 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 6273 7497 6285 7500
rect 6319 7528 6331 7531
rect 6638 7528 6644 7540
rect 6319 7500 6644 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 8527 7531 8585 7537
rect 8527 7528 8539 7531
rect 6788 7500 8539 7528
rect 6788 7488 6794 7500
rect 8527 7497 8539 7500
rect 8573 7497 8585 7531
rect 8527 7491 8585 7497
rect 8941 7531 8999 7537
rect 8941 7497 8953 7531
rect 8987 7528 8999 7531
rect 9582 7528 9588 7540
rect 8987 7500 9588 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 2225 7463 2283 7469
rect 2225 7429 2237 7463
rect 2271 7460 2283 7463
rect 2314 7460 2320 7472
rect 2271 7432 2320 7460
rect 2271 7429 2283 7432
rect 2225 7423 2283 7429
rect 2314 7420 2320 7432
rect 2372 7460 2378 7472
rect 3697 7463 3755 7469
rect 3697 7460 3709 7463
rect 2372 7432 3709 7460
rect 2372 7420 2378 7432
rect 3697 7429 3709 7432
rect 3743 7429 3755 7463
rect 8113 7463 8171 7469
rect 8113 7460 8125 7463
rect 3697 7423 3755 7429
rect 4126 7432 8125 7460
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 3050 7392 3056 7404
rect 2731 7364 3056 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 1648 7327 1706 7333
rect 1648 7293 1660 7327
rect 1694 7324 1706 7327
rect 2038 7324 2044 7336
rect 1694 7296 2044 7324
rect 1694 7293 1706 7296
rect 1648 7287 1706 7293
rect 2038 7284 2044 7296
rect 2096 7284 2102 7336
rect 2700 7256 2728 7355
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 3786 7324 3792 7336
rect 2823 7296 3792 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 3878 7284 3884 7336
rect 3936 7324 3942 7336
rect 4126 7324 4154 7432
rect 8113 7429 8125 7432
rect 8159 7460 8171 7463
rect 8386 7460 8392 7472
rect 8159 7432 8392 7460
rect 8159 7429 8171 7432
rect 8113 7423 8171 7429
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4948 7364 4997 7392
rect 4948 7352 4954 7364
rect 4985 7361 4997 7364
rect 5031 7392 5043 7395
rect 5442 7392 5448 7404
rect 5031 7364 5448 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 3936 7296 4154 7324
rect 6641 7327 6699 7333
rect 3936 7284 3942 7296
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 7006 7324 7012 7336
rect 6687 7296 7012 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7282 7324 7288 7336
rect 7243 7296 7288 7324
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 8456 7327 8514 7333
rect 8456 7293 8468 7327
rect 8502 7324 8514 7327
rect 8956 7324 8984 7491
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13320 7500 13461 7528
rect 13320 7488 13326 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14608 7500 15025 7528
rect 14608 7488 14614 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 16206 7528 16212 7540
rect 16167 7500 16212 7528
rect 15013 7491 15071 7497
rect 9490 7420 9496 7472
rect 9548 7460 9554 7472
rect 10137 7463 10195 7469
rect 10137 7460 10149 7463
rect 9548 7432 10149 7460
rect 9548 7420 9554 7432
rect 10137 7429 10149 7432
rect 10183 7429 10195 7463
rect 10137 7423 10195 7429
rect 11333 7463 11391 7469
rect 11333 7429 11345 7463
rect 11379 7460 11391 7463
rect 11606 7460 11612 7472
rect 11379 7432 11612 7460
rect 11379 7429 11391 7432
rect 11333 7423 11391 7429
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 12989 7463 13047 7469
rect 12989 7429 13001 7463
rect 13035 7460 13047 7463
rect 13630 7460 13636 7472
rect 13035 7432 13636 7460
rect 13035 7429 13047 7432
rect 12989 7423 13047 7429
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 9732 7364 10885 7392
rect 9732 7352 9738 7364
rect 10873 7361 10885 7364
rect 10919 7361 10931 7395
rect 10873 7355 10931 7361
rect 8502 7296 8984 7324
rect 8502 7293 8514 7296
rect 8456 7287 8514 7293
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 11112 7296 11161 7324
rect 11112 7284 11118 7296
rect 11149 7293 11161 7296
rect 11195 7324 11207 7327
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11195 7296 11989 7324
rect 11195 7293 11207 7296
rect 11149 7287 11207 7293
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 12504 7327 12562 7333
rect 12504 7293 12516 7327
rect 12550 7324 12562 7327
rect 12894 7324 12900 7336
rect 12550 7296 12900 7324
rect 12550 7293 12562 7296
rect 12504 7287 12562 7293
rect 12894 7284 12900 7296
rect 12952 7324 12958 7336
rect 13004 7324 13032 7423
rect 13630 7420 13636 7432
rect 13688 7420 13694 7472
rect 14274 7460 14280 7472
rect 13786 7432 14280 7460
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 13786 7392 13814 7432
rect 14274 7420 14280 7432
rect 14332 7420 14338 7472
rect 15028 7460 15056 7491
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 17083 7531 17141 7537
rect 17083 7497 17095 7531
rect 17129 7528 17141 7531
rect 17678 7528 17684 7540
rect 17129 7500 17684 7528
rect 17129 7497 17141 7500
rect 17083 7491 17141 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 18506 7488 18512 7540
rect 18564 7528 18570 7540
rect 19981 7531 20039 7537
rect 19981 7528 19993 7531
rect 18564 7500 19993 7528
rect 18564 7488 18570 7500
rect 19981 7497 19993 7500
rect 20027 7528 20039 7531
rect 20622 7528 20628 7540
rect 20027 7500 20628 7528
rect 20027 7497 20039 7500
rect 19981 7491 20039 7497
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 22830 7528 22836 7540
rect 22791 7500 22836 7528
rect 22830 7488 22836 7500
rect 22888 7488 22894 7540
rect 25038 7528 25044 7540
rect 24999 7500 25044 7528
rect 25038 7488 25044 7500
rect 25096 7488 25102 7540
rect 25590 7488 25596 7540
rect 25648 7528 25654 7540
rect 25685 7531 25743 7537
rect 25685 7528 25697 7531
rect 25648 7500 25697 7528
rect 25648 7488 25654 7500
rect 25685 7497 25697 7500
rect 25731 7497 25743 7531
rect 25685 7491 25743 7497
rect 17586 7460 17592 7472
rect 15028 7432 17592 7460
rect 13320 7364 13814 7392
rect 13320 7352 13326 7364
rect 12952 7296 13032 7324
rect 15028 7324 15056 7432
rect 17586 7420 17592 7432
rect 17644 7420 17650 7472
rect 17770 7420 17776 7472
rect 17828 7460 17834 7472
rect 17828 7432 20760 7460
rect 17828 7420 17834 7432
rect 15378 7352 15384 7404
rect 15436 7392 15442 7404
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 15436 7364 17877 7392
rect 15436 7352 15442 7364
rect 17865 7361 17877 7364
rect 17911 7392 17923 7395
rect 18414 7392 18420 7404
rect 17911 7364 18420 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 18414 7352 18420 7364
rect 18472 7352 18478 7404
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 19518 7392 19524 7404
rect 18739 7364 19524 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 19518 7352 19524 7364
rect 19576 7392 19582 7404
rect 20732 7401 20760 7432
rect 20806 7420 20812 7472
rect 20864 7460 20870 7472
rect 21082 7460 21088 7472
rect 20864 7432 21088 7460
rect 20864 7420 20870 7432
rect 21082 7420 21088 7432
rect 21140 7460 21146 7472
rect 21140 7432 25303 7460
rect 21140 7420 21146 7432
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 19576 7364 19625 7392
rect 19576 7352 19582 7364
rect 19613 7361 19625 7364
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7361 20775 7395
rect 24946 7392 24952 7404
rect 20717 7355 20775 7361
rect 20824 7364 24952 7392
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 15028 7296 15209 7324
rect 12952 7284 12958 7296
rect 15197 7293 15209 7296
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 15749 7327 15807 7333
rect 15749 7293 15761 7327
rect 15795 7324 15807 7327
rect 16758 7324 16764 7336
rect 15795 7296 16764 7324
rect 15795 7293 15807 7296
rect 15749 7287 15807 7293
rect 3098 7259 3156 7265
rect 3098 7256 3110 7259
rect 2700 7228 3110 7256
rect 3098 7225 3110 7228
rect 3144 7225 3156 7259
rect 9582 7256 9588 7268
rect 9543 7228 9588 7256
rect 3098 7219 3156 7225
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 9677 7259 9735 7265
rect 9677 7225 9689 7259
rect 9723 7256 9735 7259
rect 10042 7256 10048 7268
rect 9723 7228 10048 7256
rect 9723 7225 9735 7228
rect 9677 7219 9735 7225
rect 2866 7148 2872 7200
rect 2924 7188 2930 7200
rect 3326 7188 3332 7200
rect 2924 7160 3332 7188
rect 2924 7148 2930 7160
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 4893 7191 4951 7197
rect 4893 7188 4905 7191
rect 4580 7160 4905 7188
rect 4580 7148 4586 7160
rect 4893 7157 4905 7160
rect 4939 7188 4951 7191
rect 5350 7188 5356 7200
rect 4939 7160 5356 7188
rect 4939 7157 4951 7160
rect 4893 7151 4951 7157
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 6914 7188 6920 7200
rect 6875 7160 6920 7188
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 9401 7191 9459 7197
rect 9401 7157 9413 7191
rect 9447 7188 9459 7191
rect 9692 7188 9720 7219
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 13722 7256 13728 7268
rect 13683 7228 13728 7256
rect 13722 7216 13728 7228
rect 13780 7216 13786 7268
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 13872 7228 13917 7256
rect 13872 7216 13878 7228
rect 14642 7216 14648 7268
rect 14700 7256 14706 7268
rect 14737 7259 14795 7265
rect 14737 7256 14749 7259
rect 14700 7228 14749 7256
rect 14700 7216 14706 7228
rect 14737 7225 14749 7228
rect 14783 7256 14795 7259
rect 15764 7256 15792 7287
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 16942 7324 16948 7336
rect 17000 7333 17006 7336
rect 17000 7327 17038 7333
rect 16890 7296 16948 7324
rect 16942 7284 16948 7296
rect 17026 7324 17038 7327
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 17026 7296 17417 7324
rect 17026 7293 17038 7296
rect 17000 7287 17038 7293
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 20441 7327 20499 7333
rect 20441 7293 20453 7327
rect 20487 7293 20499 7327
rect 20622 7324 20628 7336
rect 20583 7296 20628 7324
rect 20441 7287 20499 7293
rect 17000 7284 17006 7287
rect 14783 7228 15792 7256
rect 16669 7259 16727 7265
rect 14783 7225 14795 7228
rect 14737 7219 14795 7225
rect 16669 7225 16681 7259
rect 16715 7256 16727 7259
rect 17310 7256 17316 7268
rect 16715 7228 17316 7256
rect 16715 7225 16727 7228
rect 16669 7219 16727 7225
rect 17310 7216 17316 7228
rect 17368 7256 17374 7268
rect 18138 7256 18144 7268
rect 17368 7228 18144 7256
rect 17368 7216 17374 7228
rect 18138 7216 18144 7228
rect 18196 7216 18202 7268
rect 18782 7216 18788 7268
rect 18840 7256 18846 7268
rect 18840 7228 18885 7256
rect 18840 7216 18846 7228
rect 19150 7216 19156 7268
rect 19208 7256 19214 7268
rect 19337 7259 19395 7265
rect 19337 7256 19349 7259
rect 19208 7228 19349 7256
rect 19208 7216 19214 7228
rect 19337 7225 19349 7228
rect 19383 7225 19395 7259
rect 19337 7219 19395 7225
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 20456 7256 20484 7287
rect 20622 7284 20628 7296
rect 20680 7324 20686 7336
rect 20824 7324 20852 7364
rect 24946 7352 24952 7364
rect 25004 7352 25010 7404
rect 20680 7296 20852 7324
rect 20680 7284 20686 7296
rect 21174 7284 21180 7336
rect 21232 7324 21238 7336
rect 21729 7327 21787 7333
rect 21729 7324 21741 7327
rect 21232 7296 21741 7324
rect 21232 7284 21238 7296
rect 21729 7293 21741 7296
rect 21775 7324 21787 7327
rect 22186 7324 22192 7336
rect 21775 7296 22192 7324
rect 21775 7293 21787 7296
rect 21729 7287 21787 7293
rect 22186 7284 22192 7296
rect 22244 7284 22250 7336
rect 22281 7327 22339 7333
rect 22281 7293 22293 7327
rect 22327 7324 22339 7327
rect 22830 7324 22836 7336
rect 22327 7296 22836 7324
rect 22327 7293 22339 7296
rect 22281 7287 22339 7293
rect 22830 7284 22836 7296
rect 22888 7284 22894 7336
rect 23382 7284 23388 7336
rect 23440 7324 23446 7336
rect 23474 7324 23480 7336
rect 23440 7296 23480 7324
rect 23440 7284 23446 7296
rect 23474 7284 23480 7296
rect 23532 7324 23538 7336
rect 25275 7333 25303 7432
rect 23661 7327 23719 7333
rect 23661 7324 23673 7327
rect 23532 7296 23673 7324
rect 23532 7284 23538 7296
rect 23661 7293 23673 7296
rect 23707 7293 23719 7327
rect 23661 7287 23719 7293
rect 24213 7327 24271 7333
rect 24213 7293 24225 7327
rect 24259 7324 24271 7327
rect 24673 7327 24731 7333
rect 24673 7324 24685 7327
rect 24259 7296 24685 7324
rect 24259 7293 24271 7296
rect 24213 7287 24271 7293
rect 24673 7293 24685 7296
rect 24719 7293 24731 7327
rect 24673 7287 24731 7293
rect 25260 7327 25318 7333
rect 25260 7293 25272 7327
rect 25306 7324 25318 7327
rect 26053 7327 26111 7333
rect 26053 7324 26065 7327
rect 25306 7296 26065 7324
rect 25306 7293 25318 7296
rect 25260 7287 25318 7293
rect 26053 7293 26065 7296
rect 26099 7293 26111 7327
rect 26053 7287 26111 7293
rect 22848 7256 22876 7284
rect 23106 7256 23112 7268
rect 20312 7228 21956 7256
rect 22848 7228 23112 7256
rect 20312 7216 20318 7228
rect 9447 7160 9720 7188
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10505 7191 10563 7197
rect 10505 7188 10517 7191
rect 10192 7160 10517 7188
rect 10192 7148 10198 7160
rect 10505 7157 10517 7160
rect 10551 7188 10563 7191
rect 11609 7191 11667 7197
rect 11609 7188 11621 7191
rect 10551 7160 11621 7188
rect 10551 7157 10563 7160
rect 10505 7151 10563 7157
rect 11609 7157 11621 7160
rect 11655 7188 11667 7191
rect 12526 7188 12532 7200
rect 11655 7160 12532 7188
rect 11655 7157 11667 7160
rect 11609 7151 11667 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12713 7191 12771 7197
rect 12713 7188 12725 7191
rect 12676 7160 12725 7188
rect 12676 7148 12682 7160
rect 12713 7157 12725 7160
rect 12759 7157 12771 7191
rect 15470 7188 15476 7200
rect 15431 7160 15476 7188
rect 12713 7151 12771 7157
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 18230 7188 18236 7200
rect 17920 7160 18236 7188
rect 17920 7148 17926 7160
rect 18230 7148 18236 7160
rect 18288 7188 18294 7200
rect 18417 7191 18475 7197
rect 18417 7188 18429 7191
rect 18288 7160 18429 7188
rect 18288 7148 18294 7160
rect 18417 7157 18429 7160
rect 18463 7188 18475 7191
rect 20272 7188 20300 7216
rect 21174 7188 21180 7200
rect 18463 7160 20300 7188
rect 21135 7160 21180 7188
rect 18463 7157 18475 7160
rect 18417 7151 18475 7157
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 21358 7148 21364 7200
rect 21416 7188 21422 7200
rect 21542 7188 21548 7200
rect 21416 7160 21548 7188
rect 21416 7148 21422 7160
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 21726 7148 21732 7200
rect 21784 7188 21790 7200
rect 21821 7191 21879 7197
rect 21821 7188 21833 7191
rect 21784 7160 21833 7188
rect 21784 7148 21790 7160
rect 21821 7157 21833 7160
rect 21867 7157 21879 7191
rect 21928 7188 21956 7228
rect 23106 7216 23112 7228
rect 23164 7256 23170 7268
rect 24118 7256 24124 7268
rect 23164 7228 24124 7256
rect 23164 7216 23170 7228
rect 24118 7216 24124 7228
rect 24176 7256 24182 7268
rect 24228 7256 24256 7287
rect 24176 7228 24256 7256
rect 24176 7216 24182 7228
rect 22922 7188 22928 7200
rect 21928 7160 22928 7188
rect 21821 7151 21879 7157
rect 22922 7148 22928 7160
rect 22980 7148 22986 7200
rect 23382 7188 23388 7200
rect 23343 7160 23388 7188
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 23750 7188 23756 7200
rect 23711 7160 23756 7188
rect 23750 7148 23756 7160
rect 23808 7148 23814 7200
rect 24762 7148 24768 7200
rect 24820 7188 24826 7200
rect 25363 7191 25421 7197
rect 25363 7188 25375 7191
rect 24820 7160 25375 7188
rect 24820 7148 24826 7160
rect 25363 7157 25375 7160
rect 25409 7157 25421 7191
rect 25363 7151 25421 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1946 6984 1952 6996
rect 1907 6956 1952 6984
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 3050 6984 3056 6996
rect 2648 6956 3056 6984
rect 2648 6944 2654 6956
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 3418 6984 3424 6996
rect 3379 6956 3424 6984
rect 3418 6944 3424 6956
rect 3476 6984 3482 6996
rect 4154 6984 4160 6996
rect 3476 6956 4160 6984
rect 3476 6944 3482 6956
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 5537 6987 5595 6993
rect 5537 6984 5549 6987
rect 4304 6956 5549 6984
rect 4304 6944 4310 6956
rect 5537 6953 5549 6956
rect 5583 6953 5595 6987
rect 6270 6984 6276 6996
rect 5537 6947 5595 6953
rect 5644 6956 6276 6984
rect 1464 6851 1522 6857
rect 1464 6817 1476 6851
rect 1510 6848 1522 6851
rect 1964 6848 1992 6944
rect 2222 6876 2228 6928
rect 2280 6916 2286 6928
rect 2866 6916 2872 6928
rect 2280 6888 2872 6916
rect 2280 6876 2286 6888
rect 2866 6876 2872 6888
rect 2924 6876 2930 6928
rect 3142 6916 3148 6928
rect 3103 6888 3148 6916
rect 3142 6876 3148 6888
rect 3200 6876 3206 6928
rect 4890 6916 4896 6928
rect 4851 6888 4896 6916
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 5644 6916 5672 6956
rect 6270 6944 6276 6956
rect 6328 6984 6334 6996
rect 7009 6987 7067 6993
rect 7009 6984 7021 6987
rect 6328 6956 7021 6984
rect 6328 6944 6334 6956
rect 7009 6953 7021 6956
rect 7055 6984 7067 6987
rect 7282 6984 7288 6996
rect 7055 6956 7288 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 7282 6944 7288 6956
rect 7340 6984 7346 6996
rect 8846 6984 8852 6996
rect 7340 6956 8852 6984
rect 7340 6944 7346 6956
rect 8846 6944 8852 6956
rect 8904 6944 8910 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 9769 6987 9827 6993
rect 9769 6984 9781 6987
rect 9732 6956 9781 6984
rect 9732 6944 9738 6956
rect 9769 6953 9781 6956
rect 9815 6953 9827 6987
rect 9769 6947 9827 6953
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 13725 6987 13783 6993
rect 9916 6956 13676 6984
rect 9916 6944 9922 6956
rect 5994 6916 6000 6928
rect 5460 6888 5672 6916
rect 5955 6888 6000 6916
rect 1510 6820 1992 6848
rect 2409 6851 2467 6857
rect 1510 6817 1522 6820
rect 1464 6811 1522 6817
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 2455 6820 3801 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 3789 6817 3801 6820
rect 3835 6848 3847 6851
rect 3878 6848 3884 6860
rect 3835 6820 3884 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4706 6848 4712 6860
rect 4212 6820 4257 6848
rect 4619 6820 4712 6848
rect 4212 6808 4218 6820
rect 4706 6808 4712 6820
rect 4764 6848 4770 6860
rect 5460 6848 5488 6888
rect 5994 6876 6000 6888
rect 6052 6876 6058 6928
rect 7650 6916 7656 6928
rect 6656 6888 7656 6916
rect 4764 6820 5488 6848
rect 4764 6808 4770 6820
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 6656 6857 6684 6888
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 9493 6919 9551 6925
rect 9493 6885 9505 6919
rect 9539 6916 9551 6919
rect 9582 6916 9588 6928
rect 9539 6888 9588 6916
rect 9539 6885 9551 6888
rect 9493 6879 9551 6885
rect 9582 6876 9588 6888
rect 9640 6916 9646 6928
rect 11379 6919 11437 6925
rect 11379 6916 11391 6919
rect 9640 6888 11391 6916
rect 9640 6876 9646 6888
rect 11379 6885 11391 6888
rect 11425 6885 11437 6919
rect 12710 6916 12716 6928
rect 12671 6888 12716 6916
rect 11379 6879 11437 6885
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 13262 6916 13268 6928
rect 13223 6888 13268 6916
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 13648 6916 13676 6956
rect 13725 6953 13737 6987
rect 13771 6984 13783 6987
rect 13814 6984 13820 6996
rect 13771 6956 13820 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 13814 6944 13820 6956
rect 13872 6944 13878 6996
rect 15427 6987 15485 6993
rect 15427 6953 15439 6987
rect 15473 6984 15485 6987
rect 17218 6984 17224 6996
rect 15473 6956 17224 6984
rect 15473 6953 15485 6956
rect 15427 6947 15485 6953
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 17402 6984 17408 6996
rect 17363 6956 17408 6984
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 18230 6984 18236 6996
rect 18191 6956 18236 6984
rect 18230 6944 18236 6956
rect 18288 6944 18294 6996
rect 18782 6984 18788 6996
rect 18743 6956 18788 6984
rect 18782 6944 18788 6956
rect 18840 6984 18846 6996
rect 19061 6987 19119 6993
rect 19061 6984 19073 6987
rect 18840 6956 19073 6984
rect 18840 6944 18846 6956
rect 19061 6953 19073 6956
rect 19107 6953 19119 6987
rect 19061 6947 19119 6953
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 19751 6987 19809 6993
rect 19751 6984 19763 6987
rect 19576 6956 19763 6984
rect 19576 6944 19582 6956
rect 19751 6953 19763 6956
rect 19797 6953 19809 6987
rect 20254 6984 20260 6996
rect 20215 6956 20260 6984
rect 19751 6947 19809 6953
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 22554 6944 22560 6996
rect 22612 6984 22618 6996
rect 22741 6987 22799 6993
rect 22741 6984 22753 6987
rect 22612 6956 22753 6984
rect 22612 6944 22618 6956
rect 22741 6953 22753 6956
rect 22787 6984 22799 6987
rect 22925 6987 22983 6993
rect 22925 6984 22937 6987
rect 22787 6956 22937 6984
rect 22787 6953 22799 6956
rect 22741 6947 22799 6953
rect 22925 6953 22937 6956
rect 22971 6953 22983 6987
rect 22925 6947 22983 6953
rect 23934 6944 23940 6996
rect 23992 6984 23998 6996
rect 24305 6987 24363 6993
rect 24305 6984 24317 6987
rect 23992 6956 24317 6984
rect 23992 6944 23998 6956
rect 24305 6953 24317 6956
rect 24351 6953 24363 6987
rect 24946 6984 24952 6996
rect 24907 6956 24952 6984
rect 24305 6947 24363 6953
rect 24946 6944 24952 6956
rect 25004 6944 25010 6996
rect 17862 6916 17868 6928
rect 13648 6888 17868 6916
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 21358 6876 21364 6928
rect 21416 6916 21422 6928
rect 21866 6919 21924 6925
rect 21866 6916 21878 6919
rect 21416 6888 21878 6916
rect 21416 6876 21422 6888
rect 21866 6885 21878 6888
rect 21912 6885 21924 6919
rect 23477 6919 23535 6925
rect 23477 6916 23489 6919
rect 21866 6879 21924 6885
rect 23124 6888 23489 6916
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 5592 6820 5733 6848
rect 5592 6808 5598 6820
rect 5721 6817 5733 6820
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6817 6699 6851
rect 9858 6848 9864 6860
rect 9819 6820 9864 6848
rect 6641 6811 6699 6817
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10134 6848 10140 6860
rect 10095 6820 10140 6848
rect 10134 6808 10140 6820
rect 10192 6848 10198 6860
rect 10689 6851 10747 6857
rect 10689 6848 10701 6851
rect 10192 6820 10701 6848
rect 10192 6808 10198 6820
rect 10689 6817 10701 6820
rect 10735 6817 10747 6851
rect 10689 6811 10747 6817
rect 11276 6851 11334 6857
rect 11276 6817 11288 6851
rect 11322 6817 11334 6851
rect 11276 6811 11334 6817
rect 14252 6851 14310 6857
rect 14252 6817 14264 6851
rect 14298 6848 14310 6851
rect 14550 6848 14556 6860
rect 14298 6820 14556 6848
rect 14298 6817 14310 6820
rect 14252 6811 14310 6817
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2648 6752 2789 6780
rect 2648 6740 2654 6752
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 2866 6740 2872 6792
rect 2924 6780 2930 6792
rect 2924 6752 5672 6780
rect 2924 6740 2930 6752
rect 1535 6715 1593 6721
rect 1535 6681 1547 6715
rect 1581 6712 1593 6715
rect 4890 6712 4896 6724
rect 1581 6684 4896 6712
rect 1581 6681 1593 6684
rect 1535 6675 1593 6681
rect 4890 6672 4896 6684
rect 4948 6672 4954 6724
rect 5644 6712 5672 6752
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 7190 6780 7196 6792
rect 6880 6752 7196 6780
rect 6880 6740 6886 6752
rect 7190 6740 7196 6752
rect 7248 6780 7254 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7248 6752 7573 6780
rect 7248 6740 7254 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 8849 6783 8907 6789
rect 8849 6780 8861 6783
rect 7561 6743 7619 6749
rect 7938 6752 8861 6780
rect 7938 6712 7966 6752
rect 8849 6749 8861 6752
rect 8895 6749 8907 6783
rect 8849 6743 8907 6749
rect 9950 6740 9956 6792
rect 10008 6780 10014 6792
rect 11291 6780 11319 6811
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 15197 6851 15255 6857
rect 15197 6817 15209 6851
rect 15243 6848 15255 6851
rect 15378 6848 15384 6860
rect 15243 6820 15384 6848
rect 15243 6817 15255 6820
rect 15197 6811 15255 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6817 16359 6851
rect 16758 6848 16764 6860
rect 16719 6820 16764 6848
rect 16301 6811 16359 6817
rect 11514 6780 11520 6792
rect 10008 6752 11520 6780
rect 10008 6740 10014 6752
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 12618 6780 12624 6792
rect 12579 6752 12624 6780
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 16206 6740 16212 6792
rect 16264 6780 16270 6792
rect 16316 6780 16344 6811
rect 16758 6808 16764 6820
rect 16816 6808 16822 6860
rect 19058 6808 19064 6860
rect 19116 6848 19122 6860
rect 19610 6848 19616 6860
rect 19668 6857 19674 6860
rect 19668 6851 19706 6857
rect 19116 6820 19616 6848
rect 19116 6808 19122 6820
rect 19610 6808 19616 6820
rect 19694 6817 19706 6851
rect 19668 6811 19706 6817
rect 19668 6808 19674 6811
rect 16264 6752 16344 6780
rect 17037 6783 17095 6789
rect 16264 6740 16270 6752
rect 17037 6749 17049 6783
rect 17083 6780 17095 6783
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17083 6752 17877 6780
rect 17083 6749 17095 6752
rect 17037 6743 17095 6749
rect 17865 6749 17877 6752
rect 17911 6780 17923 6783
rect 18414 6780 18420 6792
rect 17911 6752 18420 6780
rect 17911 6749 17923 6752
rect 17865 6743 17923 6749
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 22278 6780 22284 6792
rect 21591 6752 22284 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 5644 6684 7966 6712
rect 8018 6672 8024 6724
rect 8076 6712 8082 6724
rect 8113 6715 8171 6721
rect 8113 6712 8125 6715
rect 8076 6684 8125 6712
rect 8076 6672 8082 6684
rect 8113 6681 8125 6684
rect 8159 6681 8171 6715
rect 8113 6675 8171 6681
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 8573 6715 8631 6721
rect 8573 6712 8585 6715
rect 8536 6684 8585 6712
rect 8536 6672 8542 6684
rect 8573 6681 8585 6684
rect 8619 6712 8631 6715
rect 11422 6712 11428 6724
rect 8619 6684 11428 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 11532 6712 11560 6740
rect 16942 6712 16948 6724
rect 11532 6684 16948 6712
rect 16942 6672 16948 6684
rect 17000 6672 17006 6724
rect 23124 6721 23152 6888
rect 23477 6885 23489 6888
rect 23523 6885 23535 6919
rect 24026 6916 24032 6928
rect 23939 6888 24032 6916
rect 23477 6879 23535 6885
rect 24026 6876 24032 6888
rect 24084 6916 24090 6928
rect 24854 6916 24860 6928
rect 24084 6888 24860 6916
rect 24084 6876 24090 6888
rect 24854 6876 24860 6888
rect 24912 6876 24918 6928
rect 25130 6848 25136 6860
rect 25091 6820 25136 6848
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 25406 6848 25412 6860
rect 25367 6820 25412 6848
rect 25406 6808 25412 6820
rect 25464 6808 25470 6860
rect 23198 6740 23204 6792
rect 23256 6780 23262 6792
rect 23385 6783 23443 6789
rect 23385 6780 23397 6783
rect 23256 6752 23397 6780
rect 23256 6740 23262 6752
rect 23385 6749 23397 6752
rect 23431 6780 23443 6783
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 23431 6752 24685 6780
rect 23431 6749 23443 6752
rect 23385 6743 23443 6749
rect 24673 6749 24685 6752
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 22465 6715 22523 6721
rect 22465 6681 22477 6715
rect 22511 6712 22523 6715
rect 23109 6715 23167 6721
rect 23109 6712 23121 6715
rect 22511 6684 23121 6712
rect 22511 6681 22523 6684
rect 22465 6675 22523 6681
rect 23109 6681 23121 6684
rect 23155 6681 23167 6715
rect 23109 6675 23167 6681
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2406 6604 2412 6656
rect 2464 6644 2470 6656
rect 2547 6647 2605 6653
rect 2547 6644 2559 6647
rect 2464 6616 2559 6644
rect 2464 6604 2470 6616
rect 2547 6613 2559 6616
rect 2593 6613 2605 6647
rect 2682 6644 2688 6656
rect 2643 6616 2688 6644
rect 2547 6607 2605 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 7282 6644 7288 6656
rect 7243 6616 7288 6644
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11296 6616 11713 6644
rect 11296 6604 11302 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13872 6616 14105 6644
rect 13872 6604 13878 6616
rect 14093 6613 14105 6616
rect 14139 6644 14151 6647
rect 14323 6647 14381 6653
rect 14323 6644 14335 6647
rect 14139 6616 14335 6644
rect 14139 6613 14151 6616
rect 14093 6607 14151 6613
rect 14323 6613 14335 6616
rect 14369 6613 14381 6647
rect 15746 6644 15752 6656
rect 15707 6616 15752 6644
rect 14323 6607 14381 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6644 16267 6647
rect 16482 6644 16488 6656
rect 16255 6616 16488 6644
rect 16255 6613 16267 6616
rect 16209 6607 16267 6613
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 17770 6644 17776 6656
rect 17731 6616 17776 6644
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 21453 6647 21511 6653
rect 21453 6613 21465 6647
rect 21499 6644 21511 6647
rect 21542 6644 21548 6656
rect 21499 6616 21548 6644
rect 21499 6613 21511 6616
rect 21453 6607 21511 6613
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 22925 6647 22983 6653
rect 22925 6613 22937 6647
rect 22971 6644 22983 6647
rect 23750 6644 23756 6656
rect 22971 6616 23756 6644
rect 22971 6613 22983 6616
rect 22925 6607 22983 6613
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 3053 6443 3111 6449
rect 3053 6440 3065 6443
rect 2740 6412 3065 6440
rect 2740 6400 2746 6412
rect 3053 6409 3065 6412
rect 3099 6409 3111 6443
rect 4154 6440 4160 6452
rect 3053 6403 3111 6409
rect 4126 6400 4160 6440
rect 4212 6440 4218 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 4212 6412 4261 6440
rect 4212 6400 4218 6412
rect 4249 6409 4261 6412
rect 4295 6409 4307 6443
rect 4249 6403 4307 6409
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 5592 6412 6193 6440
rect 5592 6400 5598 6412
rect 6181 6409 6193 6412
rect 6227 6409 6239 6443
rect 6181 6403 6239 6409
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 7285 6443 7343 6449
rect 7285 6440 7297 6443
rect 7248 6412 7297 6440
rect 7248 6400 7254 6412
rect 7285 6409 7297 6412
rect 7331 6409 7343 6443
rect 7285 6403 7343 6409
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 7708 6412 8493 6440
rect 7708 6400 7714 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 8628 6412 8953 6440
rect 8628 6400 8634 6412
rect 8941 6409 8953 6412
rect 8987 6440 8999 6443
rect 10134 6440 10140 6452
rect 8987 6412 10140 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11514 6440 11520 6452
rect 11475 6412 11520 6440
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12710 6440 12716 6452
rect 12299 6412 12716 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 16206 6400 16212 6452
rect 16264 6440 16270 6452
rect 16301 6443 16359 6449
rect 16301 6440 16313 6443
rect 16264 6412 16313 6440
rect 16264 6400 16270 6412
rect 16301 6409 16313 6412
rect 16347 6409 16359 6443
rect 16301 6403 16359 6409
rect 16991 6443 17049 6449
rect 16991 6409 17003 6443
rect 17037 6440 17049 6443
rect 17126 6440 17132 6452
rect 17037 6412 17132 6440
rect 17037 6409 17049 6412
rect 16991 6403 17049 6409
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6440 17279 6443
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 17267 6412 17417 6440
rect 17267 6409 17279 6412
rect 17221 6403 17279 6409
rect 17405 6409 17417 6412
rect 17451 6440 17463 6443
rect 22925 6443 22983 6449
rect 22925 6440 22937 6443
rect 17451 6412 22937 6440
rect 17451 6409 17463 6412
rect 17405 6403 17463 6409
rect 22925 6409 22937 6412
rect 22971 6409 22983 6443
rect 22925 6403 22983 6409
rect 23106 6400 23112 6452
rect 23164 6440 23170 6452
rect 23164 6412 23209 6440
rect 23164 6400 23170 6412
rect 23290 6400 23296 6452
rect 23348 6440 23354 6452
rect 23385 6443 23443 6449
rect 23385 6440 23397 6443
rect 23348 6412 23397 6440
rect 23348 6400 23354 6412
rect 23385 6409 23397 6412
rect 23431 6409 23443 6443
rect 23385 6403 23443 6409
rect 23566 6400 23572 6452
rect 23624 6440 23630 6452
rect 27614 6440 27620 6452
rect 23624 6412 27620 6440
rect 23624 6400 23630 6412
rect 27614 6400 27620 6412
rect 27672 6400 27678 6452
rect 4126 6372 4154 6400
rect 4706 6372 4712 6384
rect 3712 6344 4154 6372
rect 4667 6344 4712 6372
rect 3712 6304 3740 6344
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 5074 6332 5080 6384
rect 5132 6372 5138 6384
rect 5350 6372 5356 6384
rect 5132 6344 5356 6372
rect 5132 6332 5138 6344
rect 5350 6332 5356 6344
rect 5408 6372 5414 6384
rect 5905 6375 5963 6381
rect 5905 6372 5917 6375
rect 5408 6344 5917 6372
rect 5408 6332 5414 6344
rect 5905 6341 5917 6344
rect 5951 6372 5963 6375
rect 5994 6372 6000 6384
rect 5951 6344 6000 6372
rect 5951 6341 5963 6344
rect 5905 6335 5963 6341
rect 5994 6332 6000 6344
rect 6052 6372 6058 6384
rect 7466 6372 7472 6384
rect 6052 6344 7472 6372
rect 6052 6332 6058 6344
rect 7466 6332 7472 6344
rect 7524 6332 7530 6384
rect 9398 6372 9404 6384
rect 9311 6344 9404 6372
rect 9398 6332 9404 6344
rect 9456 6372 9462 6384
rect 9858 6372 9864 6384
rect 9456 6344 9864 6372
rect 9456 6332 9462 6344
rect 9858 6332 9864 6344
rect 9916 6332 9922 6384
rect 10152 6372 10180 6400
rect 14366 6372 14372 6384
rect 10152 6344 10640 6372
rect 14327 6344 14372 6372
rect 3528 6276 3740 6304
rect 2038 6236 2044 6248
rect 1999 6208 2044 6236
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 3528 6245 3556 6276
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 4890 6304 4896 6316
rect 3844 6276 3889 6304
rect 4803 6276 4896 6304
rect 3844 6264 3850 6276
rect 4890 6264 4896 6276
rect 4948 6304 4954 6316
rect 7282 6304 7288 6316
rect 4948 6276 7288 6304
rect 4948 6264 4954 6276
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7386 6276 7573 6304
rect 3513 6239 3571 6245
rect 3513 6205 3525 6239
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6236 3755 6239
rect 4062 6236 4068 6248
rect 3743 6208 4068 6236
rect 3743 6205 3755 6208
rect 3697 6199 3755 6205
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 7386 6236 7414 6276
rect 7561 6273 7573 6276
rect 7607 6304 7619 6307
rect 8202 6304 8208 6316
rect 7607 6276 8208 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 10318 6304 10324 6316
rect 10279 6276 10324 6304
rect 10318 6264 10324 6276
rect 10376 6304 10382 6316
rect 10376 6276 10548 6304
rect 10376 6264 10382 6276
rect 9490 6236 9496 6248
rect 5592 6208 7414 6236
rect 9451 6208 9496 6236
rect 5592 6196 5598 6208
rect 9490 6196 9496 6208
rect 9548 6236 9554 6248
rect 10520 6245 10548 6276
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9548 6208 9965 6236
rect 9548 6196 9554 6208
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 10505 6239 10563 6245
rect 10505 6205 10517 6239
rect 10551 6205 10563 6239
rect 10612 6236 10640 6344
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 14734 6332 14740 6384
rect 14792 6372 14798 6384
rect 24762 6372 24768 6384
rect 14792 6344 24768 6372
rect 14792 6332 14798 6344
rect 24762 6332 24768 6344
rect 24820 6332 24826 6384
rect 24949 6375 25007 6381
rect 24949 6341 24961 6375
rect 24995 6372 25007 6375
rect 25130 6372 25136 6384
rect 24995 6344 25136 6372
rect 24995 6341 25007 6344
rect 24949 6335 25007 6341
rect 25130 6332 25136 6344
rect 25188 6332 25194 6384
rect 25409 6375 25467 6381
rect 25409 6341 25421 6375
rect 25455 6372 25467 6375
rect 26602 6372 26608 6384
rect 25455 6344 26608 6372
rect 25455 6341 25467 6344
rect 25409 6335 25467 6341
rect 26602 6332 26608 6344
rect 26660 6332 26666 6384
rect 11238 6304 11244 6316
rect 11199 6276 11244 6304
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 15194 6304 15200 6316
rect 13872 6276 13917 6304
rect 15155 6276 15200 6304
rect 13872 6264 13878 6276
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6304 15439 6307
rect 16482 6304 16488 6316
rect 15427 6276 16488 6304
rect 15427 6273 15439 6276
rect 15381 6267 15439 6273
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 17770 6264 17776 6316
rect 17828 6304 17834 6316
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 17828 6276 18153 6304
rect 17828 6264 17834 6276
rect 18141 6273 18153 6276
rect 18187 6304 18199 6307
rect 20441 6307 20499 6313
rect 20441 6304 20453 6307
rect 18187 6276 20453 6304
rect 18187 6273 18199 6276
rect 18141 6267 18199 6273
rect 20441 6273 20453 6276
rect 20487 6273 20499 6307
rect 20441 6267 20499 6273
rect 22925 6307 22983 6313
rect 22925 6273 22937 6307
rect 22971 6304 22983 6307
rect 23474 6304 23480 6316
rect 22971 6276 23480 6304
rect 22971 6273 22983 6276
rect 22925 6267 22983 6273
rect 23474 6264 23480 6276
rect 23532 6264 23538 6316
rect 24026 6264 24032 6316
rect 24084 6304 24090 6316
rect 25777 6307 25835 6313
rect 25777 6304 25789 6307
rect 24084 6276 25789 6304
rect 24084 6264 24090 6276
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10612 6208 10977 6236
rect 10505 6199 10563 6205
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 10965 6199 11023 6205
rect 12780 6239 12838 6245
rect 12780 6205 12792 6239
rect 12826 6236 12838 6239
rect 13170 6236 13176 6248
rect 12826 6208 13176 6236
rect 12826 6205 12838 6208
rect 12780 6199 12838 6205
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 14550 6196 14556 6248
rect 14608 6236 14614 6248
rect 14737 6239 14795 6245
rect 14737 6236 14749 6239
rect 14608 6208 14749 6236
rect 14608 6196 14614 6208
rect 14737 6205 14749 6208
rect 14783 6205 14795 6239
rect 14737 6199 14795 6205
rect 16920 6239 16978 6245
rect 16920 6205 16932 6239
rect 16966 6236 16978 6239
rect 17221 6239 17279 6245
rect 17221 6236 17233 6239
rect 16966 6208 17233 6236
rect 16966 6205 16978 6208
rect 16920 6199 16978 6205
rect 17221 6205 17233 6208
rect 17267 6205 17279 6239
rect 17221 6199 17279 6205
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18230 6236 18236 6248
rect 17920 6208 18236 6236
rect 17920 6196 17926 6208
rect 18230 6196 18236 6208
rect 18288 6236 18294 6248
rect 19426 6236 19432 6248
rect 18288 6208 19432 6236
rect 18288 6196 18294 6208
rect 2409 6171 2467 6177
rect 2409 6137 2421 6171
rect 2455 6168 2467 6171
rect 2590 6168 2596 6180
rect 2455 6140 2596 6168
rect 2455 6137 2467 6140
rect 2409 6131 2467 6137
rect 2590 6128 2596 6140
rect 2648 6128 2654 6180
rect 3786 6128 3792 6180
rect 3844 6168 3850 6180
rect 3970 6168 3976 6180
rect 3844 6140 3976 6168
rect 3844 6128 3850 6140
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 4985 6171 5043 6177
rect 4985 6137 4997 6171
rect 5031 6168 5043 6171
rect 5166 6168 5172 6180
rect 5031 6140 5172 6168
rect 5031 6137 5043 6140
rect 4985 6131 5043 6137
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 6641 6171 6699 6177
rect 6641 6137 6653 6171
rect 6687 6168 6699 6171
rect 7653 6171 7711 6177
rect 6687 6140 7414 6168
rect 6687 6137 6699 6140
rect 6641 6131 6699 6137
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 2866 6100 2872 6112
rect 2823 6072 2872 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 7386 6100 7414 6140
rect 7653 6137 7665 6171
rect 7699 6137 7711 6171
rect 7653 6131 7711 6137
rect 7668 6100 7696 6131
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 8205 6171 8263 6177
rect 8205 6168 8217 6171
rect 8076 6140 8217 6168
rect 8076 6128 8082 6140
rect 8205 6137 8217 6140
rect 8251 6137 8263 6171
rect 8205 6131 8263 6137
rect 11238 6128 11244 6180
rect 11296 6168 11302 6180
rect 12986 6168 12992 6180
rect 11296 6140 12992 6168
rect 11296 6128 11302 6140
rect 12986 6128 12992 6140
rect 13044 6128 13050 6180
rect 13909 6171 13967 6177
rect 13909 6137 13921 6171
rect 13955 6137 13967 6171
rect 15473 6171 15531 6177
rect 15473 6168 15485 6171
rect 13909 6131 13967 6137
rect 14568 6140 15485 6168
rect 7926 6100 7932 6112
rect 7386 6072 7932 6100
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 9950 6100 9956 6112
rect 9723 6072 9956 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 12851 6103 12909 6109
rect 12851 6069 12863 6103
rect 12897 6100 12909 6103
rect 13078 6100 13084 6112
rect 12897 6072 13084 6100
rect 12897 6069 12909 6072
rect 12851 6063 12909 6069
rect 13078 6060 13084 6072
rect 13136 6060 13142 6112
rect 13633 6103 13691 6109
rect 13633 6069 13645 6103
rect 13679 6100 13691 6103
rect 13924 6100 13952 6131
rect 14568 6100 14596 6140
rect 15473 6137 15485 6140
rect 15519 6168 15531 6171
rect 15746 6168 15752 6180
rect 15519 6140 15752 6168
rect 15519 6137 15531 6140
rect 15473 6131 15531 6137
rect 15746 6128 15752 6140
rect 15804 6128 15810 6180
rect 16025 6171 16083 6177
rect 16025 6137 16037 6171
rect 16071 6168 16083 6171
rect 16206 6168 16212 6180
rect 16071 6140 16212 6168
rect 16071 6137 16083 6140
rect 16025 6131 16083 6137
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 16758 6168 16764 6180
rect 16671 6140 16764 6168
rect 16758 6128 16764 6140
rect 16816 6168 16822 6180
rect 18477 6177 18505 6208
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 19610 6236 19616 6248
rect 19571 6208 19616 6236
rect 19610 6196 19616 6208
rect 19668 6196 19674 6248
rect 19978 6236 19984 6248
rect 19939 6208 19984 6236
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 20346 6236 20352 6248
rect 20307 6208 20352 6236
rect 20346 6196 20352 6208
rect 20404 6196 20410 6248
rect 21542 6236 21548 6248
rect 21503 6208 21548 6236
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 23290 6196 23296 6248
rect 23348 6236 23354 6248
rect 23566 6236 23572 6248
rect 23348 6208 23572 6236
rect 23348 6196 23354 6208
rect 23566 6196 23572 6208
rect 23624 6236 23630 6248
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 23624 6208 23673 6236
rect 23624 6196 23630 6208
rect 23661 6205 23673 6208
rect 23707 6205 23719 6239
rect 24118 6236 24124 6248
rect 24079 6208 24124 6236
rect 23661 6199 23719 6205
rect 24118 6196 24124 6208
rect 24176 6196 24182 6248
rect 25240 6245 25268 6276
rect 25777 6273 25789 6276
rect 25823 6273 25835 6307
rect 25777 6267 25835 6273
rect 25225 6239 25283 6245
rect 25225 6205 25237 6239
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 18462 6171 18520 6177
rect 16816 6140 18229 6168
rect 16816 6128 16822 6140
rect 17862 6100 17868 6112
rect 13679 6072 14596 6100
rect 17823 6072 17868 6100
rect 13679 6069 13691 6072
rect 13633 6063 13691 6069
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 18201 6100 18229 6140
rect 18462 6137 18474 6171
rect 18508 6137 18520 6171
rect 20364 6168 20392 6196
rect 18462 6131 18520 6137
rect 18616 6140 20392 6168
rect 21866 6171 21924 6177
rect 18616 6100 18644 6140
rect 21866 6137 21878 6171
rect 21912 6137 21924 6171
rect 21866 6131 21924 6137
rect 19058 6100 19064 6112
rect 18201 6072 18644 6100
rect 19019 6072 19064 6100
rect 19058 6060 19064 6072
rect 19116 6060 19122 6112
rect 19426 6060 19432 6112
rect 19484 6100 19490 6112
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 19484 6072 21005 6100
rect 19484 6060 19490 6072
rect 20993 6069 21005 6072
rect 21039 6100 21051 6103
rect 21082 6100 21088 6112
rect 21039 6072 21088 6100
rect 21039 6069 21051 6072
rect 20993 6063 21051 6069
rect 21082 6060 21088 6072
rect 21140 6100 21146 6112
rect 21358 6100 21364 6112
rect 21140 6072 21364 6100
rect 21140 6060 21146 6072
rect 21358 6060 21364 6072
rect 21416 6100 21422 6112
rect 21881 6100 21909 6131
rect 22462 6100 22468 6112
rect 21416 6072 21909 6100
rect 22423 6072 22468 6100
rect 21416 6060 21422 6072
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 23750 6100 23756 6112
rect 23711 6072 23756 6100
rect 23750 6060 23756 6072
rect 23808 6060 23814 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3053 5899 3111 5905
rect 3053 5896 3065 5899
rect 3016 5868 3065 5896
rect 3016 5856 3022 5868
rect 3053 5865 3065 5868
rect 3099 5865 3111 5899
rect 3053 5859 3111 5865
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 3326 5896 3332 5908
rect 3283 5868 3332 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 4709 5899 4767 5905
rect 4709 5865 4721 5899
rect 4755 5896 4767 5899
rect 5074 5896 5080 5908
rect 4755 5868 5080 5896
rect 4755 5865 4767 5868
rect 4709 5859 4767 5865
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5261 5899 5319 5905
rect 5261 5896 5273 5899
rect 5224 5868 5273 5896
rect 5224 5856 5230 5868
rect 5261 5865 5273 5868
rect 5307 5865 5319 5899
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 5261 5859 5319 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 7248 5868 7389 5896
rect 7248 5856 7254 5868
rect 7377 5865 7389 5868
rect 7423 5896 7435 5899
rect 7466 5896 7472 5908
rect 7423 5868 7472 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 7926 5896 7932 5908
rect 7887 5868 7932 5896
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 8202 5896 8208 5908
rect 8163 5868 8208 5896
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 13078 5856 13084 5908
rect 13136 5896 13142 5908
rect 13449 5899 13507 5905
rect 13449 5896 13461 5899
rect 13136 5868 13461 5896
rect 13136 5856 13142 5868
rect 13449 5865 13461 5868
rect 13495 5865 13507 5899
rect 13449 5859 13507 5865
rect 1535 5831 1593 5837
rect 1535 5797 1547 5831
rect 1581 5828 1593 5831
rect 3602 5828 3608 5840
rect 1581 5800 3608 5828
rect 1581 5797 1593 5800
rect 1535 5791 1593 5797
rect 3602 5788 3608 5800
rect 3660 5788 3666 5840
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 6273 5831 6331 5837
rect 6273 5828 6285 5831
rect 4856 5800 6285 5828
rect 4856 5788 4862 5800
rect 6273 5797 6285 5800
rect 6319 5797 6331 5831
rect 6273 5791 6331 5797
rect 9950 5788 9956 5840
rect 10008 5828 10014 5840
rect 11054 5828 11060 5840
rect 10008 5800 10732 5828
rect 11015 5800 11060 5828
rect 10008 5788 10014 5800
rect 658 5720 664 5772
rect 716 5760 722 5772
rect 1432 5763 1490 5769
rect 1432 5760 1444 5763
rect 716 5732 1444 5760
rect 716 5720 722 5732
rect 1432 5729 1444 5732
rect 1478 5760 1490 5763
rect 1670 5760 1676 5772
rect 1478 5732 1676 5760
rect 1478 5729 1490 5732
rect 1432 5723 1490 5729
rect 1670 5720 1676 5732
rect 1728 5720 1734 5772
rect 2314 5720 2320 5772
rect 2372 5760 2378 5772
rect 2409 5763 2467 5769
rect 2409 5760 2421 5763
rect 2372 5732 2421 5760
rect 2372 5720 2378 5732
rect 2409 5729 2421 5732
rect 2455 5760 2467 5763
rect 3326 5760 3332 5772
rect 2455 5732 3332 5760
rect 2455 5729 2467 5732
rect 2409 5723 2467 5729
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 3878 5720 3884 5772
rect 3936 5760 3942 5772
rect 9030 5760 9036 5772
rect 3936 5732 9036 5760
rect 3936 5720 3942 5732
rect 9030 5720 9036 5732
rect 9088 5760 9094 5772
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 9088 5732 10149 5760
rect 9088 5720 9094 5732
rect 10137 5729 10149 5732
rect 10183 5760 10195 5763
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 10183 5732 10333 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 10321 5729 10333 5732
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 2590 5652 2596 5704
rect 2648 5692 2654 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2648 5664 2789 5692
rect 2648 5652 2654 5664
rect 2777 5661 2789 5664
rect 2823 5692 2835 5695
rect 2823 5664 3924 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 2314 5624 2320 5636
rect 2227 5596 2320 5624
rect 2314 5584 2320 5596
rect 2372 5624 2378 5636
rect 2866 5624 2872 5636
rect 2372 5596 2872 5624
rect 2372 5584 2378 5596
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 2038 5556 2044 5568
rect 1995 5528 2044 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 2562 5565 2590 5596
rect 2866 5584 2872 5596
rect 2924 5624 2930 5636
rect 3602 5624 3608 5636
rect 2924 5596 3608 5624
rect 2924 5584 2930 5596
rect 3602 5584 3608 5596
rect 3660 5584 3666 5636
rect 2547 5559 2605 5565
rect 2547 5556 2559 5559
rect 2525 5528 2559 5556
rect 2547 5525 2559 5528
rect 2593 5525 2605 5559
rect 2547 5519 2605 5525
rect 2685 5559 2743 5565
rect 2685 5525 2697 5559
rect 2731 5556 2743 5559
rect 2958 5556 2964 5568
rect 2731 5528 2964 5556
rect 2731 5525 2743 5528
rect 2685 5519 2743 5525
rect 2958 5516 2964 5528
rect 3016 5556 3022 5568
rect 3237 5559 3295 5565
rect 3237 5556 3249 5559
rect 3016 5528 3249 5556
rect 3016 5516 3022 5528
rect 3237 5525 3249 5528
rect 3283 5525 3295 5559
rect 3237 5519 3295 5525
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 3896 5565 3924 5664
rect 3970 5652 3976 5704
rect 4028 5692 4034 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 4028 5664 4353 5692
rect 4028 5652 4034 5664
rect 4341 5661 4353 5664
rect 4387 5692 4399 5695
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 4387 5664 5549 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 6270 5652 6276 5704
rect 6328 5692 6334 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6328 5664 7021 5692
rect 6328 5652 6334 5664
rect 7009 5661 7021 5664
rect 7055 5692 7067 5695
rect 8662 5692 8668 5704
rect 7055 5664 8668 5692
rect 7055 5661 7067 5664
rect 7009 5655 7067 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 10704 5701 10732 5800
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 13464 5828 13492 5859
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 14550 5896 14556 5908
rect 14056 5868 14556 5896
rect 14056 5856 14062 5868
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 15654 5896 15660 5908
rect 15615 5868 15660 5896
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 16209 5899 16267 5905
rect 16209 5865 16221 5899
rect 16255 5896 16267 5899
rect 18414 5896 18420 5908
rect 16255 5868 17264 5896
rect 18375 5868 18420 5896
rect 16255 5865 16267 5868
rect 16209 5859 16267 5865
rect 17236 5840 17264 5868
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 18616 5868 21005 5896
rect 13725 5831 13783 5837
rect 13725 5828 13737 5831
rect 13464 5800 13737 5828
rect 13725 5797 13737 5800
rect 13771 5797 13783 5831
rect 13725 5791 13783 5797
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 14366 5828 14372 5840
rect 13872 5800 13917 5828
rect 14327 5800 14372 5828
rect 13872 5788 13878 5800
rect 14366 5788 14372 5800
rect 14424 5788 14430 5840
rect 17218 5828 17224 5840
rect 17131 5800 17224 5828
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 12342 5760 12348 5772
rect 12303 5732 12348 5760
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 12526 5760 12532 5772
rect 12487 5732 12532 5760
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 12618 5720 12624 5772
rect 12676 5760 12682 5772
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 12676 5732 13093 5760
rect 12676 5720 12682 5732
rect 13081 5729 13093 5732
rect 13127 5729 13139 5763
rect 13081 5723 13139 5729
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 10870 5692 10876 5704
rect 10735 5664 10876 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 14826 5692 14832 5704
rect 12851 5664 13676 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 10597 5627 10655 5633
rect 10597 5624 10609 5627
rect 9732 5596 10609 5624
rect 9732 5584 9738 5596
rect 10597 5593 10609 5596
rect 10643 5593 10655 5627
rect 13648 5624 13676 5664
rect 13786 5664 14832 5692
rect 13786 5624 13814 5664
rect 14826 5652 14832 5664
rect 14884 5692 14890 5704
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14884 5664 15301 5692
rect 14884 5652 14890 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 17126 5692 17132 5704
rect 17087 5664 17132 5692
rect 15289 5655 15347 5661
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 18616 5692 18644 5868
rect 20993 5865 21005 5868
rect 21039 5865 21051 5899
rect 20993 5859 21051 5865
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 24213 5899 24271 5905
rect 24213 5896 24225 5899
rect 21600 5868 24225 5896
rect 21600 5856 21606 5868
rect 24213 5865 24225 5868
rect 24259 5865 24271 5899
rect 24213 5859 24271 5865
rect 19058 5828 19064 5840
rect 18971 5800 19064 5828
rect 19058 5788 19064 5800
rect 19116 5828 19122 5840
rect 19610 5828 19616 5840
rect 19116 5800 19616 5828
rect 19116 5788 19122 5800
rect 19610 5788 19616 5800
rect 19668 5788 19674 5840
rect 19978 5828 19984 5840
rect 19939 5800 19984 5828
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 20346 5828 20352 5840
rect 20259 5800 20352 5828
rect 20346 5788 20352 5800
rect 20404 5828 20410 5840
rect 22278 5828 22284 5840
rect 20404 5800 21312 5828
rect 22239 5800 22284 5828
rect 20404 5788 20410 5800
rect 21284 5772 21312 5800
rect 22278 5788 22284 5800
rect 22336 5788 22342 5840
rect 22462 5788 22468 5840
rect 22520 5828 22526 5840
rect 22741 5831 22799 5837
rect 22741 5828 22753 5831
rect 22520 5800 22753 5828
rect 22520 5788 22526 5800
rect 22741 5797 22753 5800
rect 22787 5797 22799 5831
rect 22741 5791 22799 5797
rect 23293 5831 23351 5837
rect 23293 5797 23305 5831
rect 23339 5828 23351 5831
rect 23934 5828 23940 5840
rect 23339 5800 23940 5828
rect 23339 5797 23351 5800
rect 23293 5791 23351 5797
rect 23934 5788 23940 5800
rect 23992 5788 23998 5840
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 18966 5692 18972 5704
rect 17236 5664 18644 5692
rect 18927 5664 18972 5692
rect 14734 5624 14740 5636
rect 13648 5596 13814 5624
rect 14647 5596 14740 5624
rect 10597 5587 10655 5593
rect 14734 5584 14740 5596
rect 14792 5624 14798 5636
rect 17236 5624 17264 5664
rect 18966 5652 18972 5664
rect 19024 5652 19030 5704
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 17678 5624 17684 5636
rect 14792 5596 17264 5624
rect 17639 5596 17684 5624
rect 14792 5584 14798 5596
rect 17678 5584 17684 5596
rect 17736 5624 17742 5636
rect 19150 5624 19156 5636
rect 17736 5596 19156 5624
rect 17736 5584 17742 5596
rect 19150 5584 19156 5596
rect 19208 5624 19214 5636
rect 19260 5624 19288 5655
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 20714 5692 20720 5704
rect 19484 5664 20720 5692
rect 19484 5652 19490 5664
rect 20714 5652 20720 5664
rect 20772 5692 20778 5704
rect 20916 5692 20944 5723
rect 21266 5720 21272 5772
rect 21324 5760 21330 5772
rect 21361 5763 21419 5769
rect 21361 5760 21373 5763
rect 21324 5732 21373 5760
rect 21324 5720 21330 5732
rect 21361 5729 21373 5732
rect 21407 5729 21419 5763
rect 21361 5723 21419 5729
rect 23566 5720 23572 5772
rect 23624 5760 23630 5772
rect 24118 5760 24124 5772
rect 23624 5732 24124 5760
rect 23624 5720 23630 5732
rect 24118 5720 24124 5732
rect 24176 5720 24182 5772
rect 24581 5763 24639 5769
rect 24581 5729 24593 5763
rect 24627 5729 24639 5763
rect 24581 5723 24639 5729
rect 22186 5692 22192 5704
rect 20772 5664 22192 5692
rect 20772 5652 20778 5664
rect 22186 5652 22192 5664
rect 22244 5652 22250 5704
rect 22646 5692 22652 5704
rect 22607 5664 22652 5692
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 24596 5692 24624 5723
rect 23768 5664 24624 5692
rect 19208 5596 19288 5624
rect 22005 5627 22063 5633
rect 19208 5584 19214 5596
rect 22005 5593 22017 5627
rect 22051 5624 22063 5627
rect 22738 5624 22744 5636
rect 22051 5596 22744 5624
rect 22051 5593 22063 5596
rect 22005 5587 22063 5593
rect 22738 5584 22744 5596
rect 22796 5584 22802 5636
rect 23768 5568 23796 5664
rect 3421 5559 3479 5565
rect 3421 5556 3433 5559
rect 3384 5528 3433 5556
rect 3384 5516 3390 5528
rect 3421 5525 3433 5528
rect 3467 5525 3479 5559
rect 3421 5519 3479 5525
rect 3881 5559 3939 5565
rect 3881 5525 3893 5559
rect 3927 5556 3939 5559
rect 4062 5556 4068 5568
rect 3927 5528 4068 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 5350 5516 5356 5568
rect 5408 5556 5414 5568
rect 10502 5565 10508 5568
rect 5905 5559 5963 5565
rect 5905 5556 5917 5559
rect 5408 5528 5917 5556
rect 5408 5516 5414 5528
rect 5905 5525 5917 5528
rect 5951 5525 5963 5559
rect 5905 5519 5963 5525
rect 10486 5559 10508 5565
rect 10486 5525 10498 5559
rect 10486 5519 10508 5525
rect 10502 5516 10508 5519
rect 10560 5516 10566 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 10744 5528 11345 5556
rect 10744 5516 10750 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 17862 5516 17868 5568
rect 17920 5556 17926 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 17920 5528 18061 5556
rect 17920 5516 17926 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 22278 5516 22284 5568
rect 22336 5556 22342 5568
rect 23566 5556 23572 5568
rect 22336 5528 23572 5556
rect 22336 5516 22342 5528
rect 23566 5516 23572 5528
rect 23624 5516 23630 5568
rect 23750 5556 23756 5568
rect 23711 5528 23756 5556
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 25130 5556 25136 5568
rect 25091 5528 25136 5556
rect 25130 5516 25136 5528
rect 25188 5556 25194 5568
rect 25406 5556 25412 5568
rect 25188 5528 25412 5556
rect 25188 5516 25194 5528
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2038 5312 2044 5364
rect 2096 5352 2102 5364
rect 6270 5352 6276 5364
rect 2096 5324 6132 5352
rect 6231 5324 6276 5352
rect 2096 5312 2102 5324
rect 1949 5287 2007 5293
rect 1949 5253 1961 5287
rect 1995 5284 2007 5287
rect 2958 5284 2964 5296
rect 1995 5256 2964 5284
rect 1995 5253 2007 5256
rect 1949 5247 2007 5253
rect 2958 5244 2964 5256
rect 3016 5284 3022 5296
rect 3053 5287 3111 5293
rect 3053 5284 3065 5287
rect 3016 5256 3065 5284
rect 3016 5244 3022 5256
rect 3053 5253 3065 5256
rect 3099 5253 3111 5287
rect 3053 5247 3111 5253
rect 3694 5244 3700 5296
rect 3752 5284 3758 5296
rect 4433 5287 4491 5293
rect 3752 5256 4154 5284
rect 3752 5244 3758 5256
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 2038 5216 2044 5228
rect 1360 5188 2044 5216
rect 1360 5176 1366 5188
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 3970 5216 3976 5228
rect 3931 5188 3976 5216
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4126 5216 4154 5256
rect 4433 5253 4445 5287
rect 4479 5284 4491 5287
rect 4522 5284 4528 5296
rect 4479 5256 4528 5284
rect 4479 5253 4491 5256
rect 4433 5247 4491 5253
rect 4522 5244 4528 5256
rect 4580 5284 4586 5296
rect 5074 5284 5080 5296
rect 4580 5256 5080 5284
rect 4580 5244 4586 5256
rect 5074 5244 5080 5256
rect 5132 5244 5138 5296
rect 6104 5284 6132 5324
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 9674 5352 9680 5364
rect 9635 5324 9680 5352
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 9950 5352 9956 5364
rect 9911 5324 9956 5352
rect 9950 5312 9956 5324
rect 10008 5352 10014 5364
rect 10321 5355 10379 5361
rect 10321 5352 10333 5355
rect 10008 5324 10333 5352
rect 10008 5312 10014 5324
rect 10321 5321 10333 5324
rect 10367 5321 10379 5355
rect 10321 5315 10379 5321
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 10686 5361 10692 5364
rect 10643 5355 10692 5361
rect 10643 5352 10655 5355
rect 10560 5324 10655 5352
rect 10560 5312 10566 5324
rect 10643 5321 10655 5324
rect 10689 5321 10692 5355
rect 10643 5315 10692 5321
rect 10686 5312 10692 5315
rect 10744 5312 10750 5364
rect 11146 5352 11152 5364
rect 11107 5324 11152 5352
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 12161 5355 12219 5361
rect 12161 5321 12173 5355
rect 12207 5352 12219 5355
rect 12342 5352 12348 5364
rect 12207 5324 12348 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 7466 5284 7472 5296
rect 6104 5256 7472 5284
rect 7466 5244 7472 5256
rect 7524 5284 7530 5296
rect 9490 5284 9496 5296
rect 7524 5256 9496 5284
rect 7524 5244 7530 5256
rect 9490 5244 9496 5256
rect 9548 5244 9554 5296
rect 10781 5287 10839 5293
rect 10781 5253 10793 5287
rect 10827 5284 10839 5287
rect 11054 5284 11060 5296
rect 10827 5256 11060 5284
rect 10827 5253 10839 5256
rect 10781 5247 10839 5253
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 4893 5219 4951 5225
rect 4893 5216 4905 5219
rect 4126 5188 4905 5216
rect 4893 5185 4905 5188
rect 4939 5216 4951 5219
rect 5350 5216 5356 5228
rect 4939 5188 5356 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 6914 5216 6920 5228
rect 6871 5188 6920 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 9646 5188 10824 5216
rect 1820 5151 1878 5157
rect 1820 5117 1832 5151
rect 1866 5148 1878 5151
rect 2314 5148 2320 5160
rect 1866 5120 2320 5148
rect 1866 5117 1878 5120
rect 1820 5111 1878 5117
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3237 5151 3295 5157
rect 3237 5148 3249 5151
rect 3108 5120 3249 5148
rect 3108 5108 3114 5120
rect 3237 5117 3249 5120
rect 3283 5148 3295 5151
rect 3694 5148 3700 5160
rect 3283 5120 3700 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 3789 5151 3847 5157
rect 3789 5117 3801 5151
rect 3835 5148 3847 5151
rect 4706 5148 4712 5160
rect 3835 5120 4712 5148
rect 3835 5117 3847 5120
rect 3789 5111 3847 5117
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5080 1731 5083
rect 2406 5080 2412 5092
rect 1719 5052 2412 5080
rect 1719 5049 1731 5052
rect 1673 5043 1731 5049
rect 2406 5040 2412 5052
rect 2464 5040 2470 5092
rect 2774 5080 2780 5092
rect 2516 5052 2780 5080
rect 2317 5015 2375 5021
rect 2317 4981 2329 5015
rect 2363 5012 2375 5015
rect 2516 5012 2544 5052
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 3970 5040 3976 5092
rect 4028 5080 4034 5092
rect 4126 5080 4154 5120
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 8389 5151 8447 5157
rect 8389 5148 8401 5151
rect 6144 5120 8401 5148
rect 6144 5108 6150 5120
rect 8389 5117 8401 5120
rect 8435 5148 8447 5151
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 8435 5120 8585 5148
rect 8435 5117 8447 5120
rect 8389 5111 8447 5117
rect 8573 5117 8585 5120
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 4890 5080 4896 5092
rect 4028 5052 4154 5080
rect 4264 5052 4896 5080
rect 4028 5040 4034 5052
rect 2363 4984 2544 5012
rect 2685 5015 2743 5021
rect 2363 4981 2375 4984
rect 2317 4975 2375 4981
rect 2685 4981 2697 5015
rect 2731 5012 2743 5015
rect 2866 5012 2872 5024
rect 2731 4984 2872 5012
rect 2731 4981 2743 4984
rect 2685 4975 2743 4981
rect 2866 4972 2872 4984
rect 2924 4972 2930 5024
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 4264 5012 4292 5052
rect 4890 5040 4896 5052
rect 4948 5040 4954 5092
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5080 5043 5083
rect 5166 5080 5172 5092
rect 5031 5052 5172 5080
rect 5031 5049 5043 5052
rect 4985 5043 5043 5049
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 5537 5083 5595 5089
rect 5537 5049 5549 5083
rect 5583 5080 5595 5083
rect 5626 5080 5632 5092
rect 5583 5052 5632 5080
rect 5583 5049 5595 5052
rect 5537 5043 5595 5049
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 8588 5080 8616 5111
rect 8846 5108 8852 5160
rect 8904 5148 8910 5160
rect 9033 5151 9091 5157
rect 9033 5148 9045 5151
rect 8904 5120 9045 5148
rect 8904 5108 8910 5120
rect 9033 5117 9045 5120
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 9646 5080 9674 5188
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 10192 5120 10517 5148
rect 10192 5108 10198 5120
rect 10505 5117 10517 5120
rect 10551 5148 10563 5151
rect 10594 5148 10600 5160
rect 10551 5120 10600 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 10796 5148 10824 5188
rect 10870 5176 10876 5228
rect 10928 5216 10934 5228
rect 10928 5188 10973 5216
rect 10928 5176 10934 5188
rect 12176 5148 12204 5315
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12621 5355 12679 5361
rect 12621 5352 12633 5355
rect 12584 5324 12633 5352
rect 12584 5312 12590 5324
rect 12621 5321 12633 5324
rect 12667 5352 12679 5355
rect 13081 5355 13139 5361
rect 13081 5352 13093 5355
rect 12667 5324 13093 5352
rect 12667 5321 12679 5324
rect 12621 5315 12679 5321
rect 13081 5321 13093 5324
rect 13127 5352 13139 5355
rect 14642 5352 14648 5364
rect 13127 5324 14648 5352
rect 13127 5321 13139 5324
rect 13081 5315 13139 5321
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 14829 5355 14887 5361
rect 14829 5321 14841 5355
rect 14875 5352 14887 5355
rect 15746 5352 15752 5364
rect 14875 5324 15752 5352
rect 14875 5321 14887 5324
rect 14829 5315 14887 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 17218 5352 17224 5364
rect 17179 5324 17224 5352
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 18966 5312 18972 5364
rect 19024 5352 19030 5364
rect 19245 5355 19303 5361
rect 19245 5352 19257 5355
rect 19024 5324 19257 5352
rect 19024 5312 19030 5324
rect 19245 5321 19257 5324
rect 19291 5321 19303 5355
rect 19610 5352 19616 5364
rect 19571 5324 19616 5352
rect 19245 5315 19303 5321
rect 19610 5312 19616 5324
rect 19668 5312 19674 5364
rect 21082 5352 21088 5364
rect 21043 5324 21088 5352
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 22186 5312 22192 5364
rect 22244 5352 22250 5364
rect 22465 5355 22523 5361
rect 22465 5352 22477 5355
rect 22244 5324 22477 5352
rect 22244 5312 22250 5324
rect 22465 5321 22477 5324
rect 22511 5321 22523 5355
rect 22465 5315 22523 5321
rect 12802 5244 12808 5296
rect 12860 5284 12866 5296
rect 18138 5284 18144 5296
rect 12860 5256 18144 5284
rect 12860 5244 12866 5256
rect 18138 5244 18144 5256
rect 18196 5284 18202 5296
rect 20257 5287 20315 5293
rect 18196 5256 18368 5284
rect 18196 5244 18202 5256
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5216 13967 5219
rect 14734 5216 14740 5228
rect 13955 5188 14740 5216
rect 13955 5185 13967 5188
rect 13909 5179 13967 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 18340 5225 18368 5256
rect 20257 5253 20269 5287
rect 20303 5284 20315 5287
rect 22370 5284 22376 5296
rect 20303 5256 22376 5284
rect 20303 5253 20315 5256
rect 20257 5247 20315 5253
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 22480 5284 22508 5315
rect 22646 5312 22652 5364
rect 22704 5352 22710 5364
rect 22741 5355 22799 5361
rect 22741 5352 22753 5355
rect 22704 5324 22753 5352
rect 22704 5312 22710 5324
rect 22741 5321 22753 5324
rect 22787 5321 22799 5355
rect 23382 5352 23388 5364
rect 23343 5324 23388 5352
rect 22741 5315 22799 5321
rect 23382 5312 23388 5324
rect 23440 5312 23446 5364
rect 24118 5312 24124 5364
rect 24176 5352 24182 5364
rect 24673 5355 24731 5361
rect 24673 5352 24685 5355
rect 24176 5324 24685 5352
rect 24176 5312 24182 5324
rect 24673 5321 24685 5324
rect 24719 5321 24731 5355
rect 24673 5315 24731 5321
rect 24762 5284 24768 5296
rect 22480 5256 24768 5284
rect 24762 5244 24768 5256
rect 24820 5244 24826 5296
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 15528 5188 15669 5216
rect 15528 5176 15534 5188
rect 15657 5185 15669 5188
rect 15703 5216 15715 5219
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 15703 5188 16865 5216
rect 15703 5185 15715 5188
rect 15657 5179 15715 5185
rect 16853 5185 16865 5188
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5185 18383 5219
rect 18325 5179 18383 5185
rect 19242 5176 19248 5228
rect 19300 5216 19306 5228
rect 20625 5219 20683 5225
rect 20625 5216 20637 5219
rect 19300 5188 20637 5216
rect 19300 5176 19306 5188
rect 20088 5157 20116 5188
rect 20625 5185 20637 5188
rect 20671 5185 20683 5219
rect 20625 5179 20683 5185
rect 10796 5120 12204 5148
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 12943 5120 13492 5148
rect 20051 5120 20085 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 8588 5052 9674 5080
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 11514 5080 11520 5092
rect 10744 5052 11520 5080
rect 10744 5040 10750 5052
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 3016 4984 4292 5012
rect 5184 5012 5212 5040
rect 13464 5024 13492 5120
rect 20073 5117 20085 5120
rect 20119 5117 20131 5151
rect 20073 5111 20131 5117
rect 21177 5151 21235 5157
rect 21177 5117 21189 5151
rect 21223 5148 21235 5151
rect 22738 5148 22744 5160
rect 21223 5120 22744 5148
rect 21223 5117 21235 5120
rect 21177 5111 21235 5117
rect 22738 5108 22744 5120
rect 22796 5108 22802 5160
rect 23382 5108 23388 5160
rect 23440 5148 23446 5160
rect 23661 5151 23719 5157
rect 23661 5148 23673 5151
rect 23440 5120 23673 5148
rect 23440 5108 23446 5120
rect 23661 5117 23673 5120
rect 23707 5117 23719 5151
rect 23661 5111 23719 5117
rect 23750 5108 23756 5160
rect 23808 5148 23814 5160
rect 24118 5148 24124 5160
rect 23808 5120 24124 5148
rect 23808 5108 23814 5120
rect 24118 5108 24124 5120
rect 24176 5108 24182 5160
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 25222 5108 25228 5120
rect 25280 5148 25286 5160
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25280 5120 25789 5148
rect 25280 5108 25286 5120
rect 25777 5117 25789 5120
rect 25823 5117 25835 5151
rect 25777 5111 25835 5117
rect 14271 5083 14329 5089
rect 14271 5049 14283 5083
rect 14317 5049 14329 5083
rect 14271 5043 14329 5049
rect 15978 5083 16036 5089
rect 15978 5049 15990 5083
rect 16024 5049 16036 5083
rect 15978 5043 16036 5049
rect 18417 5083 18475 5089
rect 18417 5049 18429 5083
rect 18463 5049 18475 5083
rect 18417 5043 18475 5049
rect 18969 5083 19027 5089
rect 18969 5049 18981 5083
rect 19015 5080 19027 5083
rect 19058 5080 19064 5092
rect 19015 5052 19064 5080
rect 19015 5049 19027 5052
rect 18969 5043 19027 5049
rect 5813 5015 5871 5021
rect 5813 5012 5825 5015
rect 5184 4984 5825 5012
rect 3016 4972 3022 4984
rect 5813 4981 5825 4984
rect 5859 4981 5871 5015
rect 5813 4975 5871 4981
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 7190 5012 7196 5024
rect 6687 4984 7196 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7742 5012 7748 5024
rect 7703 4984 7748 5012
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 8018 5012 8024 5024
rect 7979 4984 8024 5012
rect 8018 4972 8024 4984
rect 8076 4972 8082 5024
rect 8662 5012 8668 5024
rect 8623 4984 8668 5012
rect 8662 4972 8668 4984
rect 8720 4972 8726 5024
rect 13446 5012 13452 5024
rect 13407 4984 13452 5012
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 13817 5015 13875 5021
rect 13817 4981 13829 5015
rect 13863 5012 13875 5015
rect 14286 5012 14314 5043
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 13863 4984 15301 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 15289 4981 15301 4984
rect 15335 5012 15347 5015
rect 15654 5012 15660 5024
rect 15335 4984 15660 5012
rect 15335 4981 15347 4984
rect 15289 4975 15347 4981
rect 15654 4972 15660 4984
rect 15712 5012 15718 5024
rect 15993 5012 16021 5043
rect 16574 5012 16580 5024
rect 15712 4984 16021 5012
rect 16535 4984 16580 5012
rect 15712 4972 15718 4984
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 5012 17834 5024
rect 18432 5012 18460 5043
rect 19058 5040 19064 5052
rect 19116 5040 19122 5092
rect 21082 5040 21088 5092
rect 21140 5080 21146 5092
rect 21498 5083 21556 5089
rect 21498 5080 21510 5083
rect 21140 5052 21510 5080
rect 21140 5040 21146 5052
rect 21498 5049 21510 5052
rect 21544 5049 21556 5083
rect 21498 5043 21556 5049
rect 22094 5012 22100 5024
rect 17828 4984 18460 5012
rect 22055 4984 22100 5012
rect 17828 4972 17834 4984
rect 22094 4972 22100 4984
rect 22152 4972 22158 5024
rect 23566 4972 23572 5024
rect 23624 5012 23630 5024
rect 23753 5015 23811 5021
rect 23753 5012 23765 5015
rect 23624 4984 23765 5012
rect 23624 4972 23630 4984
rect 23753 4981 23765 4984
rect 23799 4981 23811 5015
rect 25406 5012 25412 5024
rect 25367 4984 25412 5012
rect 23753 4975 23811 4981
rect 25406 4972 25412 4984
rect 25464 4972 25470 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1535 4811 1593 4817
rect 1535 4777 1547 4811
rect 1581 4808 1593 4811
rect 2222 4808 2228 4820
rect 1581 4780 2228 4808
rect 1581 4777 1593 4780
rect 1535 4771 1593 4777
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 2958 4808 2964 4820
rect 2363 4780 2964 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 3602 4808 3608 4820
rect 3559 4780 3608 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 3602 4768 3608 4780
rect 3660 4768 3666 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3752 4780 3801 4808
rect 3752 4768 3758 4780
rect 3789 4777 3801 4780
rect 3835 4808 3847 4811
rect 3878 4808 3884 4820
rect 3835 4780 3884 4808
rect 3835 4777 3847 4780
rect 3789 4771 3847 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4080 4780 4261 4808
rect 4080 4752 4108 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4706 4808 4712 4820
rect 4667 4780 4712 4808
rect 4249 4771 4307 4777
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 6454 4808 6460 4820
rect 6415 4780 6460 4808
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 6917 4811 6975 4817
rect 6917 4777 6929 4811
rect 6963 4808 6975 4811
rect 7190 4808 7196 4820
rect 6963 4780 7196 4808
rect 6963 4777 6975 4780
rect 6917 4771 6975 4777
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 7300 4780 8217 4808
rect 1670 4700 1676 4752
rect 1728 4740 1734 4752
rect 1857 4743 1915 4749
rect 1857 4740 1869 4743
rect 1728 4712 1869 4740
rect 1728 4700 1734 4712
rect 1857 4709 1869 4712
rect 1903 4709 1915 4743
rect 1857 4703 1915 4709
rect 3145 4743 3203 4749
rect 3145 4709 3157 4743
rect 3191 4740 3203 4743
rect 3234 4740 3240 4752
rect 3191 4712 3240 4740
rect 3191 4709 3203 4712
rect 3145 4703 3203 4709
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 4062 4700 4068 4752
rect 4120 4700 4126 4752
rect 5074 4740 5080 4752
rect 5035 4712 5080 4740
rect 5074 4700 5080 4712
rect 5132 4700 5138 4752
rect 5626 4740 5632 4752
rect 5587 4712 5632 4740
rect 5626 4700 5632 4712
rect 5684 4740 5690 4752
rect 7098 4740 7104 4752
rect 5684 4712 7104 4740
rect 5684 4700 5690 4712
rect 7098 4700 7104 4712
rect 7156 4740 7162 4752
rect 7300 4749 7328 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8205 4771 8263 4777
rect 8665 4811 8723 4817
rect 8665 4777 8677 4811
rect 8711 4808 8723 4811
rect 8846 4808 8852 4820
rect 8711 4780 8852 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 8938 4768 8944 4820
rect 8996 4808 9002 4820
rect 10321 4811 10379 4817
rect 10321 4808 10333 4811
rect 8996 4780 10333 4808
rect 8996 4768 9002 4780
rect 10321 4777 10333 4780
rect 10367 4777 10379 4811
rect 10686 4808 10692 4820
rect 10647 4780 10692 4808
rect 10321 4771 10379 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11330 4808 11336 4820
rect 11291 4780 11336 4808
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14461 4811 14519 4817
rect 14461 4808 14473 4811
rect 13872 4780 14473 4808
rect 13872 4768 13878 4780
rect 14461 4777 14473 4780
rect 14507 4777 14519 4811
rect 14461 4771 14519 4777
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15013 4811 15071 4817
rect 15013 4808 15025 4811
rect 14884 4780 15025 4808
rect 14884 4768 14890 4780
rect 15013 4777 15025 4780
rect 15059 4777 15071 4811
rect 17037 4811 17095 4817
rect 17037 4808 17049 4811
rect 15013 4771 15071 4777
rect 15672 4780 17049 4808
rect 7285 4743 7343 4749
rect 7285 4740 7297 4743
rect 7156 4712 7297 4740
rect 7156 4700 7162 4712
rect 7285 4709 7297 4712
rect 7331 4709 7343 4743
rect 7285 4703 7343 4709
rect 7377 4743 7435 4749
rect 7377 4709 7389 4743
rect 7423 4740 7435 4743
rect 7742 4740 7748 4752
rect 7423 4712 7748 4740
rect 7423 4709 7435 4712
rect 7377 4703 7435 4709
rect 7742 4700 7748 4712
rect 7800 4700 7806 4752
rect 9030 4740 9036 4752
rect 8991 4712 9036 4740
rect 9030 4700 9036 4712
rect 9088 4740 9094 4752
rect 9677 4743 9735 4749
rect 9677 4740 9689 4743
rect 9088 4712 9689 4740
rect 9088 4700 9094 4712
rect 9677 4709 9689 4712
rect 9723 4740 9735 4743
rect 10962 4740 10968 4752
rect 9723 4712 10968 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 13630 4740 13636 4752
rect 11480 4712 11836 4740
rect 13591 4712 13636 4740
rect 11480 4700 11486 4712
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 2222 4672 2228 4684
rect 1510 4644 2228 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 2222 4632 2228 4644
rect 2280 4632 2286 4684
rect 2406 4632 2412 4684
rect 2464 4672 2470 4684
rect 3326 4672 3332 4684
rect 2464 4644 3332 4672
rect 2464 4632 2470 4644
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 11517 4675 11575 4681
rect 9916 4644 10088 4672
rect 9916 4632 9922 4644
rect 2038 4564 2044 4616
rect 2096 4604 2102 4616
rect 2774 4604 2780 4616
rect 2096 4576 2780 4604
rect 2096 4564 2102 4576
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 4982 4604 4988 4616
rect 4943 4576 4988 4604
rect 4982 4564 4988 4576
rect 5040 4604 5046 4616
rect 5905 4607 5963 4613
rect 5905 4604 5917 4607
rect 5040 4576 5917 4604
rect 5040 4564 5046 4576
rect 5905 4573 5917 4576
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 7561 4607 7619 4613
rect 7561 4573 7573 4607
rect 7607 4604 7619 4607
rect 8018 4604 8024 4616
rect 7607 4576 8024 4604
rect 7607 4573 7619 4576
rect 7561 4567 7619 4573
rect 2682 4536 2688 4548
rect 2643 4508 2688 4536
rect 2682 4496 2688 4508
rect 2740 4496 2746 4548
rect 4706 4496 4712 4548
rect 4764 4536 4770 4548
rect 7576 4536 7604 4567
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 10060 4613 10088 4644
rect 11517 4641 11529 4675
rect 11563 4672 11575 4675
rect 11606 4672 11612 4684
rect 11563 4644 11612 4672
rect 11563 4641 11575 4644
rect 11517 4635 11575 4641
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 11808 4681 11836 4712
rect 13630 4700 13636 4712
rect 13688 4700 13694 4752
rect 14185 4743 14243 4749
rect 14185 4709 14197 4743
rect 14231 4740 14243 4743
rect 14366 4740 14372 4752
rect 14231 4712 14372 4740
rect 14231 4709 14243 4712
rect 14185 4703 14243 4709
rect 14366 4700 14372 4712
rect 14424 4740 14430 4752
rect 15672 4740 15700 4780
rect 17037 4777 17049 4780
rect 17083 4808 17095 4811
rect 17126 4808 17132 4820
rect 17083 4780 17132 4808
rect 17083 4777 17095 4780
rect 17037 4771 17095 4777
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 18138 4808 18144 4820
rect 18099 4780 18144 4808
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18322 4768 18328 4820
rect 18380 4808 18386 4820
rect 19245 4811 19303 4817
rect 19245 4808 19257 4811
rect 18380 4780 19257 4808
rect 18380 4768 18386 4780
rect 19245 4777 19257 4780
rect 19291 4777 19303 4811
rect 19245 4771 19303 4777
rect 20625 4811 20683 4817
rect 20625 4777 20637 4811
rect 20671 4808 20683 4811
rect 21266 4808 21272 4820
rect 20671 4780 21272 4808
rect 20671 4777 20683 4780
rect 20625 4771 20683 4777
rect 21266 4768 21272 4780
rect 21324 4808 21330 4820
rect 21324 4780 21541 4808
rect 21324 4768 21330 4780
rect 14424 4712 15700 4740
rect 14424 4700 14430 4712
rect 16114 4700 16120 4752
rect 16172 4740 16178 4752
rect 16209 4743 16267 4749
rect 16209 4740 16221 4743
rect 16172 4712 16221 4740
rect 16172 4700 16178 4712
rect 16209 4709 16221 4712
rect 16255 4740 16267 4743
rect 16574 4740 16580 4752
rect 16255 4712 16580 4740
rect 16255 4709 16267 4712
rect 16209 4703 16267 4709
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 16761 4743 16819 4749
rect 16761 4709 16773 4743
rect 16807 4740 16819 4743
rect 17678 4740 17684 4752
rect 16807 4712 17684 4740
rect 16807 4709 16819 4712
rect 16761 4703 16819 4709
rect 17678 4700 17684 4712
rect 17736 4700 17742 4752
rect 17770 4700 17776 4752
rect 17828 4740 17834 4752
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 17828 4712 18429 4740
rect 17828 4700 17834 4712
rect 18417 4709 18429 4712
rect 18463 4709 18475 4743
rect 18417 4703 18475 4709
rect 20714 4700 20720 4752
rect 20772 4740 20778 4752
rect 21082 4740 21088 4752
rect 20772 4712 21088 4740
rect 20772 4700 20778 4712
rect 21082 4700 21088 4712
rect 21140 4740 21146 4752
rect 21406 4743 21464 4749
rect 21406 4740 21418 4743
rect 21140 4712 21418 4740
rect 21140 4700 21146 4712
rect 21406 4709 21418 4712
rect 21452 4709 21464 4743
rect 21406 4703 21464 4709
rect 11793 4675 11851 4681
rect 11793 4641 11805 4675
rect 11839 4672 11851 4675
rect 12158 4672 12164 4684
rect 11839 4644 12164 4672
rect 11839 4641 11851 4644
rect 11793 4635 11851 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 19702 4632 19708 4684
rect 19760 4672 19766 4684
rect 19864 4675 19922 4681
rect 19864 4672 19876 4675
rect 19760 4644 19876 4672
rect 19760 4632 19766 4644
rect 19864 4641 19876 4644
rect 19910 4672 19922 4675
rect 20990 4672 20996 4684
rect 19910 4644 20996 4672
rect 19910 4641 19922 4644
rect 19864 4635 19922 4641
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 21513 4672 21541 4780
rect 22462 4768 22468 4820
rect 22520 4808 22526 4820
rect 22557 4811 22615 4817
rect 22557 4808 22569 4811
rect 22520 4780 22569 4808
rect 22520 4768 22526 4780
rect 22557 4777 22569 4780
rect 22603 4777 22615 4811
rect 22557 4771 22615 4777
rect 22738 4768 22744 4820
rect 22796 4808 22802 4820
rect 24489 4811 24547 4817
rect 24489 4808 24501 4811
rect 22796 4780 24501 4808
rect 22796 4768 22802 4780
rect 24489 4777 24501 4780
rect 24535 4777 24547 4811
rect 24489 4771 24547 4777
rect 22094 4700 22100 4752
rect 22152 4740 22158 4752
rect 22646 4740 22652 4752
rect 22152 4712 22652 4740
rect 22152 4700 22158 4712
rect 22646 4700 22652 4712
rect 22704 4740 22710 4752
rect 23017 4743 23075 4749
rect 23017 4740 23029 4743
rect 22704 4712 23029 4740
rect 22704 4700 22710 4712
rect 23017 4709 23029 4712
rect 23063 4709 23075 4743
rect 23017 4703 23075 4709
rect 23569 4743 23627 4749
rect 23569 4709 23581 4743
rect 23615 4740 23627 4743
rect 23934 4740 23940 4752
rect 23615 4712 23940 4740
rect 23615 4709 23627 4712
rect 23569 4703 23627 4709
rect 23934 4700 23940 4712
rect 23992 4700 23998 4752
rect 24118 4740 24124 4752
rect 24079 4712 24124 4740
rect 24118 4700 24124 4712
rect 24176 4740 24182 4752
rect 24176 4712 24900 4740
rect 24176 4700 24182 4712
rect 22554 4672 22560 4684
rect 21513 4644 22560 4672
rect 22554 4632 22560 4644
rect 22612 4632 22618 4684
rect 23842 4632 23848 4684
rect 23900 4672 23906 4684
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 23900 4644 24409 4672
rect 23900 4632 23906 4644
rect 24397 4641 24409 4644
rect 24443 4672 24455 4675
rect 24670 4672 24676 4684
rect 24443 4644 24676 4672
rect 24443 4641 24455 4644
rect 24397 4635 24455 4641
rect 24670 4632 24676 4644
rect 24728 4632 24734 4684
rect 24872 4681 24900 4712
rect 24857 4675 24915 4681
rect 24857 4641 24869 4675
rect 24903 4641 24915 4675
rect 24857 4635 24915 4641
rect 10045 4607 10103 4613
rect 9824 4576 9996 4604
rect 9824 4564 9830 4576
rect 9968 4545 9996 4576
rect 10045 4573 10057 4607
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4604 16175 4607
rect 16206 4604 16212 4616
rect 16163 4576 16212 4604
rect 16163 4573 16175 4576
rect 16117 4567 16175 4573
rect 4764 4508 7604 4536
rect 9953 4539 10011 4545
rect 4764 4496 4770 4508
rect 9953 4505 9965 4539
rect 9999 4505 10011 4539
rect 9953 4499 10011 4505
rect 2498 4428 2504 4480
rect 2556 4477 2562 4480
rect 2556 4471 2605 4477
rect 2556 4437 2559 4471
rect 2593 4437 2605 4471
rect 2556 4431 2605 4437
rect 2556 4428 2562 4431
rect 9306 4428 9312 4480
rect 9364 4468 9370 4480
rect 9401 4471 9459 4477
rect 9401 4468 9413 4471
rect 9364 4440 9413 4468
rect 9364 4428 9370 4440
rect 9401 4437 9413 4440
rect 9447 4437 9459 4471
rect 9401 4431 9459 4437
rect 9842 4471 9900 4477
rect 9842 4437 9854 4471
rect 9888 4468 9900 4471
rect 10778 4468 10784 4480
rect 9888 4440 10784 4468
rect 9888 4437 9900 4440
rect 9842 4431 9900 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 12250 4468 12256 4480
rect 12211 4440 12256 4468
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 13262 4468 13268 4480
rect 13223 4440 13268 4468
rect 13262 4428 13268 4440
rect 13320 4468 13326 4480
rect 13556 4468 13584 4567
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 18322 4604 18328 4616
rect 18283 4576 18328 4604
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 18966 4604 18972 4616
rect 18927 4576 18972 4604
rect 18966 4564 18972 4576
rect 19024 4564 19030 4616
rect 21082 4604 21088 4616
rect 21043 4576 21088 4604
rect 21082 4564 21088 4576
rect 21140 4564 21146 4616
rect 22922 4604 22928 4616
rect 22883 4576 22928 4604
rect 22922 4564 22928 4576
rect 22980 4564 22986 4616
rect 18230 4496 18236 4548
rect 18288 4536 18294 4548
rect 19935 4539 19993 4545
rect 19935 4536 19947 4539
rect 18288 4508 19947 4536
rect 18288 4496 18294 4508
rect 19935 4505 19947 4508
rect 19981 4505 19993 4539
rect 19935 4499 19993 4505
rect 20346 4496 20352 4548
rect 20404 4536 20410 4548
rect 20404 4508 23474 4536
rect 20404 4496 20410 4508
rect 15654 4468 15660 4480
rect 13320 4440 13584 4468
rect 15615 4440 15660 4468
rect 13320 4428 13326 4440
rect 15654 4428 15660 4440
rect 15712 4428 15718 4480
rect 17494 4468 17500 4480
rect 17407 4440 17500 4468
rect 17494 4428 17500 4440
rect 17552 4468 17558 4480
rect 20070 4468 20076 4480
rect 17552 4440 20076 4468
rect 17552 4428 17558 4440
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 22002 4468 22008 4480
rect 21963 4440 22008 4468
rect 22002 4428 22008 4440
rect 22060 4428 22066 4480
rect 23446 4468 23474 4508
rect 25130 4468 25136 4480
rect 23446 4440 25136 4468
rect 25130 4428 25136 4440
rect 25188 4428 25194 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2424 4236 7696 4264
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 2424 4128 2452 4236
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 2961 4199 3019 4205
rect 2961 4196 2973 4199
rect 2832 4168 2973 4196
rect 2832 4156 2838 4168
rect 2961 4165 2973 4168
rect 3007 4196 3019 4199
rect 3007 4168 5396 4196
rect 3007 4165 3019 4168
rect 2961 4159 3019 4165
rect 1811 4100 2452 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4029 1915 4063
rect 1857 4023 1915 4029
rect 1872 3924 1900 4023
rect 1946 4020 1952 4072
rect 2004 4060 2010 4072
rect 2424 4069 2452 4100
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 5077 4131 5135 4137
rect 5077 4128 5089 4131
rect 4856 4100 5089 4128
rect 4856 4088 4862 4100
rect 5077 4097 5089 4100
rect 5123 4097 5135 4131
rect 5368 4128 5396 4168
rect 5534 4156 5540 4208
rect 5592 4196 5598 4208
rect 5629 4199 5687 4205
rect 5629 4196 5641 4199
rect 5592 4168 5641 4196
rect 5592 4156 5598 4168
rect 5629 4165 5641 4168
rect 5675 4165 5687 4199
rect 5629 4159 5687 4165
rect 5994 4128 6000 4140
rect 5368 4100 6000 4128
rect 5077 4091 5135 4097
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6512 4100 6929 4128
rect 6512 4088 6518 4100
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 2225 4063 2283 4069
rect 2225 4060 2237 4063
rect 2004 4032 2237 4060
rect 2004 4020 2010 4032
rect 2225 4029 2237 4032
rect 2271 4029 2283 4063
rect 2225 4023 2283 4029
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4029 2467 4063
rect 3694 4060 3700 4072
rect 3655 4032 3700 4060
rect 2409 4023 2467 4029
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 3970 4060 3976 4072
rect 3931 4032 3976 4060
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 7668 4060 7696 4236
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 7837 4267 7895 4273
rect 7837 4264 7849 4267
rect 7800 4236 7849 4264
rect 7800 4224 7806 4236
rect 7837 4233 7849 4236
rect 7883 4233 7895 4267
rect 9582 4264 9588 4276
rect 9543 4236 9588 4264
rect 7837 4227 7895 4233
rect 9582 4224 9588 4236
rect 9640 4224 9646 4276
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 10134 4264 10140 4276
rect 10091 4236 10140 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 10134 4224 10140 4236
rect 10192 4264 10198 4276
rect 10594 4264 10600 4276
rect 10192 4236 10600 4264
rect 10192 4224 10198 4236
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11606 4264 11612 4276
rect 11287 4236 11612 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 12158 4264 12164 4276
rect 12119 4236 12164 4264
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 12621 4267 12679 4273
rect 12621 4233 12633 4267
rect 12667 4264 12679 4267
rect 15930 4264 15936 4276
rect 12667 4236 15936 4264
rect 12667 4233 12679 4236
rect 12621 4227 12679 4233
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 16114 4264 16120 4276
rect 16075 4236 16120 4264
rect 16114 4224 16120 4236
rect 16172 4224 16178 4276
rect 17497 4267 17555 4273
rect 17497 4233 17509 4267
rect 17543 4264 17555 4267
rect 17770 4264 17776 4276
rect 17543 4236 17776 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 17770 4224 17776 4236
rect 17828 4264 17834 4276
rect 18969 4267 19027 4273
rect 18969 4264 18981 4267
rect 17828 4236 18981 4264
rect 17828 4224 17834 4236
rect 18969 4233 18981 4236
rect 19015 4233 19027 4267
rect 18969 4227 19027 4233
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19426 4264 19432 4276
rect 19383 4236 19432 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 21821 4267 21879 4273
rect 19536 4236 20576 4264
rect 9858 4156 9864 4208
rect 9916 4205 9922 4208
rect 9916 4199 9965 4205
rect 9916 4165 9919 4199
rect 9953 4165 9965 4199
rect 11514 4196 11520 4208
rect 9916 4159 9965 4165
rect 10152 4168 11520 4196
rect 9916 4156 9922 4159
rect 10152 4140 10180 4168
rect 11514 4156 11520 4168
rect 11572 4156 11578 4208
rect 14366 4156 14372 4208
rect 14424 4196 14430 4208
rect 14553 4199 14611 4205
rect 14553 4196 14565 4199
rect 14424 4168 14565 4196
rect 14424 4156 14430 4168
rect 14553 4165 14565 4168
rect 14599 4196 14611 4199
rect 15749 4199 15807 4205
rect 15749 4196 15761 4199
rect 14599 4168 15761 4196
rect 14599 4165 14611 4168
rect 14553 4159 14611 4165
rect 15749 4165 15761 4168
rect 15795 4196 15807 4199
rect 16206 4196 16212 4208
rect 15795 4168 16212 4196
rect 15795 4165 15807 4168
rect 15749 4159 15807 4165
rect 16206 4156 16212 4168
rect 16264 4156 16270 4208
rect 17037 4199 17095 4205
rect 17037 4165 17049 4199
rect 17083 4196 17095 4199
rect 19058 4196 19064 4208
rect 17083 4168 19064 4196
rect 17083 4165 17095 4168
rect 17037 4159 17095 4165
rect 19058 4156 19064 4168
rect 19116 4156 19122 4208
rect 19536 4196 19564 4236
rect 19702 4196 19708 4208
rect 19306 4168 19564 4196
rect 19663 4168 19708 4196
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 10134 4128 10140 4140
rect 7892 4100 9674 4128
rect 10047 4100 10140 4128
rect 7892 4088 7898 4100
rect 8110 4060 8116 4072
rect 7668 4032 8116 4060
rect 8110 4020 8116 4032
rect 8168 4060 8174 4072
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 8168 4032 8585 4060
rect 8168 4020 8174 4032
rect 8573 4029 8585 4032
rect 8619 4060 8631 4063
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 8619 4032 9229 4060
rect 8619 4029 8631 4032
rect 8573 4023 8631 4029
rect 9217 4029 9229 4032
rect 9263 4060 9275 4063
rect 9306 4060 9312 4072
rect 9263 4032 9312 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 9646 4060 9674 4100
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4128 14059 4131
rect 16485 4131 16543 4137
rect 14047 4100 15424 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 9646 4032 10517 4060
rect 10505 4029 10517 4032
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 11333 4063 11391 4069
rect 11333 4060 11345 4063
rect 11204 4032 11345 4060
rect 11204 4020 11210 4032
rect 11333 4029 11345 4032
rect 11379 4060 11391 4063
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11379 4032 11805 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11793 4029 11805 4032
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 12483 4032 13032 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 3326 3992 3332 4004
rect 3287 3964 3332 3992
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 4154 3952 4160 4004
rect 4212 3992 4218 4004
rect 4893 3995 4951 4001
rect 4212 3964 4257 3992
rect 4212 3952 4218 3964
rect 4893 3961 4905 3995
rect 4939 3992 4951 3995
rect 5166 3992 5172 4004
rect 4939 3964 5172 3992
rect 4939 3961 4951 3964
rect 4893 3955 4951 3961
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 6641 3995 6699 4001
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 7006 3992 7012 4004
rect 6687 3964 7012 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 7561 3995 7619 4001
rect 7561 3992 7573 3995
rect 7156 3964 7573 3992
rect 7156 3952 7162 3964
rect 7561 3961 7573 3964
rect 7607 3992 7619 3995
rect 7650 3992 7656 4004
rect 7607 3964 7656 3992
rect 7607 3961 7619 3964
rect 7561 3955 7619 3961
rect 7650 3952 7656 3964
rect 7708 3952 7714 4004
rect 8389 3995 8447 4001
rect 8389 3961 8401 3995
rect 8435 3961 8447 3995
rect 8938 3992 8944 4004
rect 8899 3964 8944 3992
rect 8389 3955 8447 3961
rect 2130 3924 2136 3936
rect 1872 3896 2136 3924
rect 2130 3884 2136 3896
rect 2188 3924 2194 3936
rect 4525 3927 4583 3933
rect 4525 3924 4537 3927
rect 2188 3896 4537 3924
rect 2188 3884 2194 3896
rect 4525 3893 4537 3896
rect 4571 3924 4583 3927
rect 4982 3924 4988 3936
rect 4571 3896 4988 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 5997 3927 6055 3933
rect 5997 3924 6009 3927
rect 5132 3896 6009 3924
rect 5132 3884 5138 3896
rect 5997 3893 6009 3896
rect 6043 3893 6055 3927
rect 8294 3924 8300 3936
rect 8255 3896 8300 3924
rect 5997 3887 6055 3893
rect 8294 3884 8300 3896
rect 8352 3924 8358 3936
rect 8404 3924 8432 3955
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 9490 3952 9496 4004
rect 9548 3992 9554 4004
rect 9769 3995 9827 4001
rect 9769 3992 9781 3995
rect 9548 3964 9781 3992
rect 9548 3952 9554 3964
rect 9769 3961 9781 3964
rect 9815 3961 9827 3995
rect 9769 3955 9827 3961
rect 13004 3936 13032 4032
rect 14093 3995 14151 4001
rect 14093 3961 14105 3995
rect 14139 3992 14151 3995
rect 14921 3995 14979 4001
rect 14921 3992 14933 3995
rect 14139 3964 14933 3992
rect 14139 3961 14151 3964
rect 14093 3955 14151 3961
rect 14921 3961 14933 3964
rect 14967 3961 14979 3995
rect 14921 3955 14979 3961
rect 10778 3924 10784 3936
rect 8352 3896 8432 3924
rect 10739 3896 10784 3924
rect 8352 3884 8358 3896
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 12986 3924 12992 3936
rect 12947 3896 12992 3924
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13541 3927 13599 3933
rect 13541 3893 13553 3927
rect 13587 3924 13599 3927
rect 13630 3924 13636 3936
rect 13587 3896 13636 3924
rect 13587 3893 13599 3896
rect 13541 3887 13599 3893
rect 13630 3884 13636 3896
rect 13688 3924 13694 3936
rect 14108 3924 14136 3955
rect 15396 3933 15424 4100
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 17494 4128 17500 4140
rect 16531 4100 17500 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 17494 4088 17500 4100
rect 17552 4088 17558 4140
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 19076 4128 19104 4156
rect 19306 4128 19334 4168
rect 19702 4156 19708 4168
rect 19760 4156 19766 4208
rect 17920 4100 18276 4128
rect 19076 4100 19334 4128
rect 17920 4088 17926 4100
rect 17954 4060 17960 4072
rect 17880 4032 17960 4060
rect 16574 3992 16580 4004
rect 16535 3964 16580 3992
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 17880 3992 17908 4032
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18138 4060 18144 4072
rect 18095 4032 18144 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 16684 3964 17908 3992
rect 18248 3992 18276 4100
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 20070 4128 20076 4140
rect 19484 4100 20076 4128
rect 19484 4088 19490 4100
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20548 4137 20576 4236
rect 21821 4233 21833 4267
rect 21867 4264 21879 4267
rect 22002 4264 22008 4276
rect 21867 4236 22008 4264
rect 21867 4233 21879 4236
rect 21821 4227 21879 4233
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 24670 4264 24676 4276
rect 24631 4236 24676 4264
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 22557 4199 22615 4205
rect 22557 4165 22569 4199
rect 22603 4196 22615 4199
rect 23934 4196 23940 4208
rect 22603 4168 23940 4196
rect 22603 4165 22615 4168
rect 22557 4159 22615 4165
rect 23934 4156 23940 4168
rect 23992 4156 23998 4208
rect 24854 4156 24860 4208
rect 24912 4196 24918 4208
rect 25409 4199 25467 4205
rect 25409 4196 25421 4199
rect 24912 4168 25421 4196
rect 24912 4156 24918 4168
rect 25409 4165 25421 4168
rect 25455 4165 25467 4199
rect 25409 4159 25467 4165
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4128 20591 4131
rect 22462 4128 22468 4140
rect 20579 4100 22468 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 22462 4088 22468 4100
rect 22520 4128 22526 4140
rect 22922 4128 22928 4140
rect 22520 4100 22928 4128
rect 22520 4088 22526 4100
rect 22922 4088 22928 4100
rect 22980 4088 22986 4140
rect 25774 4128 25780 4140
rect 25240 4100 25780 4128
rect 23198 4020 23204 4072
rect 23256 4060 23262 4072
rect 23477 4063 23535 4069
rect 23477 4060 23489 4063
rect 23256 4032 23489 4060
rect 23256 4020 23262 4032
rect 23477 4029 23489 4032
rect 23523 4060 23535 4063
rect 23661 4063 23719 4069
rect 23661 4060 23673 4063
rect 23523 4032 23673 4060
rect 23523 4029 23535 4032
rect 23477 4023 23535 4029
rect 23661 4029 23673 4032
rect 23707 4029 23719 4063
rect 23661 4023 23719 4029
rect 24118 4020 24124 4072
rect 24176 4060 24182 4072
rect 25240 4069 25268 4100
rect 25774 4088 25780 4100
rect 25832 4088 25838 4140
rect 24213 4063 24271 4069
rect 24213 4060 24225 4063
rect 24176 4032 24225 4060
rect 24176 4020 24182 4032
rect 24213 4029 24225 4032
rect 24259 4060 24271 4063
rect 25225 4063 25283 4069
rect 24259 4032 25176 4060
rect 24259 4029 24271 4032
rect 24213 4023 24271 4029
rect 18370 3995 18428 4001
rect 18370 3992 18382 3995
rect 18248 3964 18382 3992
rect 13688 3896 14136 3924
rect 15381 3927 15439 3933
rect 13688 3884 13694 3896
rect 15381 3893 15393 3927
rect 15427 3924 15439 3927
rect 16684 3924 16712 3964
rect 18370 3961 18382 3964
rect 18416 3961 18428 3995
rect 19886 3992 19892 4004
rect 18370 3955 18428 3961
rect 19168 3964 19892 3992
rect 17862 3924 17868 3936
rect 15427 3896 16712 3924
rect 17823 3896 17868 3924
rect 15427 3893 15439 3896
rect 15381 3887 15439 3893
rect 17862 3884 17868 3896
rect 17920 3884 17926 3936
rect 18046 3884 18052 3936
rect 18104 3924 18110 3936
rect 19168 3924 19196 3964
rect 19886 3952 19892 3964
rect 19944 3952 19950 4004
rect 19981 3995 20039 4001
rect 19981 3961 19993 3995
rect 20027 3992 20039 3995
rect 20070 3992 20076 4004
rect 20027 3964 20076 3992
rect 20027 3961 20039 3964
rect 19981 3955 20039 3961
rect 20070 3952 20076 3964
rect 20128 3952 20134 4004
rect 21450 3952 21456 4004
rect 21508 3992 21514 4004
rect 22002 3992 22008 4004
rect 21508 3964 22008 3992
rect 21508 3952 21514 3964
rect 22002 3952 22008 3964
rect 22060 3952 22066 4004
rect 22094 3952 22100 4004
rect 22152 3992 22158 4004
rect 24136 3992 24164 4020
rect 22152 3964 22197 3992
rect 23446 3964 24164 3992
rect 22152 3952 22158 3964
rect 18104 3896 19196 3924
rect 18104 3884 18110 3896
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 20990 3924 20996 3936
rect 20772 3896 20996 3924
rect 20772 3884 20778 3896
rect 20990 3884 20996 3896
rect 21048 3924 21054 3936
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 21048 3896 21097 3924
rect 21048 3884 21054 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 23017 3927 23075 3933
rect 23017 3924 23029 3927
rect 22244 3896 23029 3924
rect 22244 3884 22250 3896
rect 23017 3893 23029 3896
rect 23063 3924 23075 3927
rect 23446 3924 23474 3964
rect 23750 3924 23756 3936
rect 23063 3896 23474 3924
rect 23711 3896 23756 3924
rect 23063 3893 23075 3896
rect 23017 3887 23075 3893
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 25148 3933 25176 4032
rect 25225 4029 25237 4063
rect 25271 4029 25283 4063
rect 25225 4023 25283 4029
rect 25133 3927 25191 3933
rect 25133 3893 25145 3927
rect 25179 3924 25191 3927
rect 25498 3924 25504 3936
rect 25179 3896 25504 3924
rect 25179 3893 25191 3896
rect 25133 3887 25191 3893
rect 25498 3884 25504 3896
rect 25556 3884 25562 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2682 3720 2688 3732
rect 2643 3692 2688 3720
rect 2682 3680 2688 3692
rect 2740 3720 2746 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 2740 3692 3433 3720
rect 2740 3680 2746 3692
rect 3421 3689 3433 3692
rect 3467 3720 3479 3723
rect 3605 3723 3663 3729
rect 3605 3720 3617 3723
rect 3467 3692 3617 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 3605 3689 3617 3692
rect 3651 3689 3663 3723
rect 3605 3683 3663 3689
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 3752 3692 3801 3720
rect 3752 3680 3758 3692
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 4614 3720 4620 3732
rect 3789 3683 3847 3689
rect 3896 3692 4620 3720
rect 1535 3655 1593 3661
rect 1535 3621 1547 3655
rect 1581 3652 1593 3655
rect 3896 3652 3924 3692
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5353 3723 5411 3729
rect 5353 3720 5365 3723
rect 5132 3692 5365 3720
rect 5132 3680 5138 3692
rect 5353 3689 5365 3692
rect 5399 3720 5411 3723
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 5399 3692 5641 3720
rect 5399 3689 5411 3692
rect 5353 3683 5411 3689
rect 5629 3689 5641 3692
rect 5675 3689 5687 3723
rect 5629 3683 5687 3689
rect 5736 3692 8340 3720
rect 1581 3624 3924 3652
rect 1581 3621 1593 3624
rect 1535 3615 1593 3621
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 4249 3655 4307 3661
rect 4249 3652 4261 3655
rect 4028 3624 4261 3652
rect 4028 3612 4034 3624
rect 4249 3621 4261 3624
rect 4295 3621 4307 3655
rect 4249 3615 4307 3621
rect 4522 3612 4528 3664
rect 4580 3652 4586 3664
rect 4754 3655 4812 3661
rect 4754 3652 4766 3655
rect 4580 3624 4766 3652
rect 4580 3612 4586 3624
rect 4754 3621 4766 3624
rect 4800 3621 4812 3655
rect 4754 3615 4812 3621
rect 4982 3612 4988 3664
rect 5040 3652 5046 3664
rect 5736 3652 5764 3692
rect 5040 3624 5764 3652
rect 5040 3612 5046 3624
rect 7006 3612 7012 3664
rect 7064 3652 7070 3664
rect 7374 3652 7380 3664
rect 7064 3624 7380 3652
rect 7064 3612 7070 3624
rect 7374 3612 7380 3624
rect 7432 3612 7438 3664
rect 7929 3655 7987 3661
rect 7929 3621 7941 3655
rect 7975 3652 7987 3655
rect 8202 3652 8208 3664
rect 7975 3624 8208 3652
rect 7975 3621 7987 3624
rect 7929 3615 7987 3621
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 8312 3652 8340 3692
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8904 3692 9045 3720
rect 8904 3680 8910 3692
rect 9033 3689 9045 3692
rect 9079 3720 9091 3723
rect 9217 3723 9275 3729
rect 9217 3720 9229 3723
rect 9079 3692 9229 3720
rect 9079 3689 9091 3692
rect 9033 3683 9091 3689
rect 9217 3689 9229 3692
rect 9263 3689 9275 3723
rect 9217 3683 9275 3689
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9861 3723 9919 3729
rect 9861 3720 9873 3723
rect 9732 3692 9873 3720
rect 9732 3680 9738 3692
rect 9861 3689 9873 3692
rect 9907 3689 9919 3723
rect 9861 3683 9919 3689
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 10192 3692 10241 3720
rect 10192 3680 10198 3692
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 10229 3683 10287 3689
rect 10505 3723 10563 3729
rect 10505 3689 10517 3723
rect 10551 3720 10563 3723
rect 11609 3723 11667 3729
rect 11609 3720 11621 3723
rect 10551 3692 11621 3720
rect 10551 3689 10563 3692
rect 10505 3683 10563 3689
rect 11609 3689 11621 3692
rect 11655 3689 11667 3723
rect 11609 3683 11667 3689
rect 16390 3680 16396 3732
rect 16448 3720 16454 3732
rect 16853 3723 16911 3729
rect 16853 3720 16865 3723
rect 16448 3692 16865 3720
rect 16448 3680 16454 3692
rect 16853 3689 16865 3692
rect 16899 3720 16911 3723
rect 18230 3720 18236 3732
rect 16899 3692 18236 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 19337 3723 19395 3729
rect 19337 3720 19349 3723
rect 18840 3692 19349 3720
rect 18840 3680 18846 3692
rect 19337 3689 19349 3692
rect 19383 3720 19395 3723
rect 20438 3720 20444 3732
rect 19383 3692 20444 3720
rect 19383 3689 19395 3692
rect 19337 3683 19395 3689
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 21082 3680 21088 3732
rect 21140 3720 21146 3732
rect 21177 3723 21235 3729
rect 21177 3720 21189 3723
rect 21140 3692 21189 3720
rect 21140 3680 21146 3692
rect 21177 3689 21189 3692
rect 21223 3720 21235 3723
rect 22646 3720 22652 3732
rect 21223 3692 21956 3720
rect 22607 3692 22652 3720
rect 21223 3689 21235 3692
rect 21177 3683 21235 3689
rect 12161 3655 12219 3661
rect 12161 3652 12173 3655
rect 8312 3624 12173 3652
rect 12161 3621 12173 3624
rect 12207 3652 12219 3655
rect 12989 3655 13047 3661
rect 12989 3652 13001 3655
rect 12207 3624 13001 3652
rect 12207 3621 12219 3624
rect 12161 3615 12219 3621
rect 12989 3621 13001 3624
rect 13035 3621 13047 3655
rect 12989 3615 13047 3621
rect 13814 3612 13820 3664
rect 13872 3652 13878 3664
rect 14366 3652 14372 3664
rect 13872 3624 13917 3652
rect 14327 3624 14372 3652
rect 13872 3612 13878 3624
rect 14366 3612 14372 3624
rect 14424 3612 14430 3664
rect 15470 3652 15476 3664
rect 15431 3624 15476 3652
rect 15470 3612 15476 3624
rect 15528 3612 15534 3664
rect 16025 3655 16083 3661
rect 16025 3621 16037 3655
rect 16071 3652 16083 3655
rect 16206 3652 16212 3664
rect 16071 3624 16212 3652
rect 16071 3621 16083 3624
rect 16025 3615 16083 3621
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 16485 3655 16543 3661
rect 16485 3621 16497 3655
rect 16531 3652 16543 3655
rect 16574 3652 16580 3664
rect 16531 3624 16580 3652
rect 16531 3621 16543 3624
rect 16485 3615 16543 3621
rect 16574 3612 16580 3624
rect 16632 3652 16638 3664
rect 18322 3652 18328 3664
rect 16632 3624 18328 3652
rect 16632 3612 16638 3624
rect 18322 3612 18328 3624
rect 18380 3652 18386 3664
rect 18417 3655 18475 3661
rect 18417 3652 18429 3655
rect 18380 3624 18429 3652
rect 18380 3612 18386 3624
rect 18417 3621 18429 3624
rect 18463 3621 18475 3655
rect 18966 3652 18972 3664
rect 18927 3624 18972 3652
rect 18417 3615 18475 3621
rect 18966 3612 18972 3624
rect 19024 3652 19030 3664
rect 19024 3624 19932 3652
rect 19024 3612 19030 3624
rect 106 3544 112 3596
rect 164 3584 170 3596
rect 1448 3587 1506 3593
rect 1448 3584 1460 3587
rect 164 3556 1460 3584
rect 164 3544 170 3556
rect 1448 3553 1460 3556
rect 1494 3584 1506 3587
rect 1670 3584 1676 3596
rect 1494 3556 1676 3584
rect 1494 3553 1506 3556
rect 1448 3547 1506 3553
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 3053 3587 3111 3593
rect 3053 3553 3065 3587
rect 3099 3553 3111 3587
rect 3053 3547 3111 3553
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3516 2007 3519
rect 2222 3516 2228 3528
rect 1995 3488 2228 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3068 3516 3096 3547
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 4212 3556 4445 3584
rect 4212 3544 4218 3556
rect 4433 3553 4445 3556
rect 4479 3584 4491 3587
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 4479 3556 6009 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 6086 3544 6092 3596
rect 6144 3584 6150 3596
rect 6181 3587 6239 3593
rect 6181 3584 6193 3587
rect 6144 3556 6193 3584
rect 6144 3544 6150 3556
rect 6181 3553 6193 3556
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 9217 3587 9275 3593
rect 9217 3553 9229 3587
rect 9263 3584 9275 3587
rect 10505 3587 10563 3593
rect 10505 3584 10517 3587
rect 9263 3556 10517 3584
rect 9263 3553 9275 3556
rect 9217 3547 9275 3553
rect 10505 3553 10517 3556
rect 10551 3584 10563 3587
rect 10594 3584 10600 3596
rect 10551 3556 10600 3584
rect 10551 3553 10563 3556
rect 10505 3547 10563 3553
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 12250 3584 12256 3596
rect 10777 3556 12256 3584
rect 6104 3516 6132 3544
rect 7282 3516 7288 3528
rect 2924 3488 6132 3516
rect 7195 3488 7288 3516
rect 2924 3476 2930 3488
rect 7282 3476 7288 3488
rect 7340 3516 7346 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7340 3488 8217 3516
rect 7340 3476 7346 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 10777 3516 10805 3556
rect 12250 3544 12256 3556
rect 12308 3584 12314 3596
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 12308 3556 12357 3584
rect 12308 3544 12314 3556
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 17000 3556 17141 3584
rect 17000 3544 17006 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 19242 3544 19248 3596
rect 19300 3584 19306 3596
rect 19794 3584 19800 3596
rect 19300 3556 19800 3584
rect 19300 3544 19306 3556
rect 19794 3544 19800 3556
rect 19852 3544 19858 3596
rect 19904 3584 19932 3624
rect 19978 3612 19984 3664
rect 20036 3652 20042 3664
rect 20257 3655 20315 3661
rect 20257 3652 20269 3655
rect 20036 3624 20269 3652
rect 20036 3612 20042 3624
rect 20257 3621 20269 3624
rect 20303 3621 20315 3655
rect 20257 3615 20315 3621
rect 21726 3612 21732 3664
rect 21784 3652 21790 3664
rect 21821 3655 21879 3661
rect 21821 3652 21833 3655
rect 21784 3624 21833 3652
rect 21784 3612 21790 3624
rect 21821 3621 21833 3624
rect 21867 3621 21879 3655
rect 21928 3652 21956 3692
rect 22646 3680 22652 3692
rect 22704 3680 22710 3732
rect 22738 3680 22744 3732
rect 22796 3720 22802 3732
rect 24857 3723 24915 3729
rect 24857 3720 24869 3723
rect 22796 3692 24869 3720
rect 22796 3680 22802 3692
rect 24857 3689 24869 3692
rect 24903 3689 24915 3723
rect 24857 3683 24915 3689
rect 23750 3652 23756 3664
rect 21928 3624 23756 3652
rect 21821 3615 21879 3621
rect 23750 3612 23756 3624
rect 23808 3612 23814 3664
rect 21450 3584 21456 3596
rect 19904 3556 21456 3584
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 22373 3587 22431 3593
rect 22373 3553 22385 3587
rect 22419 3584 22431 3587
rect 22462 3584 22468 3596
rect 22419 3556 22468 3584
rect 22419 3553 22431 3556
rect 22373 3547 22431 3553
rect 22462 3544 22468 3556
rect 22520 3544 22526 3596
rect 23290 3584 23296 3596
rect 23251 3556 23296 3584
rect 23290 3544 23296 3556
rect 23348 3544 23354 3596
rect 23661 3587 23719 3593
rect 23661 3584 23673 3587
rect 23492 3556 23673 3584
rect 9364 3488 10805 3516
rect 10965 3519 11023 3525
rect 9364 3476 9370 3488
rect 10965 3485 10977 3519
rect 11011 3516 11023 3519
rect 11790 3516 11796 3528
rect 11011 3488 11796 3516
rect 11011 3485 11023 3488
rect 10965 3479 11023 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 14458 3516 14464 3528
rect 13771 3488 14464 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 14458 3476 14464 3488
rect 14516 3516 14522 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 14516 3488 14657 3516
rect 14516 3476 14522 3488
rect 14645 3485 14657 3488
rect 14691 3485 14703 3519
rect 14645 3479 14703 3485
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15378 3516 15384 3528
rect 15151 3488 15384 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3516 17831 3519
rect 18325 3519 18383 3525
rect 18325 3516 18337 3519
rect 17819 3488 18337 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 18325 3485 18337 3488
rect 18371 3516 18383 3519
rect 19334 3516 19340 3528
rect 18371 3488 19340 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 21729 3519 21787 3525
rect 21729 3485 21741 3519
rect 21775 3516 21787 3519
rect 21818 3516 21824 3528
rect 21775 3488 21824 3516
rect 21775 3485 21787 3488
rect 21729 3479 21787 3485
rect 21818 3476 21824 3488
rect 21876 3476 21882 3528
rect 3605 3451 3663 3457
rect 3605 3417 3617 3451
rect 3651 3448 3663 3451
rect 3651 3420 4154 3448
rect 3651 3417 3663 3420
rect 3605 3411 3663 3417
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2096 3352 2237 3380
rect 2096 3340 2102 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 4126 3380 4154 3420
rect 4890 3408 4896 3460
rect 4948 3448 4954 3460
rect 6365 3451 6423 3457
rect 6365 3448 6377 3451
rect 4948 3420 6377 3448
rect 4948 3408 4954 3420
rect 6365 3417 6377 3420
rect 6411 3448 6423 3451
rect 6454 3448 6460 3460
rect 6411 3420 6460 3448
rect 6411 3417 6423 3420
rect 6365 3411 6423 3417
rect 6454 3408 6460 3420
rect 6512 3408 6518 3460
rect 6546 3408 6552 3460
rect 6604 3448 6610 3460
rect 8665 3451 8723 3457
rect 8665 3448 8677 3451
rect 6604 3420 8677 3448
rect 6604 3408 6610 3420
rect 8665 3417 8677 3420
rect 8711 3448 8723 3451
rect 9122 3448 9128 3460
rect 8711 3420 9128 3448
rect 8711 3417 8723 3420
rect 8665 3411 8723 3417
rect 9122 3408 9128 3420
rect 9180 3408 9186 3460
rect 10226 3408 10232 3460
rect 10284 3448 10290 3460
rect 11977 3451 12035 3457
rect 11977 3448 11989 3451
rect 10284 3420 11989 3448
rect 10284 3408 10290 3420
rect 10980 3392 11008 3420
rect 11977 3417 11989 3420
rect 12023 3448 12035 3451
rect 17313 3451 17371 3457
rect 12023 3420 12480 3448
rect 12023 3417 12035 3420
rect 11977 3411 12035 3417
rect 6730 3380 6736 3392
rect 4126 3352 6736 3380
rect 2225 3343 2283 3349
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 7006 3380 7012 3392
rect 6967 3352 7012 3380
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 9493 3383 9551 3389
rect 9493 3349 9505 3383
rect 9539 3380 9551 3383
rect 9858 3380 9864 3392
rect 9539 3352 9864 3380
rect 9539 3349 9551 3352
rect 9493 3343 9551 3349
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 10410 3340 10416 3392
rect 10468 3380 10474 3392
rect 10686 3380 10692 3392
rect 10468 3352 10692 3380
rect 10468 3340 10474 3352
rect 10686 3340 10692 3352
rect 10744 3389 10750 3392
rect 10744 3383 10793 3389
rect 10744 3349 10747 3383
rect 10781 3349 10793 3383
rect 10870 3380 10876 3392
rect 10831 3352 10876 3380
rect 10744 3343 10793 3349
rect 10744 3340 10750 3343
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 10962 3340 10968 3392
rect 11020 3340 11026 3392
rect 11241 3383 11299 3389
rect 11241 3349 11253 3383
rect 11287 3380 11299 3383
rect 11514 3380 11520 3392
rect 11287 3352 11520 3380
rect 11287 3349 11299 3352
rect 11241 3343 11299 3349
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 12452 3389 12480 3420
rect 17313 3417 17325 3451
rect 17359 3448 17371 3451
rect 19981 3451 20039 3457
rect 17359 3420 18689 3448
rect 17359 3417 17371 3420
rect 17313 3411 17371 3417
rect 12437 3383 12495 3389
rect 12437 3349 12449 3383
rect 12483 3349 12495 3383
rect 13354 3380 13360 3392
rect 13315 3352 13360 3380
rect 12437 3343 12495 3349
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 18138 3380 18144 3392
rect 18099 3352 18144 3380
rect 18138 3340 18144 3352
rect 18196 3340 18202 3392
rect 18661 3380 18689 3420
rect 19981 3417 19993 3451
rect 20027 3448 20039 3451
rect 22186 3448 22192 3460
rect 20027 3420 22192 3448
rect 20027 3417 20039 3420
rect 19981 3411 20039 3417
rect 22186 3408 22192 3420
rect 22244 3408 22250 3460
rect 22480 3448 22508 3544
rect 22554 3476 22560 3528
rect 22612 3516 22618 3528
rect 23109 3519 23167 3525
rect 23109 3516 23121 3519
rect 22612 3488 23121 3516
rect 22612 3476 22618 3488
rect 23109 3485 23121 3488
rect 23155 3516 23167 3519
rect 23492 3516 23520 3556
rect 23661 3553 23673 3556
rect 23707 3553 23719 3587
rect 23661 3547 23719 3553
rect 24762 3544 24768 3596
rect 24820 3584 24826 3596
rect 25038 3584 25044 3596
rect 24820 3556 25044 3584
rect 24820 3544 24826 3556
rect 25038 3544 25044 3556
rect 25096 3544 25102 3596
rect 25317 3587 25375 3593
rect 25317 3553 25329 3587
rect 25363 3584 25375 3587
rect 25498 3584 25504 3596
rect 25363 3556 25504 3584
rect 25363 3553 25375 3556
rect 25317 3547 25375 3553
rect 25498 3544 25504 3556
rect 25556 3544 25562 3596
rect 23750 3516 23756 3528
rect 23155 3488 23520 3516
rect 23711 3488 23756 3516
rect 23155 3485 23167 3488
rect 23109 3479 23167 3485
rect 23750 3476 23756 3488
rect 23808 3476 23814 3528
rect 24581 3451 24639 3457
rect 24581 3448 24593 3451
rect 22480 3420 24593 3448
rect 24581 3417 24593 3420
rect 24627 3417 24639 3451
rect 24581 3411 24639 3417
rect 20438 3380 20444 3392
rect 18661 3352 20444 3380
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 22646 3340 22652 3392
rect 22704 3380 22710 3392
rect 23290 3380 23296 3392
rect 22704 3352 23296 3380
rect 22704 3340 22710 3352
rect 23290 3340 23296 3352
rect 23348 3340 23354 3392
rect 24026 3340 24032 3392
rect 24084 3380 24090 3392
rect 24213 3383 24271 3389
rect 24213 3380 24225 3383
rect 24084 3352 24225 3380
rect 24084 3340 24090 3352
rect 24213 3349 24225 3352
rect 24259 3349 24271 3383
rect 24213 3343 24271 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2866 3176 2872 3188
rect 2827 3148 2872 3176
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 3602 3136 3608 3188
rect 3660 3176 3666 3188
rect 6546 3176 6552 3188
rect 3660 3148 6552 3176
rect 3660 3136 3666 3148
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 7190 3176 7196 3188
rect 6687 3148 7196 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7432 3148 7849 3176
rect 7432 3136 7438 3148
rect 7837 3145 7849 3148
rect 7883 3176 7895 3179
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 7883 3148 8125 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8113 3145 8125 3148
rect 8159 3145 8171 3179
rect 9677 3179 9735 3185
rect 9677 3176 9689 3179
rect 8113 3139 8171 3145
rect 8496 3148 9689 3176
rect 4522 3108 4528 3120
rect 4483 3080 4528 3108
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 5534 3108 5540 3120
rect 5495 3080 5540 3108
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 6730 3068 6736 3120
rect 6788 3108 6794 3120
rect 8496 3108 8524 3148
rect 9677 3145 9689 3148
rect 9723 3145 9735 3179
rect 9677 3139 9735 3145
rect 6788 3080 8524 3108
rect 8573 3111 8631 3117
rect 6788 3068 6794 3080
rect 8573 3077 8585 3111
rect 8619 3108 8631 3111
rect 8619 3080 8984 3108
rect 8619 3077 8631 3080
rect 8573 3071 8631 3077
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 4338 3040 4344 3052
rect 2547 3012 4344 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 4338 3000 4344 3012
rect 4396 3000 4402 3052
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4672 3012 4997 3040
rect 4672 3000 4678 3012
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 8018 3040 8024 3052
rect 5031 3012 8024 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 8846 3040 8852 3052
rect 8352 3012 8852 3040
rect 8352 3000 8358 3012
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 8956 3040 8984 3080
rect 9398 3040 9404 3052
rect 8956 3012 9404 3040
rect 2222 2972 2228 2984
rect 2183 2944 2228 2972
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 3418 2972 3424 2984
rect 3379 2944 3424 2972
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 3602 2932 3608 2984
rect 3660 2972 3666 2984
rect 3789 2975 3847 2981
rect 3789 2972 3801 2975
rect 3660 2944 3801 2972
rect 3660 2932 3666 2944
rect 3789 2941 3801 2944
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 6917 2975 6975 2981
rect 6917 2941 6929 2975
rect 6963 2972 6975 2975
rect 7006 2972 7012 2984
rect 6963 2944 7012 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 7006 2932 7012 2944
rect 7064 2972 7070 2984
rect 8956 2981 8984 3012
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 9692 3040 9720 3139
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 10008 3148 10057 3176
rect 10008 3136 10014 3148
rect 10045 3145 10057 3148
rect 10091 3176 10103 3179
rect 12250 3176 12256 3188
rect 10091 3148 10640 3176
rect 12211 3148 12256 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 9766 3068 9772 3120
rect 9824 3108 9830 3120
rect 10410 3117 10416 3120
rect 10367 3111 10416 3117
rect 10367 3108 10379 3111
rect 9824 3080 10379 3108
rect 9824 3068 9830 3080
rect 10367 3077 10379 3080
rect 10413 3077 10416 3111
rect 10367 3071 10416 3077
rect 10410 3068 10416 3071
rect 10468 3068 10474 3120
rect 10505 3111 10563 3117
rect 10505 3077 10517 3111
rect 10551 3077 10563 3111
rect 10505 3071 10563 3077
rect 10520 3040 10548 3071
rect 10612 3049 10640 3148
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 13725 3179 13783 3185
rect 13725 3145 13737 3179
rect 13771 3176 13783 3179
rect 13814 3176 13820 3188
rect 13771 3148 13820 3176
rect 13771 3145 13783 3148
rect 13725 3139 13783 3145
rect 13814 3136 13820 3148
rect 13872 3176 13878 3188
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 13872 3148 14013 3176
rect 13872 3136 13878 3148
rect 14001 3145 14013 3148
rect 14047 3145 14059 3179
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 14001 3139 14059 3145
rect 15470 3136 15476 3148
rect 15528 3176 15534 3188
rect 15749 3179 15807 3185
rect 15749 3176 15761 3179
rect 15528 3148 15761 3176
rect 15528 3136 15534 3148
rect 15749 3145 15761 3148
rect 15795 3176 15807 3179
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 15795 3148 16129 3176
rect 15795 3145 15807 3148
rect 15749 3139 15807 3145
rect 16117 3145 16129 3148
rect 16163 3176 16175 3179
rect 16482 3176 16488 3188
rect 16163 3148 16488 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 17000 3148 17325 3176
rect 17000 3136 17006 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 19794 3176 19800 3188
rect 19755 3148 19800 3176
rect 17313 3139 17371 3145
rect 19794 3136 19800 3148
rect 19852 3136 19858 3188
rect 21266 3136 21272 3188
rect 21324 3176 21330 3188
rect 22373 3179 22431 3185
rect 22373 3176 22385 3179
rect 21324 3148 22385 3176
rect 21324 3136 21330 3148
rect 22373 3145 22385 3148
rect 22419 3176 22431 3179
rect 22646 3176 22652 3188
rect 22419 3148 22652 3176
rect 22419 3145 22431 3148
rect 22373 3139 22431 3145
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 22830 3176 22836 3188
rect 22791 3148 22836 3176
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 23109 3179 23167 3185
rect 23109 3145 23121 3179
rect 23155 3176 23167 3179
rect 23474 3176 23480 3188
rect 23155 3148 23480 3176
rect 23155 3145 23167 3148
rect 23109 3139 23167 3145
rect 18414 3068 18420 3120
rect 18472 3108 18478 3120
rect 22278 3108 22284 3120
rect 18472 3080 22284 3108
rect 18472 3068 18478 3080
rect 22278 3068 22284 3080
rect 22336 3068 22342 3120
rect 9692 3012 10548 3040
rect 8941 2975 8999 2981
rect 7064 2944 8616 2972
rect 7064 2932 7070 2944
rect 4065 2907 4123 2913
rect 4065 2873 4077 2907
rect 4111 2904 4123 2907
rect 4798 2904 4804 2916
rect 4111 2876 4804 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 4798 2864 4804 2876
rect 4856 2864 4862 2916
rect 5074 2864 5080 2916
rect 5132 2904 5138 2916
rect 5132 2876 5177 2904
rect 5132 2864 5138 2876
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 2498 2796 2504 2848
rect 2556 2836 2562 2848
rect 3234 2836 3240 2848
rect 2556 2808 3240 2836
rect 2556 2796 2562 2808
rect 3234 2796 3240 2808
rect 3292 2796 3298 2848
rect 6086 2796 6092 2848
rect 6144 2836 6150 2848
rect 6181 2839 6239 2845
rect 6181 2836 6193 2839
rect 6144 2808 6193 2836
rect 6144 2796 6150 2808
rect 6181 2805 6193 2808
rect 6227 2805 6239 2839
rect 6181 2799 6239 2805
rect 7190 2796 7196 2848
rect 7248 2836 7254 2848
rect 7285 2839 7343 2845
rect 7285 2836 7297 2839
rect 7248 2808 7297 2836
rect 7248 2796 7254 2808
rect 7285 2805 7297 2808
rect 7331 2805 7343 2839
rect 8588 2836 8616 2944
rect 8941 2941 8953 2975
rect 8987 2941 8999 2975
rect 9122 2972 9128 2984
rect 9083 2944 9128 2972
rect 8941 2935 8999 2941
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 10226 2972 10232 2984
rect 10187 2944 10232 2972
rect 10226 2932 10232 2944
rect 10284 2932 10290 2984
rect 10520 2972 10548 3012
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 16390 3040 16396 3052
rect 16351 3012 16396 3040
rect 10597 3003 10655 3009
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 18966 3000 18972 3052
rect 19024 3040 19030 3052
rect 19061 3043 19119 3049
rect 19061 3040 19073 3043
rect 19024 3012 19073 3040
rect 19024 3000 19030 3012
rect 19061 3009 19073 3012
rect 19107 3009 19119 3043
rect 19061 3003 19119 3009
rect 20349 3043 20407 3049
rect 20349 3009 20361 3043
rect 20395 3040 20407 3043
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 20395 3012 20821 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 20809 3009 20821 3012
rect 20855 3040 20867 3043
rect 22738 3040 22744 3052
rect 20855 3012 22744 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 23124 3040 23152 3139
rect 23474 3136 23480 3148
rect 23532 3136 23538 3188
rect 24673 3179 24731 3185
rect 24673 3176 24685 3179
rect 23823 3148 24685 3176
rect 23658 3068 23664 3120
rect 23716 3108 23722 3120
rect 23823 3117 23851 3148
rect 24673 3145 24685 3148
rect 24719 3145 24731 3179
rect 25038 3176 25044 3188
rect 24999 3148 25044 3176
rect 24673 3139 24731 3145
rect 25038 3136 25044 3148
rect 25096 3136 25102 3188
rect 23799 3111 23857 3117
rect 23799 3108 23811 3111
rect 23716 3080 23811 3108
rect 23716 3068 23722 3080
rect 23799 3077 23811 3080
rect 23845 3077 23857 3111
rect 23934 3108 23940 3120
rect 23895 3080 23940 3108
rect 23799 3071 23857 3077
rect 23934 3068 23940 3080
rect 23992 3068 23998 3120
rect 25409 3111 25467 3117
rect 25409 3108 25421 3111
rect 24320 3080 25421 3108
rect 24026 3040 24032 3052
rect 23032 3012 23152 3040
rect 23987 3012 24032 3040
rect 10870 2972 10876 2984
rect 10520 2944 10876 2972
rect 10870 2932 10876 2944
rect 10928 2972 10934 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 10928 2944 11253 2972
rect 10928 2932 10934 2944
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 11698 2932 11704 2984
rect 11756 2972 11762 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 11756 2944 12817 2972
rect 11756 2932 11762 2944
rect 12805 2941 12817 2944
rect 12851 2972 12863 2975
rect 13354 2972 13360 2984
rect 12851 2944 13360 2972
rect 12851 2941 12863 2944
rect 12805 2935 12863 2941
rect 13354 2932 13360 2944
rect 13412 2932 13418 2984
rect 14553 2975 14611 2981
rect 14553 2941 14565 2975
rect 14599 2972 14611 2975
rect 14642 2972 14648 2984
rect 14599 2944 14648 2972
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 22624 2975 22682 2981
rect 22624 2941 22636 2975
rect 22670 2972 22682 2975
rect 23032 2972 23060 3012
rect 24026 3000 24032 3012
rect 24084 3000 24090 3052
rect 24118 3000 24124 3052
rect 24176 3040 24182 3052
rect 24176 3012 24221 3040
rect 24176 3000 24182 3012
rect 22670 2944 23060 2972
rect 22670 2941 22682 2944
rect 22624 2935 22682 2941
rect 23106 2932 23112 2984
rect 23164 2972 23170 2984
rect 23385 2975 23443 2981
rect 23385 2972 23397 2975
rect 23164 2944 23397 2972
rect 23164 2932 23170 2944
rect 23385 2941 23397 2944
rect 23431 2972 23443 2975
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23431 2944 23673 2972
rect 23431 2941 23443 2944
rect 23385 2935 23443 2941
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 23661 2935 23719 2941
rect 23842 2932 23848 2984
rect 23900 2972 23906 2984
rect 24320 2972 24348 3080
rect 25409 3077 25421 3080
rect 25455 3077 25467 3111
rect 25409 3071 25467 3077
rect 23900 2944 24348 2972
rect 25225 2975 25283 2981
rect 23900 2932 23906 2944
rect 25225 2941 25237 2975
rect 25271 2941 25283 2975
rect 25225 2935 25283 2941
rect 9214 2864 9220 2916
rect 9272 2904 9278 2916
rect 10965 2907 11023 2913
rect 10965 2904 10977 2907
rect 9272 2876 10977 2904
rect 9272 2864 9278 2876
rect 10965 2873 10977 2876
rect 11011 2873 11023 2907
rect 10965 2867 11023 2873
rect 13126 2907 13184 2913
rect 13126 2873 13138 2907
rect 13172 2904 13184 2907
rect 14369 2907 14427 2913
rect 14369 2904 14381 2907
rect 13172 2876 14381 2904
rect 13172 2873 13184 2876
rect 13126 2867 13184 2873
rect 14369 2873 14381 2876
rect 14415 2904 14427 2907
rect 14874 2907 14932 2913
rect 14874 2904 14886 2907
rect 14415 2876 14886 2904
rect 14415 2873 14427 2876
rect 14369 2867 14427 2873
rect 14874 2873 14886 2876
rect 14920 2904 14932 2907
rect 15654 2904 15660 2916
rect 14920 2876 15660 2904
rect 14920 2873 14932 2876
rect 14874 2867 14932 2873
rect 8757 2839 8815 2845
rect 8757 2836 8769 2839
rect 8588 2808 8769 2836
rect 7285 2799 7343 2805
rect 8757 2805 8769 2808
rect 8803 2805 8815 2839
rect 8757 2799 8815 2805
rect 9858 2796 9864 2848
rect 9916 2836 9922 2848
rect 11701 2839 11759 2845
rect 11701 2836 11713 2839
rect 9916 2808 11713 2836
rect 9916 2796 9922 2808
rect 11701 2805 11713 2808
rect 11747 2836 11759 2839
rect 11790 2836 11796 2848
rect 11747 2808 11796 2836
rect 11747 2805 11759 2808
rect 11701 2799 11759 2805
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12618 2836 12624 2848
rect 12579 2808 12624 2836
rect 12618 2796 12624 2808
rect 12676 2836 12682 2848
rect 13141 2836 13169 2867
rect 15654 2864 15660 2876
rect 15712 2904 15718 2916
rect 16206 2904 16212 2916
rect 15712 2876 16212 2904
rect 15712 2864 15718 2876
rect 16206 2864 16212 2876
rect 16264 2864 16270 2916
rect 16482 2864 16488 2916
rect 16540 2904 16546 2916
rect 18877 2907 18935 2913
rect 18877 2904 18889 2907
rect 16540 2876 16585 2904
rect 17788 2876 18889 2904
rect 16540 2864 16546 2876
rect 17788 2848 17816 2876
rect 18877 2873 18889 2876
rect 18923 2904 18935 2907
rect 19242 2904 19248 2916
rect 18923 2876 19248 2904
rect 18923 2873 18935 2876
rect 18877 2867 18935 2873
rect 19242 2864 19248 2876
rect 19300 2864 19306 2916
rect 20717 2907 20775 2913
rect 20717 2873 20729 2907
rect 20763 2904 20775 2907
rect 20990 2904 20996 2916
rect 20763 2876 20996 2904
rect 20763 2873 20775 2876
rect 20717 2867 20775 2873
rect 20990 2864 20996 2876
rect 21048 2904 21054 2916
rect 21130 2907 21188 2913
rect 21130 2904 21142 2907
rect 21048 2876 21142 2904
rect 21048 2864 21054 2876
rect 21130 2873 21142 2876
rect 21176 2873 21188 2907
rect 21130 2867 21188 2873
rect 21266 2864 21272 2916
rect 21324 2904 21330 2916
rect 25240 2904 25268 2935
rect 26145 2907 26203 2913
rect 26145 2904 26157 2907
rect 21324 2876 26157 2904
rect 21324 2864 21330 2876
rect 26145 2873 26157 2876
rect 26191 2873 26203 2907
rect 26145 2867 26203 2873
rect 17770 2836 17776 2848
rect 12676 2808 13169 2836
rect 17731 2808 17776 2836
rect 12676 2796 12682 2808
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18322 2836 18328 2848
rect 18283 2808 18328 2836
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 21726 2836 21732 2848
rect 21687 2808 21732 2836
rect 21726 2796 21732 2808
rect 21784 2836 21790 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21784 2808 22017 2836
rect 21784 2796 21790 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 23290 2796 23296 2848
rect 23348 2836 23354 2848
rect 24210 2836 24216 2848
rect 23348 2808 24216 2836
rect 23348 2796 23354 2808
rect 24210 2796 24216 2808
rect 24268 2796 24274 2848
rect 25498 2796 25504 2848
rect 25556 2836 25562 2848
rect 25777 2839 25835 2845
rect 25777 2836 25789 2839
rect 25556 2808 25789 2836
rect 25556 2796 25562 2808
rect 25777 2805 25789 2808
rect 25823 2805 25835 2839
rect 25777 2799 25835 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 3418 2632 3424 2644
rect 3379 2604 3424 2632
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3660 2604 3801 2632
rect 3660 2592 3666 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 4522 2592 4528 2644
rect 4580 2632 4586 2644
rect 4893 2635 4951 2641
rect 4893 2632 4905 2635
rect 4580 2604 4905 2632
rect 4580 2592 4586 2604
rect 4893 2601 4905 2604
rect 4939 2601 4951 2635
rect 4893 2595 4951 2601
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 3436 2564 3464 2592
rect 2363 2536 3464 2564
rect 4908 2564 4936 2595
rect 5166 2592 5172 2644
rect 5224 2632 5230 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5224 2604 6009 2632
rect 5224 2592 5230 2604
rect 5997 2601 6009 2604
rect 6043 2632 6055 2635
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 6043 2604 6653 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 6641 2601 6653 2604
rect 6687 2632 6699 2635
rect 6914 2632 6920 2644
rect 6687 2604 6920 2632
rect 6687 2601 6699 2604
rect 6641 2595 6699 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 7024 2604 7941 2632
rect 5398 2567 5456 2573
rect 5398 2564 5410 2567
rect 4908 2536 5410 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 842 2456 848 2508
rect 900 2496 906 2508
rect 2700 2505 2728 2536
rect 5398 2533 5410 2536
rect 5444 2533 5456 2567
rect 5398 2527 5456 2533
rect 6362 2524 6368 2576
rect 6420 2564 6426 2576
rect 7024 2573 7052 2604
rect 7929 2601 7941 2604
rect 7975 2601 7987 2635
rect 7929 2595 7987 2601
rect 8018 2592 8024 2644
rect 8076 2632 8082 2644
rect 8297 2635 8355 2641
rect 8297 2632 8309 2635
rect 8076 2604 8309 2632
rect 8076 2592 8082 2604
rect 8297 2601 8309 2604
rect 8343 2601 8355 2635
rect 8297 2595 8355 2601
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 8527 2604 9597 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 9585 2601 9597 2604
rect 9631 2632 9643 2635
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 9631 2604 10885 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 11882 2632 11888 2644
rect 10873 2595 10931 2601
rect 11256 2604 11888 2632
rect 7009 2567 7067 2573
rect 7009 2564 7021 2567
rect 6420 2536 7021 2564
rect 6420 2524 6426 2536
rect 7009 2533 7021 2536
rect 7055 2533 7067 2567
rect 7009 2527 7067 2533
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2564 7159 2567
rect 7190 2564 7196 2576
rect 7147 2536 7196 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 7650 2564 7656 2576
rect 7611 2536 7656 2564
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 11146 2564 11152 2576
rect 9140 2536 11152 2564
rect 1432 2499 1490 2505
rect 1432 2496 1444 2499
rect 900 2468 1444 2496
rect 900 2456 906 2468
rect 1432 2465 1444 2468
rect 1478 2496 1490 2499
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1478 2468 1869 2496
rect 1478 2465 1490 2468
rect 1432 2459 1490 2465
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2465 2743 2499
rect 2685 2459 2743 2465
rect 2961 2499 3019 2505
rect 2961 2465 2973 2499
rect 3007 2465 3019 2499
rect 2961 2459 3019 2465
rect 4132 2499 4190 2505
rect 4132 2465 4144 2499
rect 4178 2496 4190 2499
rect 4706 2496 4712 2508
rect 4178 2468 4712 2496
rect 4178 2465 4190 2468
rect 4132 2459 4190 2465
rect 2976 2360 3004 2459
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 9140 2505 9168 2536
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 5077 2499 5135 2505
rect 5077 2496 5089 2499
rect 4856 2468 5089 2496
rect 4856 2456 4862 2468
rect 5077 2465 5089 2468
rect 5123 2496 5135 2499
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5123 2468 6285 2496
rect 5123 2465 5135 2468
rect 5077 2459 5135 2465
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8711 2468 9137 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9582 2496 9588 2508
rect 9125 2459 9183 2465
rect 9232 2468 9588 2496
rect 3142 2428 3148 2440
rect 3103 2400 3148 2428
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 8680 2428 8708 2459
rect 4396 2400 8708 2428
rect 4396 2388 4402 2400
rect 4203 2363 4261 2369
rect 2976 2332 4154 2360
rect 1535 2295 1593 2301
rect 1535 2261 1547 2295
rect 1581 2292 1593 2295
rect 2130 2292 2136 2304
rect 1581 2264 2136 2292
rect 1581 2261 1593 2264
rect 1535 2255 1593 2261
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 4126 2292 4154 2332
rect 4203 2329 4215 2363
rect 4249 2360 4261 2363
rect 9232 2360 9260 2468
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 11256 2505 11284 2604
rect 11882 2592 11888 2604
rect 11940 2632 11946 2644
rect 11977 2635 12035 2641
rect 11977 2632 11989 2635
rect 11940 2604 11989 2632
rect 11940 2592 11946 2604
rect 11977 2601 11989 2604
rect 12023 2601 12035 2635
rect 13630 2632 13636 2644
rect 13591 2604 13636 2632
rect 11977 2595 12035 2601
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 16301 2635 16359 2641
rect 16301 2632 16313 2635
rect 16264 2604 16313 2632
rect 16264 2592 16270 2604
rect 16301 2601 16313 2604
rect 16347 2601 16359 2635
rect 16301 2595 16359 2601
rect 17405 2635 17463 2641
rect 17405 2601 17417 2635
rect 17451 2632 17463 2635
rect 17770 2632 17776 2644
rect 17451 2604 17776 2632
rect 17451 2601 17463 2604
rect 17405 2595 17463 2601
rect 11698 2564 11704 2576
rect 11659 2536 11704 2564
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 12618 2524 12624 2576
rect 12676 2564 12682 2576
rect 13034 2567 13092 2573
rect 13034 2564 13046 2567
rect 12676 2536 13046 2564
rect 12676 2524 12682 2536
rect 13034 2533 13046 2536
rect 13080 2533 13092 2567
rect 16316 2564 16344 2595
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 18322 2592 18328 2644
rect 18380 2632 18386 2644
rect 19245 2635 19303 2641
rect 19245 2632 19257 2635
rect 18380 2604 19257 2632
rect 18380 2592 18386 2604
rect 19245 2601 19257 2604
rect 19291 2601 19303 2635
rect 19245 2595 19303 2601
rect 20211 2635 20269 2641
rect 20211 2601 20223 2635
rect 20257 2632 20269 2635
rect 21266 2632 21272 2644
rect 20257 2604 21272 2632
rect 20257 2601 20269 2604
rect 20211 2595 20269 2601
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 21818 2592 21824 2644
rect 21876 2632 21882 2644
rect 22281 2635 22339 2641
rect 22281 2632 22293 2635
rect 21876 2604 22293 2632
rect 21876 2592 21882 2604
rect 22281 2601 22293 2604
rect 22327 2601 22339 2635
rect 22281 2595 22339 2601
rect 23845 2635 23903 2641
rect 23845 2601 23857 2635
rect 23891 2632 23903 2635
rect 23934 2632 23940 2644
rect 23891 2604 23940 2632
rect 23891 2601 23903 2604
rect 23845 2595 23903 2601
rect 16806 2567 16864 2573
rect 16806 2564 16818 2567
rect 16316 2536 16818 2564
rect 13034 2527 13092 2533
rect 16806 2533 16818 2536
rect 16852 2564 16864 2567
rect 17862 2564 17868 2576
rect 16852 2536 17868 2564
rect 16852 2533 16864 2536
rect 16806 2527 16864 2533
rect 17862 2524 17868 2536
rect 17920 2564 17926 2576
rect 18049 2567 18107 2573
rect 18049 2564 18061 2567
rect 17920 2536 18061 2564
rect 17920 2524 17926 2536
rect 18049 2533 18061 2536
rect 18095 2564 18107 2567
rect 18646 2567 18704 2573
rect 18646 2564 18658 2567
rect 18095 2536 18658 2564
rect 18095 2533 18107 2536
rect 18049 2527 18107 2533
rect 18646 2533 18658 2536
rect 18692 2533 18704 2567
rect 18646 2527 18704 2533
rect 20993 2567 21051 2573
rect 20993 2533 21005 2567
rect 21039 2564 21051 2567
rect 21453 2567 21511 2573
rect 21453 2564 21465 2567
rect 21039 2536 21465 2564
rect 21039 2533 21051 2536
rect 20993 2527 21051 2533
rect 21453 2533 21465 2536
rect 21499 2564 21511 2567
rect 21726 2564 21732 2576
rect 21499 2536 21732 2564
rect 21499 2533 21511 2536
rect 21453 2527 21511 2533
rect 21726 2524 21732 2536
rect 21784 2524 21790 2576
rect 22002 2564 22008 2576
rect 21963 2536 22008 2564
rect 22002 2524 22008 2536
rect 22060 2524 22066 2576
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9732 2468 9781 2496
rect 9732 2456 9738 2468
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 11241 2499 11299 2505
rect 11241 2465 11253 2499
rect 11287 2465 11299 2499
rect 11422 2496 11428 2508
rect 11383 2468 11428 2496
rect 11241 2459 11299 2465
rect 9784 2428 9812 2459
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 11572 2468 15485 2496
rect 11572 2456 11578 2468
rect 15473 2465 15485 2468
rect 15519 2496 15531 2499
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 15519 2468 15945 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 15933 2465 15945 2468
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 17819 2468 18337 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 18325 2465 18337 2468
rect 18371 2496 18383 2499
rect 18414 2496 18420 2508
rect 18371 2468 18420 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 19150 2456 19156 2508
rect 19208 2496 19214 2508
rect 20108 2499 20166 2505
rect 20108 2496 20120 2499
rect 19208 2468 20120 2496
rect 19208 2456 19214 2468
rect 20108 2465 20120 2468
rect 20154 2496 20166 2499
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20154 2468 20545 2496
rect 20154 2465 20166 2468
rect 20108 2459 20166 2465
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2496 22891 2499
rect 23477 2499 23535 2505
rect 23477 2496 23489 2499
rect 22879 2468 23489 2496
rect 22879 2465 22891 2468
rect 22833 2459 22891 2465
rect 23477 2465 23489 2468
rect 23523 2496 23535 2499
rect 23566 2496 23572 2508
rect 23523 2468 23572 2496
rect 23523 2465 23535 2468
rect 23477 2459 23535 2465
rect 23566 2456 23572 2468
rect 23624 2456 23630 2508
rect 12158 2428 12164 2440
rect 9784 2400 12164 2428
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 12710 2428 12716 2440
rect 12671 2400 12716 2428
rect 12710 2388 12716 2400
rect 12768 2428 12774 2440
rect 13909 2431 13967 2437
rect 13909 2428 13921 2431
rect 12768 2400 13921 2428
rect 12768 2388 12774 2400
rect 13909 2397 13921 2400
rect 13955 2397 13967 2431
rect 13909 2391 13967 2397
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 16482 2428 16488 2440
rect 15335 2400 16488 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 21358 2428 21364 2440
rect 21319 2400 21364 2428
rect 21358 2388 21364 2400
rect 21416 2388 21422 2440
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 23860 2428 23888 2595
rect 23934 2592 23940 2604
rect 23992 2592 23998 2644
rect 24118 2632 24124 2644
rect 24079 2604 24124 2632
rect 24118 2592 24124 2604
rect 24176 2592 24182 2644
rect 24857 2635 24915 2641
rect 24857 2601 24869 2635
rect 24903 2632 24915 2635
rect 25498 2632 25504 2644
rect 24903 2604 25504 2632
rect 24903 2601 24915 2604
rect 24857 2595 24915 2601
rect 25498 2592 25504 2604
rect 25556 2592 25562 2644
rect 25041 2567 25099 2573
rect 25041 2564 25053 2567
rect 24228 2536 25053 2564
rect 24228 2508 24256 2536
rect 25041 2533 25053 2536
rect 25087 2533 25099 2567
rect 25041 2527 25099 2533
rect 24210 2496 24216 2508
rect 24171 2468 24216 2496
rect 24210 2456 24216 2468
rect 24268 2456 24274 2508
rect 24581 2499 24639 2505
rect 24581 2465 24593 2499
rect 24627 2496 24639 2499
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 24627 2468 24869 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 24857 2459 24915 2465
rect 25314 2456 25320 2508
rect 25372 2496 25378 2508
rect 25660 2499 25718 2505
rect 25660 2496 25672 2499
rect 25372 2468 25672 2496
rect 25372 2456 25378 2468
rect 25660 2465 25672 2468
rect 25706 2496 25718 2499
rect 25706 2468 26188 2496
rect 25706 2465 25718 2468
rect 25660 2459 25718 2465
rect 21508 2400 23888 2428
rect 21508 2388 21514 2400
rect 9766 2360 9772 2372
rect 4249 2332 9260 2360
rect 9679 2332 9772 2360
rect 4249 2329 4261 2332
rect 4203 2323 4261 2329
rect 9766 2320 9772 2332
rect 9824 2360 9830 2372
rect 9824 2332 10088 2360
rect 9824 2320 9830 2332
rect 4617 2295 4675 2301
rect 4617 2292 4629 2295
rect 4126 2264 4629 2292
rect 4617 2261 4629 2264
rect 4663 2292 4675 2295
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 4663 2264 8493 2292
rect 4663 2261 4675 2264
rect 4617 2255 4675 2261
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 8754 2252 8760 2304
rect 8812 2292 8818 2304
rect 8849 2295 8907 2301
rect 8849 2292 8861 2295
rect 8812 2264 8861 2292
rect 8812 2252 8818 2264
rect 8849 2261 8861 2264
rect 8895 2292 8907 2295
rect 9784 2292 9812 2320
rect 9950 2292 9956 2304
rect 8895 2264 9812 2292
rect 9911 2264 9956 2292
rect 8895 2261 8907 2264
rect 8849 2255 8907 2261
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 10060 2292 10088 2332
rect 10226 2320 10232 2372
rect 10284 2360 10290 2372
rect 12345 2363 12403 2369
rect 12345 2360 12357 2363
rect 10284 2332 12357 2360
rect 10284 2320 10290 2332
rect 12345 2329 12357 2332
rect 12391 2360 12403 2363
rect 12618 2360 12624 2372
rect 12391 2332 12624 2360
rect 12391 2329 12403 2332
rect 12345 2323 12403 2329
rect 12618 2320 12624 2332
rect 12676 2320 12682 2372
rect 13446 2320 13452 2372
rect 13504 2360 13510 2372
rect 15657 2363 15715 2369
rect 15657 2360 15669 2363
rect 13504 2332 15669 2360
rect 13504 2320 13510 2332
rect 15657 2329 15669 2332
rect 15703 2329 15715 2363
rect 15657 2323 15715 2329
rect 10321 2295 10379 2301
rect 10321 2292 10333 2295
rect 10060 2264 10333 2292
rect 10321 2261 10333 2264
rect 10367 2292 10379 2295
rect 10686 2292 10692 2304
rect 10367 2264 10692 2292
rect 10367 2261 10379 2264
rect 10321 2255 10379 2261
rect 10686 2252 10692 2264
rect 10744 2252 10750 2304
rect 10873 2295 10931 2301
rect 10873 2261 10885 2295
rect 10919 2292 10931 2295
rect 11422 2292 11428 2304
rect 10919 2264 11428 2292
rect 10919 2261 10931 2264
rect 10873 2255 10931 2261
rect 11422 2252 11428 2264
rect 11480 2292 11486 2304
rect 13464 2292 13492 2320
rect 14642 2292 14648 2304
rect 11480 2264 13492 2292
rect 14603 2264 14648 2292
rect 11480 2252 11486 2264
rect 14642 2252 14648 2264
rect 14700 2252 14706 2304
rect 21376 2292 21404 2388
rect 22002 2320 22008 2372
rect 22060 2360 22066 2372
rect 23017 2363 23075 2369
rect 23017 2360 23029 2363
rect 22060 2332 23029 2360
rect 22060 2320 22066 2332
rect 23017 2329 23029 2332
rect 23063 2329 23075 2363
rect 23017 2323 23075 2329
rect 23106 2320 23112 2372
rect 23164 2360 23170 2372
rect 25731 2363 25789 2369
rect 25731 2360 25743 2363
rect 23164 2332 25743 2360
rect 23164 2320 23170 2332
rect 25731 2329 25743 2332
rect 25777 2329 25789 2363
rect 25731 2323 25789 2329
rect 26160 2301 26188 2468
rect 22649 2295 22707 2301
rect 22649 2292 22661 2295
rect 21376 2264 22661 2292
rect 22649 2261 22661 2264
rect 22695 2261 22707 2295
rect 22649 2255 22707 2261
rect 26145 2295 26203 2301
rect 26145 2261 26157 2295
rect 26191 2292 26203 2295
rect 27706 2292 27712 2304
rect 26191 2264 27712 2292
rect 26191 2261 26203 2264
rect 26145 2255 26203 2261
rect 27706 2252 27712 2264
rect 27764 2252 27770 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 15378 2048 15384 2100
rect 15436 2088 15442 2100
rect 23106 2088 23112 2100
rect 15436 2060 23112 2088
rect 15436 2048 15442 2060
rect 23106 2048 23112 2060
rect 23164 2048 23170 2100
rect 11974 76 11980 128
rect 12032 116 12038 128
rect 16298 116 16304 128
rect 12032 88 16304 116
rect 12032 76 12038 88
rect 16298 76 16304 88
rect 16356 76 16362 128
rect 16758 76 16764 128
rect 16816 116 16822 128
rect 17770 116 17776 128
rect 16816 88 17776 116
rect 16816 76 16822 88
rect 17770 76 17776 88
rect 17828 76 17834 128
<< via1 >>
rect 5540 27480 5592 27532
rect 6184 27480 6236 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 18328 24828 18380 24880
rect 27620 24828 27672 24880
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 20168 24352 20220 24404
rect 10692 24259 10744 24268
rect 10692 24225 10710 24259
rect 10710 24225 10744 24259
rect 10692 24216 10744 24225
rect 11520 24216 11572 24268
rect 11704 24216 11756 24268
rect 16948 24259 17000 24268
rect 16948 24225 16957 24259
rect 16957 24225 16991 24259
rect 16991 24225 17000 24259
rect 16948 24216 17000 24225
rect 18052 24259 18104 24268
rect 18052 24225 18061 24259
rect 18061 24225 18095 24259
rect 18095 24225 18104 24259
rect 18052 24216 18104 24225
rect 18788 24080 18840 24132
rect 9772 24012 9824 24064
rect 11336 24012 11388 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 10692 23851 10744 23860
rect 10692 23817 10701 23851
rect 10701 23817 10735 23851
rect 10735 23817 10744 23851
rect 10692 23808 10744 23817
rect 16028 23808 16080 23860
rect 17408 23808 17460 23860
rect 18052 23808 18104 23860
rect 18512 23808 18564 23860
rect 21640 23808 21692 23860
rect 24216 23808 24268 23860
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 22652 23740 22704 23792
rect 24216 23672 24268 23724
rect 27160 23672 27212 23724
rect 1952 23647 2004 23656
rect 1952 23613 1961 23647
rect 1961 23613 1995 23647
rect 1995 23613 2004 23647
rect 1952 23604 2004 23613
rect 7196 23604 7248 23656
rect 11244 23604 11296 23656
rect 11520 23604 11572 23656
rect 14372 23647 14424 23656
rect 14372 23613 14381 23647
rect 14381 23613 14415 23647
rect 14415 23613 14424 23647
rect 14372 23604 14424 23613
rect 12992 23536 13044 23588
rect 18144 23604 18196 23656
rect 21272 23647 21324 23656
rect 15292 23536 15344 23588
rect 16948 23579 17000 23588
rect 16948 23545 16957 23579
rect 16957 23545 16991 23579
rect 16991 23545 17000 23579
rect 16948 23536 17000 23545
rect 5264 23468 5316 23520
rect 9956 23511 10008 23520
rect 9956 23477 9965 23511
rect 9965 23477 9999 23511
rect 9999 23477 10008 23511
rect 9956 23468 10008 23477
rect 10692 23468 10744 23520
rect 11704 23511 11756 23520
rect 11704 23477 11713 23511
rect 11713 23477 11747 23511
rect 11747 23477 11756 23511
rect 11704 23468 11756 23477
rect 12256 23468 12308 23520
rect 12716 23468 12768 23520
rect 18236 23511 18288 23520
rect 18236 23477 18245 23511
rect 18245 23477 18279 23511
rect 18279 23477 18288 23511
rect 18236 23468 18288 23477
rect 21272 23613 21281 23647
rect 21281 23613 21315 23647
rect 21315 23613 21324 23647
rect 21272 23604 21324 23613
rect 21916 23604 21968 23656
rect 21088 23468 21140 23520
rect 22376 23468 22428 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1124 23264 1176 23316
rect 11152 23307 11204 23316
rect 11152 23273 11161 23307
rect 11161 23273 11195 23307
rect 11195 23273 11204 23307
rect 11152 23264 11204 23273
rect 13176 23264 13228 23316
rect 14372 23264 14424 23316
rect 18328 23264 18380 23316
rect 24860 23264 24912 23316
rect 1952 23196 2004 23248
rect 8576 23196 8628 23248
rect 9864 23239 9916 23248
rect 9864 23205 9873 23239
rect 9873 23205 9907 23239
rect 9907 23205 9916 23239
rect 9864 23196 9916 23205
rect 14648 23196 14700 23248
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 7196 23128 7248 23180
rect 11336 23128 11388 23180
rect 12164 23128 12216 23180
rect 13820 23128 13872 23180
rect 15384 23171 15436 23180
rect 15384 23137 15393 23171
rect 15393 23137 15427 23171
rect 15427 23137 15436 23171
rect 15384 23128 15436 23137
rect 16764 23171 16816 23180
rect 16764 23137 16808 23171
rect 16808 23137 16816 23171
rect 18052 23171 18104 23180
rect 16764 23128 16816 23137
rect 18052 23137 18061 23171
rect 18061 23137 18095 23171
rect 18095 23137 18104 23171
rect 18052 23128 18104 23137
rect 24676 23128 24728 23180
rect 9220 23060 9272 23112
rect 10048 23103 10100 23112
rect 10048 23069 10057 23103
rect 10057 23069 10091 23103
rect 10091 23069 10100 23103
rect 10048 23060 10100 23069
rect 6276 22992 6328 23044
rect 12992 22992 13044 23044
rect 7288 22924 7340 22976
rect 7748 22967 7800 22976
rect 7748 22933 7757 22967
rect 7757 22933 7791 22967
rect 7791 22933 7800 22967
rect 7748 22924 7800 22933
rect 8852 22924 8904 22976
rect 11060 22924 11112 22976
rect 12532 22924 12584 22976
rect 15936 22924 15988 22976
rect 17592 22924 17644 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1216 22720 1268 22772
rect 7196 22763 7248 22772
rect 7196 22729 7205 22763
rect 7205 22729 7239 22763
rect 7239 22729 7248 22763
rect 7196 22720 7248 22729
rect 8208 22720 8260 22772
rect 8576 22763 8628 22772
rect 8576 22729 8585 22763
rect 8585 22729 8619 22763
rect 8619 22729 8628 22763
rect 8576 22720 8628 22729
rect 9864 22720 9916 22772
rect 11520 22720 11572 22772
rect 13084 22720 13136 22772
rect 1032 22584 1084 22636
rect 7748 22652 7800 22704
rect 9220 22652 9272 22704
rect 11336 22695 11388 22704
rect 11336 22661 11345 22695
rect 11345 22661 11379 22695
rect 11379 22661 11388 22695
rect 11336 22652 11388 22661
rect 13452 22652 13504 22704
rect 1952 22559 2004 22568
rect 1952 22525 1961 22559
rect 1961 22525 1995 22559
rect 1995 22525 2004 22559
rect 1952 22516 2004 22525
rect 7564 22584 7616 22636
rect 9588 22627 9640 22636
rect 9588 22593 9597 22627
rect 9597 22593 9631 22627
rect 9631 22593 9640 22627
rect 9588 22584 9640 22593
rect 10048 22584 10100 22636
rect 13820 22584 13872 22636
rect 10876 22559 10928 22568
rect 10876 22525 10894 22559
rect 10894 22525 10928 22559
rect 10876 22516 10928 22525
rect 12164 22516 12216 22568
rect 12440 22559 12492 22568
rect 6460 22448 6512 22500
rect 7104 22380 7156 22432
rect 7748 22448 7800 22500
rect 9312 22491 9364 22500
rect 9312 22457 9321 22491
rect 9321 22457 9355 22491
rect 9355 22457 9364 22491
rect 9312 22448 9364 22457
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 12440 22516 12492 22525
rect 14004 22559 14056 22568
rect 14004 22525 14013 22559
rect 14013 22525 14047 22559
rect 14047 22525 14056 22559
rect 14004 22516 14056 22525
rect 16764 22763 16816 22772
rect 16764 22729 16773 22763
rect 16773 22729 16807 22763
rect 16807 22729 16816 22763
rect 16764 22720 16816 22729
rect 18052 22652 18104 22704
rect 16856 22516 16908 22568
rect 9036 22423 9088 22432
rect 9036 22389 9045 22423
rect 9045 22389 9079 22423
rect 9079 22389 9088 22423
rect 13728 22448 13780 22500
rect 15384 22448 15436 22500
rect 22376 22448 22428 22500
rect 9036 22380 9088 22389
rect 10784 22380 10836 22432
rect 12624 22423 12676 22432
rect 12624 22389 12633 22423
rect 12633 22389 12667 22423
rect 12667 22389 12676 22423
rect 12624 22380 12676 22389
rect 13360 22380 13412 22432
rect 15660 22423 15712 22432
rect 15660 22389 15669 22423
rect 15669 22389 15703 22423
rect 15703 22389 15712 22423
rect 15660 22380 15712 22389
rect 23480 22380 23532 22432
rect 24676 22380 24728 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1400 22176 1452 22228
rect 8852 22219 8904 22228
rect 8852 22185 8861 22219
rect 8861 22185 8895 22219
rect 8895 22185 8904 22219
rect 8852 22176 8904 22185
rect 11060 22219 11112 22228
rect 11060 22185 11069 22219
rect 11069 22185 11103 22219
rect 11103 22185 11112 22219
rect 11060 22176 11112 22185
rect 12532 22176 12584 22228
rect 6828 22108 6880 22160
rect 10140 22151 10192 22160
rect 10140 22117 10149 22151
rect 10149 22117 10183 22151
rect 10183 22117 10192 22151
rect 10140 22108 10192 22117
rect 13452 22176 13504 22228
rect 15292 22176 15344 22228
rect 13268 22151 13320 22160
rect 13268 22117 13277 22151
rect 13277 22117 13311 22151
rect 13311 22117 13320 22151
rect 13268 22108 13320 22117
rect 15752 22108 15804 22160
rect 6184 22083 6236 22092
rect 6184 22049 6193 22083
rect 6193 22049 6227 22083
rect 6227 22049 6236 22083
rect 6184 22040 6236 22049
rect 11520 22083 11572 22092
rect 11520 22049 11529 22083
rect 11529 22049 11563 22083
rect 11563 22049 11572 22083
rect 11520 22040 11572 22049
rect 6644 21972 6696 22024
rect 7380 21972 7432 22024
rect 7564 22015 7616 22024
rect 7564 21981 7573 22015
rect 7573 21981 7607 22015
rect 7607 21981 7616 22015
rect 7564 21972 7616 21981
rect 9496 21972 9548 22024
rect 10784 21972 10836 22024
rect 16948 21972 17000 22024
rect 8668 21904 8720 21956
rect 9588 21904 9640 21956
rect 13728 21947 13780 21956
rect 13728 21913 13737 21947
rect 13737 21913 13771 21947
rect 13771 21913 13780 21947
rect 13728 21904 13780 21913
rect 16488 21904 16540 21956
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 12808 21879 12860 21888
rect 12808 21845 12817 21879
rect 12817 21845 12851 21879
rect 12851 21845 12860 21879
rect 12808 21836 12860 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 7656 21632 7708 21684
rect 11520 21675 11572 21684
rect 11520 21641 11529 21675
rect 11529 21641 11563 21675
rect 11563 21641 11572 21675
rect 11520 21632 11572 21641
rect 13268 21632 13320 21684
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 7012 21564 7064 21616
rect 6184 21496 6236 21548
rect 7564 21539 7616 21548
rect 7564 21505 7573 21539
rect 7573 21505 7607 21539
rect 7607 21505 7616 21539
rect 7564 21496 7616 21505
rect 7840 21564 7892 21616
rect 8668 21496 8720 21548
rect 8852 21539 8904 21548
rect 8852 21505 8861 21539
rect 8861 21505 8895 21539
rect 8895 21505 8904 21539
rect 8852 21496 8904 21505
rect 9128 21539 9180 21548
rect 9128 21505 9137 21539
rect 9137 21505 9171 21539
rect 9171 21505 9180 21539
rect 9128 21496 9180 21505
rect 11060 21496 11112 21548
rect 13360 21564 13412 21616
rect 13544 21564 13596 21616
rect 13728 21496 13780 21548
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 16856 21564 16908 21616
rect 15752 21496 15804 21548
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 664 21428 716 21480
rect 4988 21428 5040 21480
rect 6276 21471 6328 21480
rect 6276 21437 6285 21471
rect 6285 21437 6319 21471
rect 6319 21437 6328 21471
rect 6276 21428 6328 21437
rect 18144 21471 18196 21480
rect 18144 21437 18162 21471
rect 18162 21437 18196 21471
rect 18144 21428 18196 21437
rect 22008 21428 22060 21480
rect 25136 21471 25188 21480
rect 25136 21437 25145 21471
rect 25145 21437 25179 21471
rect 25179 21437 25188 21471
rect 25136 21428 25188 21437
rect 6920 21360 6972 21412
rect 7012 21360 7064 21412
rect 7380 21403 7432 21412
rect 7380 21369 7389 21403
rect 7389 21369 7423 21403
rect 7423 21369 7432 21403
rect 7380 21360 7432 21369
rect 5080 21335 5132 21344
rect 5080 21301 5089 21335
rect 5089 21301 5123 21335
rect 5123 21301 5132 21335
rect 5080 21292 5132 21301
rect 6828 21292 6880 21344
rect 7196 21292 7248 21344
rect 8576 21335 8628 21344
rect 8576 21301 8585 21335
rect 8585 21301 8619 21335
rect 8619 21301 8628 21335
rect 9036 21360 9088 21412
rect 12808 21360 12860 21412
rect 13544 21360 13596 21412
rect 16028 21403 16080 21412
rect 8576 21292 8628 21301
rect 10140 21335 10192 21344
rect 10140 21301 10149 21335
rect 10149 21301 10183 21335
rect 10183 21301 10192 21335
rect 10140 21292 10192 21301
rect 14188 21335 14240 21344
rect 14188 21301 14197 21335
rect 14197 21301 14231 21335
rect 14231 21301 14240 21335
rect 14188 21292 14240 21301
rect 14556 21292 14608 21344
rect 16028 21369 16037 21403
rect 16037 21369 16071 21403
rect 16071 21369 16080 21403
rect 16028 21360 16080 21369
rect 16396 21360 16448 21412
rect 16948 21335 17000 21344
rect 16948 21301 16957 21335
rect 16957 21301 16991 21335
rect 16991 21301 17000 21335
rect 16948 21292 17000 21301
rect 17500 21292 17552 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 5264 21131 5316 21140
rect 5264 21097 5273 21131
rect 5273 21097 5307 21131
rect 5307 21097 5316 21131
rect 5264 21088 5316 21097
rect 6552 21088 6604 21140
rect 7196 21088 7248 21140
rect 7380 21131 7432 21140
rect 7380 21097 7389 21131
rect 7389 21097 7423 21131
rect 7423 21097 7432 21131
rect 7380 21088 7432 21097
rect 7472 21088 7524 21140
rect 2044 21020 2096 21072
rect 9220 21088 9272 21140
rect 9496 21131 9548 21140
rect 9496 21097 9505 21131
rect 9505 21097 9539 21131
rect 9539 21097 9548 21131
rect 9496 21088 9548 21097
rect 13268 21088 13320 21140
rect 13912 21088 13964 21140
rect 15844 21088 15896 21140
rect 4436 20995 4488 21004
rect 4436 20961 4445 20995
rect 4445 20961 4479 20995
rect 4479 20961 4488 20995
rect 4436 20952 4488 20961
rect 5080 20952 5132 21004
rect 6184 20952 6236 21004
rect 8484 20952 8536 21004
rect 4620 20791 4672 20800
rect 4620 20757 4629 20791
rect 4629 20757 4663 20791
rect 4663 20757 4672 20791
rect 4620 20748 4672 20757
rect 6000 20748 6052 20800
rect 6276 20791 6328 20800
rect 6276 20757 6285 20791
rect 6285 20757 6319 20791
rect 6319 20757 6328 20791
rect 9496 20884 9548 20936
rect 9864 21020 9916 21072
rect 11152 21020 11204 21072
rect 13728 21063 13780 21072
rect 13728 21029 13737 21063
rect 13737 21029 13771 21063
rect 13771 21029 13780 21063
rect 13728 21020 13780 21029
rect 13820 21063 13872 21072
rect 13820 21029 13829 21063
rect 13829 21029 13863 21063
rect 13863 21029 13872 21063
rect 14372 21063 14424 21072
rect 13820 21020 13872 21029
rect 14372 21029 14381 21063
rect 14381 21029 14415 21063
rect 14415 21029 14424 21063
rect 14372 21020 14424 21029
rect 15660 21020 15712 21072
rect 17408 21088 17460 21140
rect 17500 21063 17552 21072
rect 17500 21029 17509 21063
rect 17509 21029 17543 21063
rect 17543 21029 17552 21063
rect 17500 21020 17552 21029
rect 12072 20995 12124 21004
rect 12072 20961 12081 20995
rect 12081 20961 12115 20995
rect 12115 20961 12124 20995
rect 12072 20952 12124 20961
rect 12532 20995 12584 21004
rect 12532 20961 12541 20995
rect 12541 20961 12575 20995
rect 12575 20961 12584 20995
rect 12532 20952 12584 20961
rect 9680 20884 9732 20936
rect 10784 20884 10836 20936
rect 13268 20927 13320 20936
rect 13268 20893 13277 20927
rect 13277 20893 13311 20927
rect 13311 20893 13320 20927
rect 13268 20884 13320 20893
rect 16396 20927 16448 20936
rect 16396 20893 16405 20927
rect 16405 20893 16439 20927
rect 16439 20893 16448 20927
rect 16396 20884 16448 20893
rect 10600 20816 10652 20868
rect 16488 20816 16540 20868
rect 7656 20791 7708 20800
rect 6276 20748 6328 20757
rect 7656 20757 7665 20791
rect 7665 20757 7699 20791
rect 7699 20757 7708 20791
rect 7656 20748 7708 20757
rect 9036 20791 9088 20800
rect 9036 20757 9045 20791
rect 9045 20757 9079 20791
rect 9079 20757 9088 20791
rect 9036 20748 9088 20757
rect 10140 20791 10192 20800
rect 10140 20757 10149 20791
rect 10149 20757 10183 20791
rect 10183 20757 10192 20791
rect 10140 20748 10192 20757
rect 16304 20748 16356 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1860 20408 1912 20460
rect 1400 20204 1452 20256
rect 5540 20544 5592 20596
rect 7748 20587 7800 20596
rect 7748 20553 7757 20587
rect 7757 20553 7791 20587
rect 7791 20553 7800 20587
rect 7748 20544 7800 20553
rect 8484 20587 8536 20596
rect 8484 20553 8493 20587
rect 8493 20553 8527 20587
rect 8527 20553 8536 20587
rect 8484 20544 8536 20553
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 9956 20587 10008 20596
rect 9956 20553 9965 20587
rect 9965 20553 9999 20587
rect 9999 20553 10008 20587
rect 11152 20587 11204 20596
rect 9956 20544 10008 20553
rect 3976 20476 4028 20528
rect 4436 20476 4488 20528
rect 4896 20476 4948 20528
rect 8944 20476 8996 20528
rect 9036 20408 9088 20460
rect 9128 20451 9180 20460
rect 9128 20417 9137 20451
rect 9137 20417 9171 20451
rect 9171 20417 9180 20451
rect 11152 20553 11161 20587
rect 11161 20553 11195 20587
rect 11195 20553 11204 20587
rect 11152 20544 11204 20553
rect 12072 20587 12124 20596
rect 12072 20553 12081 20587
rect 12081 20553 12115 20587
rect 12115 20553 12124 20587
rect 12072 20544 12124 20553
rect 12532 20544 12584 20596
rect 14188 20587 14240 20596
rect 14188 20553 14197 20587
rect 14197 20553 14231 20587
rect 14231 20553 14240 20587
rect 14188 20544 14240 20553
rect 15660 20544 15712 20596
rect 16028 20544 16080 20596
rect 17408 20587 17460 20596
rect 17408 20553 17417 20587
rect 17417 20553 17451 20587
rect 17451 20553 17460 20587
rect 17408 20544 17460 20553
rect 17500 20544 17552 20596
rect 16948 20476 17000 20528
rect 9128 20408 9180 20417
rect 10600 20451 10652 20460
rect 10600 20417 10609 20451
rect 10609 20417 10643 20451
rect 10643 20417 10652 20451
rect 10600 20408 10652 20417
rect 10876 20408 10928 20460
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 16488 20408 16540 20460
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 5080 20383 5132 20392
rect 5080 20349 5089 20383
rect 5089 20349 5123 20383
rect 5123 20349 5132 20383
rect 5080 20340 5132 20349
rect 5264 20340 5316 20392
rect 6092 20340 6144 20392
rect 7656 20340 7708 20392
rect 14556 20340 14608 20392
rect 15568 20340 15620 20392
rect 18512 20408 18564 20460
rect 20352 20408 20404 20460
rect 19524 20383 19576 20392
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 7012 20272 7064 20324
rect 2504 20204 2556 20256
rect 3516 20204 3568 20256
rect 3792 20204 3844 20256
rect 6184 20247 6236 20256
rect 6184 20213 6193 20247
rect 6193 20213 6227 20247
rect 6227 20213 6236 20247
rect 6184 20204 6236 20213
rect 6552 20247 6604 20256
rect 6552 20213 6561 20247
rect 6561 20213 6595 20247
rect 6595 20213 6604 20247
rect 9128 20272 9180 20324
rect 6552 20204 6604 20213
rect 10140 20204 10192 20256
rect 13176 20247 13228 20256
rect 13176 20213 13185 20247
rect 13185 20213 13219 20247
rect 13219 20213 13228 20247
rect 16304 20315 16356 20324
rect 16304 20281 16313 20315
rect 16313 20281 16347 20315
rect 16347 20281 16356 20315
rect 16304 20272 16356 20281
rect 14464 20247 14516 20256
rect 13176 20204 13228 20213
rect 14464 20213 14473 20247
rect 14473 20213 14507 20247
rect 14507 20213 14516 20247
rect 14464 20204 14516 20213
rect 15384 20204 15436 20256
rect 15568 20247 15620 20256
rect 15568 20213 15577 20247
rect 15577 20213 15611 20247
rect 15611 20213 15620 20247
rect 15568 20204 15620 20213
rect 18052 20204 18104 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 6828 20000 6880 20052
rect 9036 20000 9088 20052
rect 9128 20043 9180 20052
rect 9128 20009 9137 20043
rect 9137 20009 9171 20043
rect 9171 20009 9180 20043
rect 9128 20000 9180 20009
rect 9864 20000 9916 20052
rect 10784 20000 10836 20052
rect 13176 20000 13228 20052
rect 13728 20000 13780 20052
rect 15844 20043 15896 20052
rect 15844 20009 15853 20043
rect 15853 20009 15887 20043
rect 15887 20009 15896 20043
rect 15844 20000 15896 20009
rect 6276 19932 6328 19984
rect 6552 19932 6604 19984
rect 9588 19932 9640 19984
rect 15752 19932 15804 19984
rect 16212 19975 16264 19984
rect 16212 19941 16221 19975
rect 16221 19941 16255 19975
rect 16255 19941 16264 19975
rect 16212 19932 16264 19941
rect 16856 19932 16908 19984
rect 17776 19975 17828 19984
rect 17776 19941 17785 19975
rect 17785 19941 17819 19975
rect 17819 19941 17828 19975
rect 17776 19932 17828 19941
rect 1492 19864 1544 19916
rect 2688 19864 2740 19916
rect 4620 19864 4672 19916
rect 5264 19907 5316 19916
rect 4712 19796 4764 19848
rect 5264 19873 5273 19907
rect 5273 19873 5307 19907
rect 5307 19873 5316 19907
rect 5264 19864 5316 19873
rect 5448 19864 5500 19916
rect 8944 19864 8996 19916
rect 11888 19864 11940 19916
rect 13820 19907 13872 19916
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 14464 19864 14516 19916
rect 18880 19864 18932 19916
rect 6368 19839 6420 19848
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 7012 19796 7064 19848
rect 10600 19796 10652 19848
rect 12808 19796 12860 19848
rect 16396 19796 16448 19848
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 17960 19839 18012 19848
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 12072 19728 12124 19780
rect 1676 19660 1728 19712
rect 2412 19660 2464 19712
rect 7748 19703 7800 19712
rect 7748 19669 7757 19703
rect 7757 19669 7791 19703
rect 7791 19669 7800 19703
rect 7748 19660 7800 19669
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 16580 19660 16632 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 4712 19499 4764 19508
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 10140 19456 10192 19508
rect 10600 19456 10652 19508
rect 16212 19499 16264 19508
rect 16212 19465 16221 19499
rect 16221 19465 16255 19499
rect 16255 19465 16264 19499
rect 16212 19456 16264 19465
rect 16396 19456 16448 19508
rect 17960 19456 18012 19508
rect 24768 19499 24820 19508
rect 8576 19388 8628 19440
rect 6368 19320 6420 19372
rect 11336 19388 11388 19440
rect 12440 19388 12492 19440
rect 17776 19388 17828 19440
rect 10140 19320 10192 19372
rect 2044 19227 2096 19236
rect 2044 19193 2053 19227
rect 2053 19193 2087 19227
rect 2087 19193 2096 19227
rect 2044 19184 2096 19193
rect 3424 19252 3476 19304
rect 4068 19295 4120 19304
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 5264 19295 5316 19304
rect 5264 19261 5273 19295
rect 5273 19261 5307 19295
rect 5307 19261 5316 19295
rect 5264 19252 5316 19261
rect 5448 19252 5500 19304
rect 7748 19295 7800 19304
rect 7748 19261 7757 19295
rect 7757 19261 7791 19295
rect 7791 19261 7800 19295
rect 7748 19252 7800 19261
rect 4252 19184 4304 19236
rect 9404 19252 9456 19304
rect 8944 19227 8996 19236
rect 8944 19193 8953 19227
rect 8953 19193 8987 19227
rect 8987 19193 8996 19227
rect 8944 19184 8996 19193
rect 2596 19116 2648 19168
rect 3240 19116 3292 19168
rect 3424 19159 3476 19168
rect 3424 19125 3433 19159
rect 3433 19125 3467 19159
rect 3467 19125 3476 19159
rect 3424 19116 3476 19125
rect 6368 19159 6420 19168
rect 6368 19125 6377 19159
rect 6377 19125 6411 19159
rect 6411 19125 6420 19159
rect 6368 19116 6420 19125
rect 6552 19116 6604 19168
rect 7932 19116 7984 19168
rect 8024 19116 8076 19168
rect 9588 19116 9640 19168
rect 11152 19159 11204 19168
rect 11152 19125 11161 19159
rect 11161 19125 11195 19159
rect 11195 19125 11204 19159
rect 11152 19116 11204 19125
rect 11888 19159 11940 19168
rect 11888 19125 11897 19159
rect 11897 19125 11931 19159
rect 11931 19125 11940 19159
rect 11888 19116 11940 19125
rect 13820 19320 13872 19372
rect 24768 19465 24777 19499
rect 24777 19465 24811 19499
rect 24811 19465 24820 19499
rect 24768 19456 24820 19465
rect 12532 19295 12584 19304
rect 12532 19261 12541 19295
rect 12541 19261 12575 19295
rect 12575 19261 12584 19295
rect 12532 19252 12584 19261
rect 12808 19252 12860 19304
rect 13268 19252 13320 19304
rect 13912 19252 13964 19304
rect 14740 19252 14792 19304
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 17316 19252 17368 19304
rect 18972 19252 19024 19304
rect 19432 19252 19484 19304
rect 20536 19252 20588 19304
rect 23112 19252 23164 19304
rect 13176 19184 13228 19236
rect 13268 19116 13320 19168
rect 17684 19184 17736 19236
rect 18880 19184 18932 19236
rect 17776 19116 17828 19168
rect 19064 19116 19116 19168
rect 19432 19116 19484 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 4252 18912 4304 18964
rect 9404 18955 9456 18964
rect 9404 18921 9413 18955
rect 9413 18921 9447 18955
rect 9447 18921 9456 18955
rect 9404 18912 9456 18921
rect 12440 18955 12492 18964
rect 12440 18921 12449 18955
rect 12449 18921 12483 18955
rect 12483 18921 12492 18955
rect 12440 18912 12492 18921
rect 13176 18955 13228 18964
rect 13176 18921 13185 18955
rect 13185 18921 13219 18955
rect 13219 18921 13228 18955
rect 13176 18912 13228 18921
rect 13544 18912 13596 18964
rect 16304 18912 16356 18964
rect 16580 18955 16632 18964
rect 16580 18921 16589 18955
rect 16589 18921 16623 18955
rect 16623 18921 16632 18955
rect 16580 18912 16632 18921
rect 17132 18955 17184 18964
rect 17132 18921 17141 18955
rect 17141 18921 17175 18955
rect 17175 18921 17184 18955
rect 17132 18912 17184 18921
rect 17684 18912 17736 18964
rect 24216 18912 24268 18964
rect 6092 18887 6144 18896
rect 1952 18776 2004 18828
rect 2964 18819 3016 18828
rect 2964 18785 3008 18819
rect 3008 18785 3016 18819
rect 2964 18776 3016 18785
rect 3700 18708 3752 18760
rect 4528 18640 4580 18692
rect 1492 18572 1544 18624
rect 3608 18572 3660 18624
rect 4068 18572 4120 18624
rect 6092 18853 6101 18887
rect 6101 18853 6135 18887
rect 6135 18853 6144 18887
rect 6092 18844 6144 18853
rect 10232 18844 10284 18896
rect 10876 18887 10928 18896
rect 10876 18853 10885 18887
rect 10885 18853 10919 18887
rect 10919 18853 10928 18887
rect 10876 18844 10928 18853
rect 15476 18844 15528 18896
rect 5356 18819 5408 18828
rect 5356 18785 5365 18819
rect 5365 18785 5399 18819
rect 5399 18785 5408 18819
rect 5356 18776 5408 18785
rect 5448 18776 5500 18828
rect 7012 18819 7064 18828
rect 7012 18785 7021 18819
rect 7021 18785 7055 18819
rect 7055 18785 7064 18819
rect 7012 18776 7064 18785
rect 7196 18776 7248 18828
rect 11796 18776 11848 18828
rect 11888 18776 11940 18828
rect 17040 18819 17092 18828
rect 8024 18708 8076 18760
rect 8668 18708 8720 18760
rect 5080 18640 5132 18692
rect 9036 18640 9088 18692
rect 13176 18708 13228 18760
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 17040 18785 17049 18819
rect 17049 18785 17083 18819
rect 17083 18785 17092 18819
rect 17040 18776 17092 18785
rect 17408 18776 17460 18828
rect 18788 18776 18840 18828
rect 18972 18776 19024 18828
rect 20076 18776 20128 18828
rect 24124 18776 24176 18828
rect 18512 18708 18564 18760
rect 20444 18708 20496 18760
rect 17776 18640 17828 18692
rect 18420 18640 18472 18692
rect 5264 18615 5316 18624
rect 5264 18581 5273 18615
rect 5273 18581 5307 18615
rect 5307 18581 5316 18615
rect 5264 18572 5316 18581
rect 8300 18572 8352 18624
rect 9220 18572 9272 18624
rect 9588 18572 9640 18624
rect 12164 18572 12216 18624
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 14740 18572 14792 18624
rect 18604 18572 18656 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1952 18368 2004 18420
rect 4896 18368 4948 18420
rect 5172 18368 5224 18420
rect 7012 18411 7064 18420
rect 7012 18377 7021 18411
rect 7021 18377 7055 18411
rect 7055 18377 7064 18411
rect 7012 18368 7064 18377
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 13268 18368 13320 18420
rect 13912 18368 13964 18420
rect 17040 18411 17092 18420
rect 2964 18300 3016 18352
rect 4436 18300 4488 18352
rect 7196 18300 7248 18352
rect 12440 18300 12492 18352
rect 1952 18028 2004 18080
rect 2964 18028 3016 18080
rect 7748 18232 7800 18284
rect 8116 18232 8168 18284
rect 12808 18232 12860 18284
rect 14740 18275 14792 18284
rect 4068 18207 4120 18216
rect 4068 18173 4077 18207
rect 4077 18173 4111 18207
rect 4111 18173 4120 18207
rect 4068 18164 4120 18173
rect 5172 18207 5224 18216
rect 5172 18173 5181 18207
rect 5181 18173 5215 18207
rect 5215 18173 5224 18207
rect 5172 18164 5224 18173
rect 5264 18164 5316 18216
rect 6092 18164 6144 18216
rect 9036 18164 9088 18216
rect 9680 18207 9732 18216
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 11336 18207 11388 18216
rect 5448 18096 5500 18148
rect 6736 18096 6788 18148
rect 4436 18028 4488 18080
rect 6552 18028 6604 18080
rect 7472 18139 7524 18148
rect 7472 18105 7481 18139
rect 7481 18105 7515 18139
rect 7515 18105 7524 18139
rect 9956 18139 10008 18148
rect 7472 18096 7524 18105
rect 9956 18105 9965 18139
rect 9965 18105 9999 18139
rect 9999 18105 10008 18139
rect 9956 18096 10008 18105
rect 8300 18028 8352 18080
rect 8668 18071 8720 18080
rect 8668 18037 8677 18071
rect 8677 18037 8711 18071
rect 8711 18037 8720 18071
rect 8668 18028 8720 18037
rect 11336 18173 11345 18207
rect 11345 18173 11379 18207
rect 11379 18173 11388 18207
rect 11336 18164 11388 18173
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 13176 18139 13228 18148
rect 13176 18105 13185 18139
rect 13185 18105 13219 18139
rect 13219 18105 13228 18139
rect 13176 18096 13228 18105
rect 11336 18028 11388 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 13544 18028 13596 18080
rect 14096 18164 14148 18216
rect 17040 18377 17049 18411
rect 17049 18377 17083 18411
rect 17083 18377 17092 18411
rect 17040 18368 17092 18377
rect 18788 18368 18840 18420
rect 19524 18368 19576 18420
rect 20076 18411 20128 18420
rect 20076 18377 20085 18411
rect 20085 18377 20119 18411
rect 20119 18377 20128 18411
rect 20076 18368 20128 18377
rect 16580 18300 16632 18352
rect 16488 18275 16540 18284
rect 16488 18241 16497 18275
rect 16497 18241 16531 18275
rect 16531 18241 16540 18275
rect 16488 18232 16540 18241
rect 16672 18232 16724 18284
rect 18788 18164 18840 18216
rect 20536 18164 20588 18216
rect 17960 18096 18012 18148
rect 15476 18028 15528 18080
rect 17408 18071 17460 18080
rect 17408 18037 17417 18071
rect 17417 18037 17451 18071
rect 17451 18037 17460 18071
rect 17408 18028 17460 18037
rect 18972 18028 19024 18080
rect 20628 18071 20680 18080
rect 20628 18037 20637 18071
rect 20637 18037 20671 18071
rect 20671 18037 20680 18071
rect 20628 18028 20680 18037
rect 21180 18028 21232 18080
rect 24124 18028 24176 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 4068 17824 4120 17876
rect 6368 17867 6420 17876
rect 6368 17833 6377 17867
rect 6377 17833 6411 17867
rect 6411 17833 6420 17867
rect 6368 17824 6420 17833
rect 7472 17824 7524 17876
rect 10140 17867 10192 17876
rect 10140 17833 10149 17867
rect 10149 17833 10183 17867
rect 10183 17833 10192 17867
rect 10140 17824 10192 17833
rect 13176 17824 13228 17876
rect 16120 17824 16172 17876
rect 5172 17756 5224 17808
rect 7932 17799 7984 17808
rect 7932 17765 7941 17799
rect 7941 17765 7975 17799
rect 7975 17765 7984 17799
rect 7932 17756 7984 17765
rect 8116 17756 8168 17808
rect 10784 17756 10836 17808
rect 15292 17756 15344 17808
rect 16856 17799 16908 17808
rect 16856 17765 16865 17799
rect 16865 17765 16899 17799
rect 16899 17765 16908 17799
rect 16856 17756 16908 17765
rect 17408 17756 17460 17808
rect 2320 17688 2372 17740
rect 4712 17731 4764 17740
rect 4712 17697 4721 17731
rect 4721 17697 4755 17731
rect 4755 17697 4764 17731
rect 4712 17688 4764 17697
rect 5356 17688 5408 17740
rect 6552 17688 6604 17740
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 12440 17731 12492 17740
rect 12440 17697 12449 17731
rect 12449 17697 12483 17731
rect 12483 17697 12492 17731
rect 12440 17688 12492 17697
rect 14096 17731 14148 17740
rect 3332 17620 3384 17672
rect 6828 17620 6880 17672
rect 8668 17620 8720 17672
rect 10692 17620 10744 17672
rect 12532 17663 12584 17672
rect 8300 17552 8352 17604
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 14096 17697 14105 17731
rect 14105 17697 14139 17731
rect 14139 17697 14148 17731
rect 14096 17688 14148 17697
rect 15936 17688 15988 17740
rect 16672 17688 16724 17740
rect 17132 17688 17184 17740
rect 18696 17688 18748 17740
rect 13912 17620 13964 17672
rect 16764 17620 16816 17672
rect 17040 17620 17092 17672
rect 17224 17620 17276 17672
rect 20996 17688 21048 17740
rect 22560 17688 22612 17740
rect 23572 17688 23624 17740
rect 11704 17552 11756 17604
rect 19248 17552 19300 17604
rect 1768 17484 1820 17536
rect 4804 17484 4856 17536
rect 9680 17484 9732 17536
rect 10140 17484 10192 17536
rect 14372 17484 14424 17536
rect 15568 17484 15620 17536
rect 17224 17484 17276 17536
rect 17500 17527 17552 17536
rect 17500 17493 17509 17527
rect 17509 17493 17543 17527
rect 17543 17493 17552 17527
rect 17500 17484 17552 17493
rect 18236 17484 18288 17536
rect 20260 17484 20312 17536
rect 21732 17484 21784 17536
rect 22468 17484 22520 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 4712 17280 4764 17332
rect 7932 17280 7984 17332
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 12440 17280 12492 17332
rect 13268 17280 13320 17332
rect 13912 17323 13964 17332
rect 6184 17212 6236 17264
rect 2964 17144 3016 17196
rect 4160 17119 4212 17128
rect 4160 17085 4169 17119
rect 4169 17085 4203 17119
rect 4203 17085 4212 17119
rect 4160 17076 4212 17085
rect 4344 17008 4396 17060
rect 6552 17144 6604 17196
rect 6736 17144 6788 17196
rect 13912 17289 13921 17323
rect 13921 17289 13955 17323
rect 13955 17289 13964 17323
rect 13912 17280 13964 17289
rect 17408 17280 17460 17332
rect 24768 17323 24820 17332
rect 24768 17289 24777 17323
rect 24777 17289 24811 17323
rect 24811 17289 24820 17323
rect 24768 17280 24820 17289
rect 18236 17212 18288 17264
rect 18512 17212 18564 17264
rect 11244 17144 11296 17196
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 16120 17187 16172 17196
rect 16120 17153 16129 17187
rect 16129 17153 16163 17187
rect 16163 17153 16172 17187
rect 16120 17144 16172 17153
rect 18328 17144 18380 17196
rect 20996 17144 21048 17196
rect 21824 17144 21876 17196
rect 6000 17076 6052 17128
rect 9128 17076 9180 17128
rect 13268 17119 13320 17128
rect 4712 17051 4764 17060
rect 4712 17017 4721 17051
rect 4721 17017 4755 17051
rect 4755 17017 4764 17051
rect 4712 17008 4764 17017
rect 4804 17051 4856 17060
rect 4804 17017 4813 17051
rect 4813 17017 4847 17051
rect 4847 17017 4856 17051
rect 5356 17051 5408 17060
rect 4804 17008 4856 17017
rect 5356 17017 5365 17051
rect 5365 17017 5399 17051
rect 5399 17017 5408 17051
rect 5356 17008 5408 17017
rect 2320 16983 2372 16992
rect 2320 16949 2329 16983
rect 2329 16949 2363 16983
rect 2363 16949 2372 16983
rect 2320 16940 2372 16949
rect 2780 16983 2832 16992
rect 2780 16949 2789 16983
rect 2789 16949 2823 16983
rect 2823 16949 2832 16983
rect 2780 16940 2832 16949
rect 2964 16940 3016 16992
rect 4252 16940 4304 16992
rect 6368 16940 6420 16992
rect 7012 16940 7064 16992
rect 8576 17008 8628 17060
rect 9680 17008 9732 17060
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 10784 17008 10836 17060
rect 10876 17008 10928 17060
rect 13268 17085 13277 17119
rect 13277 17085 13311 17119
rect 13311 17085 13320 17119
rect 13268 17076 13320 17085
rect 15936 17076 15988 17128
rect 19432 17076 19484 17128
rect 20352 17076 20404 17128
rect 22560 17119 22612 17128
rect 22560 17085 22569 17119
rect 22569 17085 22603 17119
rect 22603 17085 22612 17119
rect 22560 17076 22612 17085
rect 23296 17076 23348 17128
rect 24584 17119 24636 17128
rect 24584 17085 24593 17119
rect 24593 17085 24627 17119
rect 24627 17085 24636 17119
rect 24584 17076 24636 17085
rect 13544 17008 13596 17060
rect 15476 17008 15528 17060
rect 16856 17008 16908 17060
rect 18144 17051 18196 17060
rect 18144 17017 18153 17051
rect 18153 17017 18187 17051
rect 18187 17017 18196 17051
rect 18144 17008 18196 17017
rect 18236 17051 18288 17060
rect 18236 17017 18245 17051
rect 18245 17017 18279 17051
rect 18279 17017 18288 17051
rect 18788 17051 18840 17060
rect 18236 17008 18288 17017
rect 18788 17017 18797 17051
rect 18797 17017 18831 17051
rect 18831 17017 18840 17051
rect 18788 17008 18840 17017
rect 21364 17008 21416 17060
rect 10968 16940 11020 16992
rect 11980 16983 12032 16992
rect 11980 16949 11989 16983
rect 11989 16949 12023 16983
rect 12023 16949 12032 16983
rect 11980 16940 12032 16949
rect 12808 16940 12860 16992
rect 14188 16983 14240 16992
rect 14188 16949 14197 16983
rect 14197 16949 14231 16983
rect 14231 16949 14240 16983
rect 14188 16940 14240 16949
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 18696 16940 18748 16992
rect 19524 16940 19576 16992
rect 23572 16940 23624 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 6828 16779 6880 16788
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 7932 16736 7984 16788
rect 8668 16779 8720 16788
rect 8668 16745 8677 16779
rect 8677 16745 8711 16779
rect 8711 16745 8720 16779
rect 8668 16736 8720 16745
rect 9496 16736 9548 16788
rect 10692 16779 10744 16788
rect 4252 16668 4304 16720
rect 4712 16668 4764 16720
rect 6000 16711 6052 16720
rect 6000 16677 6009 16711
rect 6009 16677 6043 16711
rect 6043 16677 6052 16711
rect 6000 16668 6052 16677
rect 7840 16711 7892 16720
rect 7840 16677 7849 16711
rect 7849 16677 7883 16711
rect 7883 16677 7892 16711
rect 7840 16668 7892 16677
rect 9220 16668 9272 16720
rect 10692 16745 10701 16779
rect 10701 16745 10735 16779
rect 10735 16745 10744 16779
rect 10692 16736 10744 16745
rect 14096 16736 14148 16788
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 18144 16736 18196 16788
rect 21088 16779 21140 16788
rect 11428 16711 11480 16720
rect 11428 16677 11437 16711
rect 11437 16677 11471 16711
rect 11471 16677 11480 16711
rect 11428 16668 11480 16677
rect 13728 16668 13780 16720
rect 14188 16668 14240 16720
rect 15292 16668 15344 16720
rect 15844 16668 15896 16720
rect 17500 16668 17552 16720
rect 19340 16711 19392 16720
rect 19340 16677 19349 16711
rect 19349 16677 19383 16711
rect 19383 16677 19392 16711
rect 19340 16668 19392 16677
rect 21088 16745 21097 16779
rect 21097 16745 21131 16779
rect 21131 16745 21140 16779
rect 21088 16736 21140 16745
rect 19984 16668 20036 16720
rect 2596 16600 2648 16652
rect 3148 16600 3200 16652
rect 4344 16600 4396 16652
rect 4620 16532 4672 16584
rect 21088 16600 21140 16652
rect 22100 16600 22152 16652
rect 22928 16643 22980 16652
rect 22928 16609 22937 16643
rect 22937 16609 22971 16643
rect 22971 16609 22980 16643
rect 22928 16600 22980 16609
rect 25228 16600 25280 16652
rect 6184 16532 6236 16584
rect 7748 16575 7800 16584
rect 7748 16541 7757 16575
rect 7757 16541 7791 16575
rect 7791 16541 7800 16575
rect 7748 16532 7800 16541
rect 8668 16532 8720 16584
rect 10876 16532 10928 16584
rect 11612 16532 11664 16584
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 13176 16575 13228 16584
rect 11704 16532 11756 16541
rect 13176 16541 13185 16575
rect 13185 16541 13219 16575
rect 13219 16541 13228 16575
rect 13176 16532 13228 16541
rect 15476 16532 15528 16584
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 5356 16464 5408 16516
rect 8116 16464 8168 16516
rect 8300 16507 8352 16516
rect 8300 16473 8309 16507
rect 8309 16473 8343 16507
rect 8343 16473 8352 16507
rect 8300 16464 8352 16473
rect 18788 16532 18840 16584
rect 19248 16575 19300 16584
rect 19248 16541 19257 16575
rect 19257 16541 19291 16575
rect 19291 16541 19300 16575
rect 19248 16532 19300 16541
rect 22652 16532 22704 16584
rect 24676 16464 24728 16516
rect 2136 16439 2188 16448
rect 2136 16405 2145 16439
rect 2145 16405 2179 16439
rect 2179 16405 2188 16439
rect 2136 16396 2188 16405
rect 7564 16396 7616 16448
rect 9036 16396 9088 16448
rect 10876 16396 10928 16448
rect 11244 16396 11296 16448
rect 11888 16396 11940 16448
rect 13268 16396 13320 16448
rect 14096 16439 14148 16448
rect 14096 16405 14105 16439
rect 14105 16405 14139 16439
rect 14139 16405 14148 16439
rect 14096 16396 14148 16405
rect 15292 16396 15344 16448
rect 20628 16396 20680 16448
rect 22284 16396 22336 16448
rect 24860 16396 24912 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 4804 16192 4856 16244
rect 6000 16192 6052 16244
rect 6184 16235 6236 16244
rect 6184 16201 6193 16235
rect 6193 16201 6227 16235
rect 6227 16201 6236 16235
rect 6184 16192 6236 16201
rect 6736 16192 6788 16244
rect 7840 16192 7892 16244
rect 9496 16192 9548 16244
rect 9680 16235 9732 16244
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 15844 16235 15896 16244
rect 15844 16201 15853 16235
rect 15853 16201 15887 16235
rect 15887 16201 15896 16235
rect 15844 16192 15896 16201
rect 17500 16235 17552 16244
rect 11428 16124 11480 16176
rect 15476 16167 15528 16176
rect 15476 16133 15485 16167
rect 15485 16133 15519 16167
rect 15519 16133 15528 16167
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 19248 16192 19300 16244
rect 21088 16235 21140 16244
rect 21088 16201 21097 16235
rect 21097 16201 21131 16235
rect 21131 16201 21140 16235
rect 21088 16192 21140 16201
rect 22008 16235 22060 16244
rect 22008 16201 22017 16235
rect 22017 16201 22051 16235
rect 22051 16201 22060 16235
rect 22008 16192 22060 16201
rect 24768 16235 24820 16244
rect 24768 16201 24777 16235
rect 24777 16201 24811 16235
rect 24811 16201 24820 16235
rect 24768 16192 24820 16201
rect 15476 16124 15528 16133
rect 5540 16056 5592 16108
rect 6736 16056 6788 16108
rect 7564 16056 7616 16108
rect 8668 16056 8720 16108
rect 9772 16056 9824 16108
rect 10784 16056 10836 16108
rect 15292 16056 15344 16108
rect 15384 16056 15436 16108
rect 16488 16099 16540 16108
rect 16488 16065 16497 16099
rect 16497 16065 16531 16099
rect 16531 16065 16540 16099
rect 16488 16056 16540 16065
rect 2044 16031 2096 16040
rect 2044 15997 2053 16031
rect 2053 15997 2087 16031
rect 2087 15997 2096 16031
rect 2044 15988 2096 15997
rect 2872 15988 2924 16040
rect 2228 15920 2280 15972
rect 3424 15988 3476 16040
rect 5264 15920 5316 15972
rect 13084 16031 13136 16040
rect 7840 15963 7892 15972
rect 7840 15929 7849 15963
rect 7849 15929 7883 15963
rect 7883 15929 7892 15963
rect 7840 15920 7892 15929
rect 8484 15920 8536 15972
rect 13084 15997 13093 16031
rect 13093 15997 13127 16031
rect 13127 15997 13136 16031
rect 13084 15988 13136 15997
rect 1216 15852 1268 15904
rect 3148 15852 3200 15904
rect 4252 15852 4304 15904
rect 5356 15895 5408 15904
rect 5356 15861 5365 15895
rect 5365 15861 5399 15895
rect 5399 15861 5408 15895
rect 5356 15852 5408 15861
rect 9680 15852 9732 15904
rect 12992 15920 13044 15972
rect 13268 15920 13320 15972
rect 13728 15920 13780 15972
rect 14096 15920 14148 15972
rect 14924 15920 14976 15972
rect 16580 15963 16632 15972
rect 16580 15929 16589 15963
rect 16589 15929 16623 15963
rect 16623 15929 16632 15963
rect 16580 15920 16632 15929
rect 20076 16124 20128 16176
rect 18604 16056 18656 16108
rect 19524 16056 19576 16108
rect 19984 16099 20036 16108
rect 19984 16065 19993 16099
rect 19993 16065 20027 16099
rect 20027 16065 20036 16099
rect 19984 16056 20036 16065
rect 20168 16056 20220 16108
rect 18788 15963 18840 15972
rect 11612 15895 11664 15904
rect 11612 15861 11621 15895
rect 11621 15861 11655 15895
rect 11655 15861 11664 15895
rect 11612 15852 11664 15861
rect 15568 15852 15620 15904
rect 16304 15852 16356 15904
rect 18788 15929 18797 15963
rect 18797 15929 18831 15963
rect 18831 15929 18840 15963
rect 18788 15920 18840 15929
rect 19248 15920 19300 15972
rect 19340 15852 19392 15904
rect 22008 15988 22060 16040
rect 22928 15988 22980 16040
rect 22192 15852 22244 15904
rect 22928 15895 22980 15904
rect 22928 15861 22937 15895
rect 22937 15861 22971 15895
rect 22971 15861 22980 15895
rect 22928 15852 22980 15861
rect 25228 15852 25280 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1124 15648 1176 15700
rect 2872 15648 2924 15700
rect 3148 15691 3200 15700
rect 3148 15657 3157 15691
rect 3157 15657 3191 15691
rect 3191 15657 3200 15691
rect 3148 15648 3200 15657
rect 3516 15648 3568 15700
rect 4620 15691 4672 15700
rect 4252 15623 4304 15632
rect 4252 15589 4261 15623
rect 4261 15589 4295 15623
rect 4295 15589 4304 15623
rect 4252 15580 4304 15589
rect 4620 15657 4629 15691
rect 4629 15657 4663 15691
rect 4663 15657 4672 15691
rect 4620 15648 4672 15657
rect 5080 15648 5132 15700
rect 5540 15648 5592 15700
rect 7840 15648 7892 15700
rect 9220 15648 9272 15700
rect 11520 15648 11572 15700
rect 13176 15648 13228 15700
rect 13268 15648 13320 15700
rect 14924 15691 14976 15700
rect 14924 15657 14933 15691
rect 14933 15657 14967 15691
rect 14967 15657 14976 15691
rect 14924 15648 14976 15657
rect 16488 15691 16540 15700
rect 16488 15657 16497 15691
rect 16497 15657 16531 15691
rect 16531 15657 16540 15691
rect 16488 15648 16540 15657
rect 18328 15648 18380 15700
rect 18604 15691 18656 15700
rect 18604 15657 18613 15691
rect 18613 15657 18647 15691
rect 18647 15657 18656 15691
rect 18604 15648 18656 15657
rect 19524 15648 19576 15700
rect 20812 15648 20864 15700
rect 22008 15648 22060 15700
rect 23848 15648 23900 15700
rect 6184 15580 6236 15632
rect 7012 15580 7064 15632
rect 7564 15580 7616 15632
rect 11612 15580 11664 15632
rect 13084 15580 13136 15632
rect 14740 15580 14792 15632
rect 17316 15623 17368 15632
rect 17316 15589 17325 15623
rect 17325 15589 17359 15623
rect 17359 15589 17368 15623
rect 17316 15580 17368 15589
rect 17684 15580 17736 15632
rect 18788 15580 18840 15632
rect 18972 15580 19024 15632
rect 19984 15580 20036 15632
rect 21272 15623 21324 15632
rect 21272 15589 21281 15623
rect 21281 15589 21315 15623
rect 21315 15589 21324 15623
rect 21272 15580 21324 15589
rect 21456 15580 21508 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 3424 15512 3476 15564
rect 5080 15555 5132 15564
rect 5080 15521 5089 15555
rect 5089 15521 5123 15555
rect 5123 15521 5132 15555
rect 5080 15512 5132 15521
rect 5540 15555 5592 15564
rect 5540 15521 5549 15555
rect 5549 15521 5583 15555
rect 5583 15521 5592 15555
rect 5540 15512 5592 15521
rect 8484 15512 8536 15564
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 2596 15444 2648 15496
rect 5264 15444 5316 15496
rect 8024 15444 8076 15496
rect 10140 15512 10192 15564
rect 10876 15512 10928 15564
rect 11428 15555 11480 15564
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 11888 15555 11940 15564
rect 11888 15521 11897 15555
rect 11897 15521 11931 15555
rect 11931 15521 11940 15555
rect 11888 15512 11940 15521
rect 22928 15512 22980 15564
rect 24216 15512 24268 15564
rect 25136 15512 25188 15564
rect 12348 15444 12400 15496
rect 2228 15308 2280 15360
rect 9864 15376 9916 15428
rect 4068 15308 4120 15360
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 7840 15351 7892 15360
rect 7840 15317 7849 15351
rect 7849 15317 7883 15351
rect 7883 15317 7892 15351
rect 7840 15308 7892 15317
rect 12624 15308 12676 15360
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 15476 15444 15528 15496
rect 14740 15308 14792 15360
rect 18604 15444 18656 15496
rect 21180 15487 21232 15496
rect 21180 15453 21189 15487
rect 21189 15453 21223 15487
rect 21223 15453 21232 15487
rect 21180 15444 21232 15453
rect 22100 15487 22152 15496
rect 17224 15308 17276 15360
rect 20168 15376 20220 15428
rect 21088 15376 21140 15428
rect 22100 15453 22109 15487
rect 22109 15453 22143 15487
rect 22143 15453 22152 15487
rect 22100 15444 22152 15453
rect 21640 15376 21692 15428
rect 17500 15308 17552 15360
rect 21916 15308 21968 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2136 15147 2188 15156
rect 2136 15113 2145 15147
rect 2145 15113 2179 15147
rect 2179 15113 2188 15147
rect 2136 15104 2188 15113
rect 3056 15147 3108 15156
rect 3056 15113 3065 15147
rect 3065 15113 3099 15147
rect 3099 15113 3108 15147
rect 3056 15104 3108 15113
rect 3424 15147 3476 15156
rect 3424 15113 3433 15147
rect 3433 15113 3467 15147
rect 3467 15113 3476 15147
rect 3424 15104 3476 15113
rect 4896 15104 4948 15156
rect 7104 15104 7156 15156
rect 8024 15147 8076 15156
rect 1400 15036 1452 15088
rect 7564 15036 7616 15088
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 9864 15147 9916 15156
rect 9864 15113 9873 15147
rect 9873 15113 9907 15147
rect 9907 15113 9916 15147
rect 9864 15104 9916 15113
rect 9680 15036 9732 15088
rect 10140 15036 10192 15088
rect 2136 14900 2188 14952
rect 3056 14900 3108 14952
rect 3148 14900 3200 14952
rect 3516 14900 3568 14952
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 4620 14968 4672 15020
rect 4896 14968 4948 15020
rect 5172 14943 5224 14952
rect 5172 14909 5181 14943
rect 5181 14909 5215 14943
rect 5215 14909 5224 14943
rect 5172 14900 5224 14909
rect 6368 14968 6420 15020
rect 8668 14968 8720 15020
rect 8024 14900 8076 14952
rect 10968 15104 11020 15156
rect 11244 15104 11296 15156
rect 12992 15104 13044 15156
rect 14740 15147 14792 15156
rect 14740 15113 14749 15147
rect 14749 15113 14783 15147
rect 14783 15113 14792 15147
rect 14740 15104 14792 15113
rect 17316 15104 17368 15156
rect 18972 15104 19024 15156
rect 21272 15104 21324 15156
rect 22928 15104 22980 15156
rect 23112 15147 23164 15156
rect 23112 15113 23121 15147
rect 23121 15113 23155 15147
rect 23155 15113 23164 15147
rect 23112 15104 23164 15113
rect 25136 15147 25188 15156
rect 25136 15113 25145 15147
rect 25145 15113 25179 15147
rect 25179 15113 25188 15147
rect 25136 15104 25188 15113
rect 11428 15036 11480 15088
rect 17132 15036 17184 15088
rect 18604 15036 18656 15088
rect 21180 15036 21232 15088
rect 10692 14968 10744 15020
rect 11520 15011 11572 15020
rect 11520 14977 11529 15011
rect 11529 14977 11563 15011
rect 11563 14977 11572 15011
rect 11520 14968 11572 14977
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 15844 15011 15896 15020
rect 15844 14977 15853 15011
rect 15853 14977 15887 15011
rect 15887 14977 15896 15011
rect 15844 14968 15896 14977
rect 16580 14968 16632 15020
rect 11888 14900 11940 14952
rect 12900 14900 12952 14952
rect 2780 14832 2832 14884
rect 3424 14832 3476 14884
rect 6828 14832 6880 14884
rect 8668 14875 8720 14884
rect 8668 14841 8677 14875
rect 8677 14841 8711 14875
rect 8711 14841 8720 14875
rect 8668 14832 8720 14841
rect 8760 14875 8812 14884
rect 8760 14841 8769 14875
rect 8769 14841 8803 14875
rect 8803 14841 8812 14875
rect 8760 14832 8812 14841
rect 3884 14764 3936 14816
rect 4160 14764 4212 14816
rect 5080 14807 5132 14816
rect 5080 14773 5089 14807
rect 5089 14773 5123 14807
rect 5123 14773 5132 14807
rect 5080 14764 5132 14773
rect 5264 14764 5316 14816
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 8576 14764 8628 14816
rect 16488 14900 16540 14952
rect 14188 14832 14240 14884
rect 13176 14764 13228 14816
rect 15292 14764 15344 14816
rect 15476 14875 15528 14884
rect 15476 14841 15485 14875
rect 15485 14841 15519 14875
rect 15519 14841 15528 14875
rect 15476 14832 15528 14841
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 17316 14764 17368 14816
rect 18328 14968 18380 15020
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 20168 14968 20220 15020
rect 22468 14968 22520 15020
rect 19432 14900 19484 14952
rect 20536 14943 20588 14952
rect 19248 14832 19300 14884
rect 20536 14909 20545 14943
rect 20545 14909 20579 14943
rect 20579 14909 20588 14943
rect 20536 14900 20588 14909
rect 20720 14900 20772 14952
rect 23112 14900 23164 14952
rect 21180 14832 21232 14884
rect 24032 14832 24084 14884
rect 18512 14764 18564 14816
rect 20996 14764 21048 14816
rect 23204 14764 23256 14816
rect 24216 14764 24268 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 2688 14560 2740 14612
rect 3424 14560 3476 14612
rect 3516 14560 3568 14612
rect 4160 14603 4212 14612
rect 4160 14569 4169 14603
rect 4169 14569 4203 14603
rect 4203 14569 4212 14603
rect 4160 14560 4212 14569
rect 8668 14560 8720 14612
rect 10692 14560 10744 14612
rect 13820 14603 13872 14612
rect 7748 14535 7800 14544
rect 7748 14501 7757 14535
rect 7757 14501 7791 14535
rect 7791 14501 7800 14535
rect 7748 14492 7800 14501
rect 8116 14492 8168 14544
rect 8760 14492 8812 14544
rect 13820 14569 13829 14603
rect 13829 14569 13863 14603
rect 13863 14569 13872 14603
rect 13820 14560 13872 14569
rect 14188 14603 14240 14612
rect 14188 14569 14197 14603
rect 14197 14569 14231 14603
rect 14231 14569 14240 14603
rect 14188 14560 14240 14569
rect 14832 14560 14884 14612
rect 15384 14560 15436 14612
rect 17224 14603 17276 14612
rect 17224 14569 17233 14603
rect 17233 14569 17267 14603
rect 17267 14569 17276 14603
rect 17224 14560 17276 14569
rect 19432 14603 19484 14612
rect 19432 14569 19441 14603
rect 19441 14569 19475 14603
rect 19475 14569 19484 14603
rect 19432 14560 19484 14569
rect 20536 14560 20588 14612
rect 24768 14603 24820 14612
rect 24768 14569 24777 14603
rect 24777 14569 24811 14603
rect 24811 14569 24820 14603
rect 24768 14560 24820 14569
rect 12624 14492 12676 14544
rect 12992 14535 13044 14544
rect 12992 14501 13001 14535
rect 13001 14501 13035 14535
rect 13035 14501 13044 14535
rect 12992 14492 13044 14501
rect 14096 14492 14148 14544
rect 17592 14535 17644 14544
rect 17592 14501 17601 14535
rect 17601 14501 17635 14535
rect 17635 14501 17644 14535
rect 17592 14492 17644 14501
rect 18236 14492 18288 14544
rect 21088 14535 21140 14544
rect 21088 14501 21097 14535
rect 21097 14501 21131 14535
rect 21131 14501 21140 14535
rect 21088 14492 21140 14501
rect 1584 14424 1636 14476
rect 2688 14424 2740 14476
rect 4068 14467 4120 14476
rect 4068 14433 4077 14467
rect 4077 14433 4111 14467
rect 4111 14433 4120 14467
rect 4068 14424 4120 14433
rect 4528 14467 4580 14476
rect 4528 14433 4537 14467
rect 4537 14433 4571 14467
rect 4571 14433 4580 14467
rect 4528 14424 4580 14433
rect 5172 14467 5224 14476
rect 5172 14433 5181 14467
rect 5181 14433 5215 14467
rect 5215 14433 5224 14467
rect 5172 14424 5224 14433
rect 5540 14467 5592 14476
rect 5540 14433 5549 14467
rect 5549 14433 5583 14467
rect 5583 14433 5592 14467
rect 5540 14424 5592 14433
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 9864 14467 9916 14476
rect 9864 14433 9873 14467
rect 9873 14433 9907 14467
rect 9907 14433 9916 14467
rect 9864 14424 9916 14433
rect 10048 14424 10100 14476
rect 11244 14467 11296 14476
rect 11244 14433 11253 14467
rect 11253 14433 11287 14467
rect 11287 14433 11296 14467
rect 11244 14424 11296 14433
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 20536 14424 20588 14476
rect 20720 14424 20772 14476
rect 22468 14467 22520 14476
rect 22468 14433 22477 14467
rect 22477 14433 22511 14467
rect 22511 14433 22520 14467
rect 22468 14424 22520 14433
rect 23020 14467 23072 14476
rect 23020 14433 23029 14467
rect 23029 14433 23063 14467
rect 23063 14433 23072 14467
rect 23020 14424 23072 14433
rect 24860 14424 24912 14476
rect 6368 14399 6420 14408
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 7932 14356 7984 14408
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 9404 14356 9456 14408
rect 12164 14356 12216 14408
rect 14004 14356 14056 14408
rect 2320 14288 2372 14340
rect 5172 14220 5224 14272
rect 5540 14220 5592 14272
rect 7288 14220 7340 14272
rect 8208 14288 8260 14340
rect 10968 14288 11020 14340
rect 15568 14356 15620 14408
rect 19156 14356 19208 14408
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 15476 14288 15528 14340
rect 17500 14288 17552 14340
rect 19248 14288 19300 14340
rect 8944 14220 8996 14272
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 16672 14220 16724 14272
rect 20352 14288 20404 14340
rect 21548 14288 21600 14340
rect 22928 14288 22980 14340
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 21824 14220 21876 14272
rect 23664 14263 23716 14272
rect 23664 14229 23673 14263
rect 23673 14229 23707 14263
rect 23707 14229 23716 14263
rect 23664 14220 23716 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1768 14059 1820 14068
rect 1768 14025 1777 14059
rect 1777 14025 1811 14059
rect 1811 14025 1820 14059
rect 1768 14016 1820 14025
rect 3424 14016 3476 14068
rect 4068 14016 4120 14068
rect 6276 14016 6328 14068
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 9864 14016 9916 14068
rect 9956 14016 10008 14068
rect 5540 13948 5592 14000
rect 6552 13948 6604 14000
rect 6828 13948 6880 14000
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 5356 13923 5408 13932
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 4896 13812 4948 13821
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 5448 13880 5500 13932
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 7840 13948 7892 14000
rect 9036 13948 9088 14000
rect 10140 13948 10192 14000
rect 11704 13991 11756 14000
rect 11704 13957 11713 13991
rect 11713 13957 11747 13991
rect 11747 13957 11756 13991
rect 11704 13948 11756 13957
rect 12992 14016 13044 14068
rect 14004 14059 14056 14068
rect 14004 14025 14013 14059
rect 14013 14025 14047 14059
rect 14047 14025 14056 14059
rect 14004 14016 14056 14025
rect 14188 14016 14240 14068
rect 18236 14016 18288 14068
rect 19984 14016 20036 14068
rect 21088 14016 21140 14068
rect 22468 14059 22520 14068
rect 22468 14025 22477 14059
rect 22477 14025 22511 14059
rect 22511 14025 22520 14059
rect 22468 14016 22520 14025
rect 24860 14016 24912 14068
rect 15384 13948 15436 14000
rect 15844 13948 15896 14000
rect 17224 13948 17276 14000
rect 19248 13948 19300 14000
rect 5264 13812 5316 13864
rect 11888 13880 11940 13932
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 15200 13880 15252 13932
rect 20076 13880 20128 13932
rect 21548 13880 21600 13932
rect 21640 13880 21692 13932
rect 22376 13880 22428 13932
rect 24768 13880 24820 13932
rect 9220 13812 9272 13864
rect 11428 13812 11480 13864
rect 11704 13812 11756 13864
rect 16304 13812 16356 13864
rect 4344 13744 4396 13796
rect 6092 13787 6144 13796
rect 6092 13753 6101 13787
rect 6101 13753 6135 13787
rect 6135 13753 6144 13787
rect 6092 13744 6144 13753
rect 2044 13719 2096 13728
rect 2044 13685 2053 13719
rect 2053 13685 2087 13719
rect 2087 13685 2096 13719
rect 2044 13676 2096 13685
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 3792 13676 3844 13685
rect 7288 13787 7340 13796
rect 7288 13753 7297 13787
rect 7297 13753 7331 13787
rect 7331 13753 7340 13787
rect 7288 13744 7340 13753
rect 9864 13744 9916 13796
rect 10140 13787 10192 13796
rect 10140 13753 10149 13787
rect 10149 13753 10183 13787
rect 10183 13753 10192 13787
rect 10692 13787 10744 13796
rect 10140 13744 10192 13753
rect 10692 13753 10701 13787
rect 10701 13753 10735 13787
rect 10735 13753 10744 13787
rect 10692 13744 10744 13753
rect 11244 13787 11296 13796
rect 11244 13753 11253 13787
rect 11253 13753 11287 13787
rect 11287 13753 11296 13787
rect 11244 13744 11296 13753
rect 15200 13787 15252 13796
rect 7748 13676 7800 13728
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 9496 13676 9548 13728
rect 9956 13676 10008 13728
rect 12164 13719 12216 13728
rect 12164 13685 12173 13719
rect 12173 13685 12207 13719
rect 12207 13685 12216 13719
rect 15200 13753 15209 13787
rect 15209 13753 15243 13787
rect 15243 13753 15252 13787
rect 15200 13744 15252 13753
rect 15292 13787 15344 13796
rect 15292 13753 15301 13787
rect 15301 13753 15335 13787
rect 15335 13753 15344 13787
rect 15292 13744 15344 13753
rect 18144 13787 18196 13796
rect 18144 13753 18153 13787
rect 18153 13753 18187 13787
rect 18187 13753 18196 13787
rect 18144 13744 18196 13753
rect 18236 13787 18288 13796
rect 18236 13753 18245 13787
rect 18245 13753 18279 13787
rect 18279 13753 18288 13787
rect 18236 13744 18288 13753
rect 18972 13744 19024 13796
rect 22744 13812 22796 13864
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 19524 13744 19576 13796
rect 19984 13787 20036 13796
rect 19984 13753 19993 13787
rect 19993 13753 20027 13787
rect 20027 13753 20036 13787
rect 19984 13744 20036 13753
rect 21824 13744 21876 13796
rect 24676 13812 24728 13864
rect 24860 13812 24912 13864
rect 25688 13855 25740 13864
rect 25688 13821 25697 13855
rect 25697 13821 25731 13855
rect 25731 13821 25740 13855
rect 25688 13812 25740 13821
rect 12164 13676 12216 13685
rect 12992 13676 13044 13728
rect 19064 13676 19116 13728
rect 20352 13676 20404 13728
rect 23020 13676 23072 13728
rect 23480 13719 23532 13728
rect 23480 13685 23489 13719
rect 23489 13685 23523 13719
rect 23523 13685 23532 13719
rect 23480 13676 23532 13685
rect 23756 13719 23808 13728
rect 23756 13685 23765 13719
rect 23765 13685 23799 13719
rect 23799 13685 23808 13719
rect 23756 13676 23808 13685
rect 24124 13676 24176 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2044 13472 2096 13524
rect 2688 13404 2740 13456
rect 3792 13404 3844 13456
rect 3976 13472 4028 13524
rect 4160 13472 4212 13524
rect 4344 13472 4396 13524
rect 4804 13472 4856 13524
rect 1676 13268 1728 13320
rect 2504 13268 2556 13320
rect 4528 13336 4580 13388
rect 6368 13472 6420 13524
rect 6552 13472 6604 13524
rect 7288 13472 7340 13524
rect 7472 13472 7524 13524
rect 8208 13447 8260 13456
rect 8208 13413 8217 13447
rect 8217 13413 8251 13447
rect 8251 13413 8260 13447
rect 8208 13404 8260 13413
rect 3240 13268 3292 13320
rect 3792 13268 3844 13320
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 4068 13268 4120 13277
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 9864 13472 9916 13524
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 12992 13515 13044 13524
rect 12992 13481 13001 13515
rect 13001 13481 13035 13515
rect 13035 13481 13044 13515
rect 12992 13472 13044 13481
rect 14188 13472 14240 13524
rect 17592 13472 17644 13524
rect 18144 13472 18196 13524
rect 19064 13472 19116 13524
rect 9588 13404 9640 13456
rect 15384 13404 15436 13456
rect 17040 13447 17092 13456
rect 17040 13413 17049 13447
rect 17049 13413 17083 13447
rect 17083 13413 17092 13447
rect 17040 13404 17092 13413
rect 18512 13404 18564 13456
rect 19248 13404 19300 13456
rect 20076 13472 20128 13524
rect 20996 13472 21048 13524
rect 23756 13472 23808 13524
rect 21548 13447 21600 13456
rect 21548 13413 21557 13447
rect 21557 13413 21591 13447
rect 21591 13413 21600 13447
rect 21548 13404 21600 13413
rect 22836 13404 22888 13456
rect 9404 13336 9456 13388
rect 9864 13336 9916 13388
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 9956 13268 10008 13320
rect 10140 13268 10192 13320
rect 12072 13336 12124 13388
rect 24768 13336 24820 13388
rect 12440 13268 12492 13320
rect 14556 13268 14608 13320
rect 16948 13311 17000 13320
rect 16948 13277 16957 13311
rect 16957 13277 16991 13311
rect 16991 13277 17000 13311
rect 16948 13268 17000 13277
rect 17224 13311 17276 13320
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 18972 13268 19024 13320
rect 21456 13311 21508 13320
rect 21456 13277 21465 13311
rect 21465 13277 21499 13311
rect 21499 13277 21508 13311
rect 21456 13268 21508 13277
rect 21640 13268 21692 13320
rect 23020 13311 23072 13320
rect 23020 13277 23029 13311
rect 23029 13277 23063 13311
rect 23063 13277 23072 13311
rect 23020 13268 23072 13277
rect 8576 13200 8628 13252
rect 10048 13200 10100 13252
rect 15476 13200 15528 13252
rect 15568 13200 15620 13252
rect 16028 13200 16080 13252
rect 22100 13200 22152 13252
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 2780 13132 2832 13184
rect 3976 13132 4028 13184
rect 4344 13132 4396 13184
rect 7748 13132 7800 13184
rect 7932 13175 7984 13184
rect 7932 13141 7941 13175
rect 7941 13141 7975 13175
rect 7975 13141 7984 13175
rect 7932 13132 7984 13141
rect 8300 13132 8352 13184
rect 8760 13132 8812 13184
rect 12808 13132 12860 13184
rect 13636 13132 13688 13184
rect 20996 13132 21048 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1676 12971 1728 12980
rect 1676 12937 1685 12971
rect 1685 12937 1719 12971
rect 1719 12937 1728 12971
rect 1676 12928 1728 12937
rect 2320 12928 2372 12980
rect 2688 12971 2740 12980
rect 2688 12937 2697 12971
rect 2697 12937 2731 12971
rect 2731 12937 2740 12971
rect 2688 12928 2740 12937
rect 3700 12971 3752 12980
rect 3700 12937 3709 12971
rect 3709 12937 3743 12971
rect 3743 12937 3752 12971
rect 3700 12928 3752 12937
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 6092 12928 6144 12980
rect 2412 12792 2464 12844
rect 3056 12792 3108 12844
rect 3792 12860 3844 12912
rect 7472 12860 7524 12912
rect 8208 12928 8260 12980
rect 8300 12928 8352 12980
rect 12992 12928 13044 12980
rect 13728 12928 13780 12980
rect 15384 12971 15436 12980
rect 15384 12937 15393 12971
rect 15393 12937 15427 12971
rect 15427 12937 15436 12971
rect 15384 12928 15436 12937
rect 21548 12928 21600 12980
rect 23020 12928 23072 12980
rect 24952 12971 25004 12980
rect 24952 12937 24961 12971
rect 24961 12937 24995 12971
rect 24995 12937 25004 12971
rect 24952 12928 25004 12937
rect 8760 12903 8812 12912
rect 8760 12869 8769 12903
rect 8769 12869 8803 12903
rect 8803 12869 8812 12903
rect 8760 12860 8812 12869
rect 10968 12860 11020 12912
rect 4068 12792 4120 12844
rect 6552 12792 6604 12844
rect 9128 12792 9180 12844
rect 3700 12724 3752 12776
rect 6828 12767 6880 12776
rect 4344 12656 4396 12708
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 6920 12724 6972 12776
rect 14832 12860 14884 12912
rect 12992 12792 13044 12844
rect 13636 12835 13688 12844
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 16396 12860 16448 12912
rect 25596 12903 25648 12912
rect 25596 12869 25605 12903
rect 25605 12869 25639 12903
rect 25639 12869 25648 12903
rect 25596 12860 25648 12869
rect 16028 12792 16080 12844
rect 17316 12792 17368 12844
rect 18788 12792 18840 12844
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 21180 12792 21232 12844
rect 6000 12656 6052 12708
rect 6552 12656 6604 12708
rect 9956 12699 10008 12708
rect 9956 12665 9965 12699
rect 9965 12665 9999 12699
rect 9999 12665 10008 12699
rect 9956 12656 10008 12665
rect 10968 12656 11020 12708
rect 3332 12631 3384 12640
rect 3332 12597 3341 12631
rect 3341 12597 3375 12631
rect 3375 12597 3384 12631
rect 3332 12588 3384 12597
rect 5908 12631 5960 12640
rect 5908 12597 5917 12631
rect 5917 12597 5951 12631
rect 5951 12597 5960 12631
rect 5908 12588 5960 12597
rect 8116 12588 8168 12640
rect 8484 12631 8536 12640
rect 8484 12597 8493 12631
rect 8493 12597 8527 12631
rect 8527 12597 8536 12631
rect 8484 12588 8536 12597
rect 9404 12588 9456 12640
rect 9588 12631 9640 12640
rect 9588 12597 9597 12631
rect 9597 12597 9631 12631
rect 9631 12597 9640 12631
rect 9588 12588 9640 12597
rect 9680 12588 9732 12640
rect 13728 12699 13780 12708
rect 13728 12665 13737 12699
rect 13737 12665 13771 12699
rect 13771 12665 13780 12699
rect 13728 12656 13780 12665
rect 11980 12588 12032 12640
rect 12072 12588 12124 12640
rect 12900 12588 12952 12640
rect 13912 12588 13964 12640
rect 14556 12631 14608 12640
rect 14556 12597 14565 12631
rect 14565 12597 14599 12631
rect 14599 12597 14608 12631
rect 14556 12588 14608 12597
rect 16948 12656 17000 12708
rect 18420 12699 18472 12708
rect 18420 12665 18429 12699
rect 18429 12665 18463 12699
rect 18463 12665 18472 12699
rect 18420 12656 18472 12665
rect 18696 12656 18748 12708
rect 19984 12724 20036 12776
rect 20996 12724 21048 12776
rect 21456 12724 21508 12776
rect 22284 12724 22336 12776
rect 24952 12724 25004 12776
rect 17040 12588 17092 12640
rect 17224 12631 17276 12640
rect 17224 12597 17233 12631
rect 17233 12597 17267 12631
rect 17267 12597 17276 12631
rect 17224 12588 17276 12597
rect 19340 12588 19392 12640
rect 22836 12656 22888 12708
rect 21272 12588 21324 12640
rect 22284 12588 22336 12640
rect 22560 12588 22612 12640
rect 23664 12588 23716 12640
rect 24768 12588 24820 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1952 12384 2004 12436
rect 3976 12384 4028 12436
rect 4068 12384 4120 12436
rect 6552 12384 6604 12436
rect 9864 12427 9916 12436
rect 9864 12393 9873 12427
rect 9873 12393 9907 12427
rect 9907 12393 9916 12427
rect 9864 12384 9916 12393
rect 9956 12384 10008 12436
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 16396 12427 16448 12436
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 18236 12384 18288 12436
rect 18512 12427 18564 12436
rect 18512 12393 18521 12427
rect 18521 12393 18555 12427
rect 18555 12393 18564 12427
rect 18512 12384 18564 12393
rect 19340 12384 19392 12436
rect 20812 12384 20864 12436
rect 21088 12384 21140 12436
rect 21272 12427 21324 12436
rect 21272 12393 21281 12427
rect 21281 12393 21315 12427
rect 21315 12393 21324 12427
rect 21272 12384 21324 12393
rect 21824 12427 21876 12436
rect 21824 12393 21833 12427
rect 21833 12393 21867 12427
rect 21867 12393 21876 12427
rect 21824 12384 21876 12393
rect 22100 12427 22152 12436
rect 22100 12393 22109 12427
rect 22109 12393 22143 12427
rect 22143 12393 22152 12427
rect 22100 12384 22152 12393
rect 22284 12384 22336 12436
rect 1492 12248 1544 12300
rect 2320 12248 2372 12300
rect 2872 12291 2924 12300
rect 2872 12257 2881 12291
rect 2881 12257 2915 12291
rect 2915 12257 2924 12291
rect 2872 12248 2924 12257
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 4252 12316 4304 12368
rect 4528 12316 4580 12368
rect 4436 12248 4488 12300
rect 6828 12316 6880 12368
rect 9680 12316 9732 12368
rect 10876 12316 10928 12368
rect 12164 12316 12216 12368
rect 15384 12316 15436 12368
rect 16120 12316 16172 12368
rect 16948 12316 17000 12368
rect 18788 12359 18840 12368
rect 18788 12325 18797 12359
rect 18797 12325 18831 12359
rect 18831 12325 18840 12359
rect 18788 12316 18840 12325
rect 19432 12359 19484 12368
rect 19432 12325 19441 12359
rect 19441 12325 19475 12359
rect 19475 12325 19484 12359
rect 19432 12316 19484 12325
rect 20536 12316 20588 12368
rect 20996 12316 21048 12368
rect 22560 12316 22612 12368
rect 23204 12384 23256 12436
rect 23848 12384 23900 12436
rect 5448 12248 5500 12300
rect 6092 12291 6144 12300
rect 6092 12257 6101 12291
rect 6101 12257 6135 12291
rect 6135 12257 6144 12291
rect 6092 12248 6144 12257
rect 8024 12248 8076 12300
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 8576 12291 8628 12300
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 21640 12248 21692 12300
rect 24584 12248 24636 12300
rect 25412 12248 25464 12300
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 4344 12180 4396 12232
rect 5908 12180 5960 12232
rect 6828 12180 6880 12232
rect 10784 12180 10836 12232
rect 10968 12223 11020 12232
rect 10968 12189 10977 12223
rect 10977 12189 11011 12223
rect 11011 12189 11020 12223
rect 10968 12180 11020 12189
rect 13084 12180 13136 12232
rect 14096 12180 14148 12232
rect 14832 12180 14884 12232
rect 17776 12180 17828 12232
rect 20076 12180 20128 12232
rect 20904 12223 20956 12232
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 22928 12180 22980 12232
rect 4160 12112 4212 12164
rect 4528 12112 4580 12164
rect 4896 12112 4948 12164
rect 6736 12112 6788 12164
rect 13728 12112 13780 12164
rect 22376 12112 22428 12164
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 2044 12044 2096 12096
rect 4620 12044 4672 12096
rect 8024 12044 8076 12096
rect 12900 12044 12952 12096
rect 13176 12044 13228 12096
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 20720 12087 20772 12096
rect 20720 12053 20729 12087
rect 20729 12053 20763 12087
rect 20763 12053 20772 12087
rect 20720 12044 20772 12053
rect 23572 12044 23624 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2320 11840 2372 11892
rect 3424 11840 3476 11892
rect 5448 11840 5500 11892
rect 7104 11840 7156 11892
rect 8300 11840 8352 11892
rect 10784 11840 10836 11892
rect 7748 11772 7800 11824
rect 10692 11772 10744 11824
rect 2412 11636 2464 11688
rect 3424 11636 3476 11688
rect 4344 11679 4396 11688
rect 4344 11645 4353 11679
rect 4353 11645 4387 11679
rect 4387 11645 4396 11679
rect 4344 11636 4396 11645
rect 4620 11679 4672 11688
rect 1492 11500 1544 11552
rect 4068 11568 4120 11620
rect 2596 11500 2648 11552
rect 3424 11500 3476 11552
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 5540 11636 5592 11688
rect 9864 11704 9916 11756
rect 12348 11772 12400 11824
rect 17316 11840 17368 11892
rect 21548 11840 21600 11892
rect 22284 11883 22336 11892
rect 22284 11849 22293 11883
rect 22293 11849 22327 11883
rect 22327 11849 22336 11883
rect 22284 11840 22336 11849
rect 24676 11883 24728 11892
rect 11612 11704 11664 11756
rect 11888 11704 11940 11756
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 14188 11704 14240 11756
rect 15752 11704 15804 11756
rect 19432 11772 19484 11824
rect 20076 11772 20128 11824
rect 16120 11704 16172 11756
rect 20720 11747 20772 11756
rect 20720 11713 20729 11747
rect 20729 11713 20763 11747
rect 20763 11713 20772 11747
rect 20720 11704 20772 11713
rect 22100 11704 22152 11756
rect 22928 11747 22980 11756
rect 22928 11713 22937 11747
rect 22937 11713 22971 11747
rect 22971 11713 22980 11747
rect 22928 11704 22980 11713
rect 14740 11636 14792 11688
rect 6092 11611 6144 11620
rect 6092 11577 6101 11611
rect 6101 11577 6135 11611
rect 6135 11577 6144 11611
rect 6092 11568 6144 11577
rect 4528 11500 4580 11552
rect 7748 11568 7800 11620
rect 8024 11611 8076 11620
rect 8024 11577 8033 11611
rect 8033 11577 8067 11611
rect 8067 11577 8076 11611
rect 8024 11568 8076 11577
rect 12164 11611 12216 11620
rect 12164 11577 12173 11611
rect 12173 11577 12207 11611
rect 12207 11577 12216 11611
rect 12164 11568 12216 11577
rect 13268 11611 13320 11620
rect 13268 11577 13277 11611
rect 13277 11577 13311 11611
rect 13311 11577 13320 11611
rect 13268 11568 13320 11577
rect 8576 11500 8628 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10876 11543 10928 11552
rect 10876 11509 10885 11543
rect 10885 11509 10919 11543
rect 10919 11509 10928 11543
rect 10876 11500 10928 11509
rect 13912 11500 13964 11552
rect 14188 11500 14240 11552
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 18972 11636 19024 11688
rect 20904 11636 20956 11688
rect 23020 11636 23072 11688
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 23940 11772 23992 11824
rect 23572 11636 23624 11688
rect 16948 11500 17000 11552
rect 19524 11568 19576 11620
rect 21272 11568 21324 11620
rect 23112 11568 23164 11620
rect 23480 11611 23532 11620
rect 23480 11577 23489 11611
rect 23489 11577 23523 11611
rect 23523 11577 23532 11611
rect 25504 11636 25556 11688
rect 23480 11568 23532 11577
rect 17776 11500 17828 11552
rect 21180 11500 21232 11552
rect 21824 11500 21876 11552
rect 23756 11543 23808 11552
rect 23756 11509 23765 11543
rect 23765 11509 23799 11543
rect 23799 11509 23808 11543
rect 23756 11500 23808 11509
rect 25412 11500 25464 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2412 11296 2464 11348
rect 3332 11296 3384 11348
rect 6552 11296 6604 11348
rect 7656 11296 7708 11348
rect 8024 11296 8076 11348
rect 12808 11339 12860 11348
rect 12808 11305 12817 11339
rect 12817 11305 12851 11339
rect 12851 11305 12860 11339
rect 12808 11296 12860 11305
rect 13084 11339 13136 11348
rect 13084 11305 13093 11339
rect 13093 11305 13127 11339
rect 13127 11305 13136 11339
rect 13084 11296 13136 11305
rect 2044 11228 2096 11280
rect 4344 11228 4396 11280
rect 4804 11228 4856 11280
rect 7748 11228 7800 11280
rect 10876 11271 10928 11280
rect 10876 11237 10885 11271
rect 10885 11237 10919 11271
rect 10919 11237 10928 11271
rect 10876 11228 10928 11237
rect 15292 11296 15344 11348
rect 18420 11296 18472 11348
rect 20076 11296 20128 11348
rect 20352 11296 20404 11348
rect 20904 11296 20956 11348
rect 22560 11296 22612 11348
rect 24952 11339 25004 11348
rect 24952 11305 24961 11339
rect 24961 11305 24995 11339
rect 24995 11305 25004 11339
rect 24952 11296 25004 11305
rect 14188 11228 14240 11280
rect 14832 11228 14884 11280
rect 15660 11271 15712 11280
rect 15660 11237 15669 11271
rect 15669 11237 15703 11271
rect 15703 11237 15712 11271
rect 15660 11228 15712 11237
rect 16948 11228 17000 11280
rect 19984 11271 20036 11280
rect 19984 11237 19993 11271
rect 19993 11237 20027 11271
rect 20027 11237 20036 11271
rect 19984 11228 20036 11237
rect 23480 11271 23532 11280
rect 23480 11237 23489 11271
rect 23489 11237 23523 11271
rect 23523 11237 23532 11271
rect 23480 11228 23532 11237
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 2688 11203 2740 11212
rect 2688 11169 2697 11203
rect 2697 11169 2731 11203
rect 2731 11169 2740 11203
rect 2688 11160 2740 11169
rect 4252 11203 4304 11212
rect 4252 11169 4261 11203
rect 4261 11169 4295 11203
rect 4295 11169 4304 11203
rect 4252 11160 4304 11169
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 4620 11160 4672 11212
rect 5172 11160 5224 11212
rect 6368 11160 6420 11212
rect 1676 11092 1728 11144
rect 5448 11092 5500 11144
rect 8392 11160 8444 11212
rect 8668 11160 8720 11212
rect 10508 11160 10560 11212
rect 12164 11160 12216 11212
rect 13268 11160 13320 11212
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 19524 11160 19576 11212
rect 20904 11203 20956 11212
rect 7196 11092 7248 11144
rect 11060 11092 11112 11144
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 16028 11092 16080 11144
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 25136 11203 25188 11212
rect 25136 11169 25145 11203
rect 25145 11169 25179 11203
rect 25179 11169 25188 11203
rect 25136 11160 25188 11169
rect 21548 11092 21600 11144
rect 22008 11092 22060 11144
rect 23664 11092 23716 11144
rect 2504 11067 2556 11076
rect 2504 11033 2513 11067
rect 2513 11033 2547 11067
rect 2547 11033 2556 11067
rect 2504 11024 2556 11033
rect 4068 11024 4120 11076
rect 4528 11067 4580 11076
rect 4528 11033 4537 11067
rect 4537 11033 4571 11067
rect 4571 11033 4580 11067
rect 4528 11024 4580 11033
rect 10692 11024 10744 11076
rect 12532 11024 12584 11076
rect 16120 11067 16172 11076
rect 16120 11033 16129 11067
rect 16129 11033 16163 11067
rect 16163 11033 16172 11067
rect 16120 11024 16172 11033
rect 23940 11067 23992 11076
rect 23940 11033 23949 11067
rect 23949 11033 23983 11067
rect 23983 11033 23992 11067
rect 23940 11024 23992 11033
rect 24952 11092 25004 11144
rect 25320 11024 25372 11076
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 2320 10999 2372 11008
rect 2320 10965 2329 10999
rect 2329 10965 2363 10999
rect 2363 10965 2372 10999
rect 2320 10956 2372 10965
rect 9864 10999 9916 11008
rect 9864 10965 9873 10999
rect 9873 10965 9907 10999
rect 9907 10965 9916 10999
rect 9864 10956 9916 10965
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12440 10956 12492 10965
rect 13636 10956 13688 11008
rect 16672 10956 16724 11008
rect 18972 10999 19024 11008
rect 18972 10965 18981 10999
rect 18981 10965 19015 10999
rect 19015 10965 19024 10999
rect 18972 10956 19024 10965
rect 22192 10956 22244 11008
rect 23848 10956 23900 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 2412 10752 2464 10804
rect 5448 10752 5500 10804
rect 6368 10752 6420 10804
rect 7196 10795 7248 10804
rect 7196 10761 7205 10795
rect 7205 10761 7239 10795
rect 7239 10761 7248 10795
rect 7196 10752 7248 10761
rect 7656 10795 7708 10804
rect 7656 10761 7665 10795
rect 7665 10761 7699 10795
rect 7699 10761 7708 10795
rect 7656 10752 7708 10761
rect 9404 10752 9456 10804
rect 10508 10795 10560 10804
rect 10508 10761 10517 10795
rect 10517 10761 10551 10795
rect 10551 10761 10560 10795
rect 10508 10752 10560 10761
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 11704 10752 11756 10804
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 12440 10752 12492 10804
rect 2504 10684 2556 10736
rect 2044 10548 2096 10600
rect 2320 10548 2372 10600
rect 5080 10616 5132 10668
rect 4528 10548 4580 10600
rect 4436 10480 4488 10532
rect 6920 10684 6972 10736
rect 8484 10684 8536 10736
rect 10968 10684 11020 10736
rect 7564 10616 7616 10668
rect 9036 10616 9088 10668
rect 12348 10684 12400 10736
rect 13820 10684 13872 10736
rect 14740 10684 14792 10736
rect 15384 10684 15436 10736
rect 13544 10616 13596 10668
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 10508 10548 10560 10600
rect 14372 10548 14424 10600
rect 16764 10752 16816 10804
rect 21548 10795 21600 10804
rect 21548 10761 21557 10795
rect 21557 10761 21591 10795
rect 21591 10761 21600 10795
rect 21548 10752 21600 10761
rect 25504 10795 25556 10804
rect 17592 10684 17644 10736
rect 20904 10684 20956 10736
rect 8024 10480 8076 10532
rect 9404 10480 9456 10532
rect 12532 10523 12584 10532
rect 12532 10489 12541 10523
rect 12541 10489 12575 10523
rect 12575 10489 12584 10523
rect 12532 10480 12584 10489
rect 12624 10523 12676 10532
rect 12624 10489 12633 10523
rect 12633 10489 12667 10523
rect 12667 10489 12676 10523
rect 12624 10480 12676 10489
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 4712 10412 4764 10464
rect 4896 10412 4948 10464
rect 6092 10412 6144 10464
rect 10140 10412 10192 10464
rect 14188 10455 14240 10464
rect 14188 10421 14197 10455
rect 14197 10421 14231 10455
rect 14231 10421 14240 10455
rect 14188 10412 14240 10421
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 16396 10548 16448 10600
rect 18420 10616 18472 10668
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 20352 10616 20404 10668
rect 25504 10761 25513 10795
rect 25513 10761 25547 10795
rect 25547 10761 25556 10795
rect 25504 10752 25556 10761
rect 23388 10684 23440 10736
rect 25596 10684 25648 10736
rect 17868 10548 17920 10557
rect 22192 10591 22244 10600
rect 15752 10480 15804 10532
rect 16948 10412 17000 10464
rect 18604 10480 18656 10532
rect 19432 10480 19484 10532
rect 18236 10412 18288 10464
rect 19524 10412 19576 10464
rect 22192 10557 22201 10591
rect 22201 10557 22235 10591
rect 22235 10557 22244 10591
rect 22192 10548 22244 10557
rect 22836 10616 22888 10668
rect 25136 10616 25188 10668
rect 23112 10548 23164 10600
rect 24400 10548 24452 10600
rect 21180 10523 21232 10532
rect 21180 10489 21189 10523
rect 21189 10489 21223 10523
rect 21223 10489 21232 10523
rect 21180 10480 21232 10489
rect 21272 10480 21324 10532
rect 23756 10523 23808 10532
rect 23756 10489 23765 10523
rect 23765 10489 23799 10523
rect 23799 10489 23808 10523
rect 23756 10480 23808 10489
rect 20720 10412 20772 10464
rect 22100 10455 22152 10464
rect 22100 10421 22109 10455
rect 22109 10421 22143 10455
rect 22143 10421 22152 10455
rect 22100 10412 22152 10421
rect 23020 10455 23072 10464
rect 23020 10421 23029 10455
rect 23029 10421 23063 10455
rect 23063 10421 23072 10455
rect 23020 10412 23072 10421
rect 23480 10412 23532 10464
rect 24952 10455 25004 10464
rect 24952 10421 24961 10455
rect 24961 10421 24995 10455
rect 24995 10421 25004 10455
rect 24952 10412 25004 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2872 10140 2924 10192
rect 2136 10072 2188 10124
rect 2320 10072 2372 10124
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 3792 10072 3844 10124
rect 4620 10208 4672 10260
rect 8024 10208 8076 10260
rect 11060 10208 11112 10260
rect 12624 10208 12676 10260
rect 13268 10208 13320 10260
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 15200 10208 15252 10260
rect 15660 10208 15712 10260
rect 17316 10208 17368 10260
rect 18420 10251 18472 10260
rect 18420 10217 18429 10251
rect 18429 10217 18463 10251
rect 18463 10217 18472 10251
rect 18420 10208 18472 10217
rect 18604 10208 18656 10260
rect 21180 10208 21232 10260
rect 21824 10208 21876 10260
rect 22284 10251 22336 10260
rect 22284 10217 22293 10251
rect 22293 10217 22327 10251
rect 22327 10217 22336 10251
rect 22284 10208 22336 10217
rect 4712 10072 4764 10124
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 8668 10140 8720 10192
rect 9312 10183 9364 10192
rect 9312 10149 9321 10183
rect 9321 10149 9355 10183
rect 9355 10149 9364 10183
rect 9312 10140 9364 10149
rect 10140 10140 10192 10192
rect 10692 10140 10744 10192
rect 13176 10183 13228 10192
rect 13176 10149 13185 10183
rect 13185 10149 13219 10183
rect 13219 10149 13228 10183
rect 13176 10140 13228 10149
rect 15568 10140 15620 10192
rect 17500 10183 17552 10192
rect 17500 10149 17509 10183
rect 17509 10149 17543 10183
rect 17543 10149 17552 10183
rect 17500 10140 17552 10149
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 6552 10072 6604 10124
rect 7196 10072 7248 10124
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 8392 10072 8444 10124
rect 11980 10115 12032 10124
rect 11980 10081 11989 10115
rect 11989 10081 12023 10115
rect 12023 10081 12032 10115
rect 11980 10072 12032 10081
rect 1952 10004 2004 10056
rect 4068 10004 4120 10056
rect 1400 9868 1452 9920
rect 1676 9868 1728 9920
rect 2412 9868 2464 9920
rect 3148 9868 3200 9920
rect 4896 9979 4948 9988
rect 4896 9945 4905 9979
rect 4905 9945 4939 9979
rect 4939 9945 4948 9979
rect 4896 9936 4948 9945
rect 6000 10004 6052 10056
rect 9036 10004 9088 10056
rect 7012 9936 7064 9988
rect 13452 10004 13504 10056
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 15384 10072 15436 10124
rect 16212 10072 16264 10124
rect 19340 10140 19392 10192
rect 19984 10072 20036 10124
rect 20352 10072 20404 10124
rect 20812 10115 20864 10124
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 21272 10140 21324 10192
rect 23572 10140 23624 10192
rect 23848 10183 23900 10192
rect 23848 10149 23857 10183
rect 23857 10149 23891 10183
rect 23891 10149 23900 10183
rect 23848 10140 23900 10149
rect 24400 10183 24452 10192
rect 24400 10149 24409 10183
rect 24409 10149 24443 10183
rect 24443 10149 24452 10183
rect 24400 10140 24452 10149
rect 22744 10072 22796 10124
rect 24860 10072 24912 10124
rect 26056 10072 26108 10124
rect 15844 10047 15896 10056
rect 13544 10004 13596 10013
rect 10692 9936 10744 9988
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 17684 10004 17736 10056
rect 18972 10004 19024 10056
rect 20444 10004 20496 10056
rect 21272 10004 21324 10056
rect 22100 10004 22152 10056
rect 23112 10004 23164 10056
rect 23940 10004 23992 10056
rect 15936 9936 15988 9988
rect 16856 9936 16908 9988
rect 19524 9936 19576 9988
rect 14556 9868 14608 9920
rect 16120 9868 16172 9920
rect 19248 9868 19300 9920
rect 20720 9868 20772 9920
rect 27528 9868 27580 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2228 9707 2280 9716
rect 2228 9673 2237 9707
rect 2237 9673 2271 9707
rect 2271 9673 2280 9707
rect 2228 9664 2280 9673
rect 2872 9664 2924 9716
rect 4712 9707 4764 9716
rect 4712 9673 4721 9707
rect 4721 9673 4755 9707
rect 4755 9673 4764 9707
rect 4712 9664 4764 9673
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 8024 9707 8076 9716
rect 8024 9673 8033 9707
rect 8033 9673 8067 9707
rect 8067 9673 8076 9707
rect 8024 9664 8076 9673
rect 8392 9707 8444 9716
rect 8392 9673 8401 9707
rect 8401 9673 8435 9707
rect 8435 9673 8444 9707
rect 8392 9664 8444 9673
rect 10140 9664 10192 9716
rect 1676 9596 1728 9648
rect 2136 9596 2188 9648
rect 1308 9528 1360 9580
rect 10968 9596 11020 9648
rect 2320 9528 2372 9580
rect 4896 9571 4948 9580
rect 2504 9460 2556 9512
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 5264 9528 5316 9580
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 9496 9528 9548 9580
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 13176 9664 13228 9716
rect 17500 9664 17552 9716
rect 18236 9707 18288 9716
rect 18236 9673 18245 9707
rect 18245 9673 18279 9707
rect 18279 9673 18288 9707
rect 18236 9664 18288 9673
rect 18696 9664 18748 9716
rect 19340 9664 19392 9716
rect 20168 9664 20220 9716
rect 20812 9664 20864 9716
rect 23020 9664 23072 9716
rect 23848 9664 23900 9716
rect 24860 9664 24912 9716
rect 25228 9664 25280 9716
rect 26056 9707 26108 9716
rect 26056 9673 26065 9707
rect 26065 9673 26099 9707
rect 26099 9673 26108 9707
rect 26056 9664 26108 9673
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 13544 9528 13596 9580
rect 4804 9503 4856 9512
rect 1860 9392 1912 9444
rect 1492 9324 1544 9376
rect 1676 9324 1728 9376
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 6920 9503 6972 9512
rect 6920 9469 6929 9503
rect 6929 9469 6963 9503
rect 6963 9469 6972 9503
rect 6920 9460 6972 9469
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 6552 9392 6604 9444
rect 8760 9435 8812 9444
rect 8760 9401 8769 9435
rect 8769 9401 8803 9435
rect 8803 9401 8812 9435
rect 9312 9435 9364 9444
rect 8760 9392 8812 9401
rect 9312 9401 9321 9435
rect 9321 9401 9355 9435
rect 9355 9401 9364 9435
rect 9312 9392 9364 9401
rect 13084 9435 13136 9444
rect 3240 9367 3292 9376
rect 3240 9333 3249 9367
rect 3249 9333 3283 9367
rect 3283 9333 3292 9367
rect 3240 9324 3292 9333
rect 3608 9324 3660 9376
rect 4436 9324 4488 9376
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7012 9324 7064 9333
rect 10140 9324 10192 9376
rect 13084 9401 13093 9435
rect 13093 9401 13127 9435
rect 13127 9401 13136 9435
rect 13084 9392 13136 9401
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 13452 9324 13504 9376
rect 20352 9596 20404 9648
rect 20904 9596 20956 9648
rect 23388 9596 23440 9648
rect 15384 9528 15436 9580
rect 19248 9571 19300 9580
rect 19248 9537 19257 9571
rect 19257 9537 19291 9571
rect 19291 9537 19300 9571
rect 19248 9528 19300 9537
rect 19432 9528 19484 9580
rect 20260 9528 20312 9580
rect 21824 9571 21876 9580
rect 21824 9537 21833 9571
rect 21833 9537 21867 9571
rect 21867 9537 21876 9571
rect 21824 9528 21876 9537
rect 14832 9460 14884 9512
rect 18512 9503 18564 9512
rect 18512 9469 18521 9503
rect 18521 9469 18555 9503
rect 18555 9469 18564 9503
rect 18512 9460 18564 9469
rect 19984 9460 20036 9512
rect 20628 9460 20680 9512
rect 21548 9503 21600 9512
rect 21548 9469 21557 9503
rect 21557 9469 21591 9503
rect 21591 9469 21600 9503
rect 25044 9596 25096 9648
rect 24216 9571 24268 9580
rect 24216 9537 24225 9571
rect 24225 9537 24259 9571
rect 24259 9537 24268 9571
rect 24216 9528 24268 9537
rect 21548 9460 21600 9469
rect 25688 9503 25740 9512
rect 25688 9469 25697 9503
rect 25697 9469 25731 9503
rect 25731 9469 25740 9503
rect 25688 9460 25740 9469
rect 15752 9392 15804 9444
rect 16120 9435 16172 9444
rect 16120 9401 16129 9435
rect 16129 9401 16163 9435
rect 16163 9401 16172 9435
rect 16120 9392 16172 9401
rect 16212 9435 16264 9444
rect 16212 9401 16221 9435
rect 16221 9401 16255 9435
rect 16255 9401 16264 9435
rect 16212 9392 16264 9401
rect 17316 9392 17368 9444
rect 15936 9367 15988 9376
rect 15936 9333 15945 9367
rect 15945 9333 15979 9367
rect 15979 9333 15988 9367
rect 15936 9324 15988 9333
rect 17684 9367 17736 9376
rect 17684 9333 17693 9367
rect 17693 9333 17727 9367
rect 17727 9333 17736 9367
rect 17684 9324 17736 9333
rect 19340 9435 19392 9444
rect 19340 9401 19349 9435
rect 19349 9401 19383 9435
rect 19383 9401 19392 9435
rect 19340 9392 19392 9401
rect 22008 9392 22060 9444
rect 20260 9324 20312 9376
rect 21824 9324 21876 9376
rect 22836 9392 22888 9444
rect 22284 9324 22336 9376
rect 23572 9324 23624 9376
rect 24676 9324 24728 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1676 9120 1728 9172
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2136 9120 2188 9172
rect 3608 9120 3660 9172
rect 3792 9163 3844 9172
rect 3792 9129 3801 9163
rect 3801 9129 3835 9163
rect 3835 9129 3844 9163
rect 3792 9120 3844 9129
rect 3976 9052 4028 9104
rect 4804 9120 4856 9172
rect 7932 9163 7984 9172
rect 7932 9129 7941 9163
rect 7941 9129 7975 9163
rect 7975 9129 7984 9163
rect 7932 9120 7984 9129
rect 10692 9163 10744 9172
rect 10692 9129 10701 9163
rect 10701 9129 10735 9163
rect 10735 9129 10744 9163
rect 10692 9120 10744 9129
rect 12348 9120 12400 9172
rect 13084 9120 13136 9172
rect 16028 9120 16080 9172
rect 16488 9120 16540 9172
rect 22100 9120 22152 9172
rect 4160 9052 4212 9104
rect 10048 9052 10100 9104
rect 16212 9052 16264 9104
rect 17040 9052 17092 9104
rect 17500 9052 17552 9104
rect 18788 9052 18840 9104
rect 21824 9052 21876 9104
rect 23572 9120 23624 9172
rect 24032 9120 24084 9172
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 4436 9027 4488 9036
rect 2688 8984 2740 8993
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 6092 9027 6144 9036
rect 6092 8993 6101 9027
rect 6101 8993 6135 9027
rect 6135 8993 6144 9027
rect 6092 8984 6144 8993
rect 6552 9027 6604 9036
rect 6552 8993 6561 9027
rect 6561 8993 6595 9027
rect 6595 8993 6604 9027
rect 6552 8984 6604 8993
rect 7472 8984 7524 9036
rect 13360 8984 13412 9036
rect 13912 8984 13964 9036
rect 16856 8984 16908 9036
rect 18604 9027 18656 9036
rect 18604 8993 18613 9027
rect 18613 8993 18647 9027
rect 18647 8993 18656 9027
rect 18604 8984 18656 8993
rect 19524 8984 19576 9036
rect 23112 8984 23164 9036
rect 23388 9027 23440 9036
rect 23388 8993 23397 9027
rect 23397 8993 23431 9027
rect 23431 8993 23440 9027
rect 23388 8984 23440 8993
rect 23848 9027 23900 9036
rect 23848 8993 23857 9027
rect 23857 8993 23891 9027
rect 23891 8993 23900 9027
rect 23848 8984 23900 8993
rect 25320 8984 25372 9036
rect 4712 8916 4764 8968
rect 8852 8916 8904 8968
rect 9220 8916 9272 8968
rect 3056 8848 3108 8900
rect 5356 8848 5408 8900
rect 9036 8848 9088 8900
rect 9404 8848 9456 8900
rect 11336 8916 11388 8968
rect 13176 8848 13228 8900
rect 13820 8848 13872 8900
rect 5264 8780 5316 8832
rect 6920 8780 6972 8832
rect 7472 8823 7524 8832
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 7472 8780 7524 8789
rect 8392 8780 8444 8832
rect 8760 8823 8812 8832
rect 8760 8789 8769 8823
rect 8769 8789 8803 8823
rect 8803 8789 8812 8823
rect 8760 8780 8812 8789
rect 9496 8780 9548 8832
rect 16120 8780 16172 8832
rect 16764 8916 16816 8968
rect 17316 8959 17368 8968
rect 17316 8925 17325 8959
rect 17325 8925 17359 8959
rect 17359 8925 17368 8959
rect 17316 8916 17368 8925
rect 20444 8916 20496 8968
rect 21364 8916 21416 8968
rect 21732 8916 21784 8968
rect 22008 8916 22060 8968
rect 22836 8959 22888 8968
rect 22836 8925 22845 8959
rect 22845 8925 22879 8959
rect 22879 8925 22888 8959
rect 22836 8916 22888 8925
rect 23296 8916 23348 8968
rect 23572 8916 23624 8968
rect 23664 8916 23716 8968
rect 24124 8916 24176 8968
rect 16856 8848 16908 8900
rect 17408 8848 17460 8900
rect 19340 8780 19392 8832
rect 21180 8823 21232 8832
rect 21180 8789 21189 8823
rect 21189 8789 21223 8823
rect 21223 8789 21232 8823
rect 21180 8780 21232 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 4068 8576 4120 8628
rect 6092 8619 6144 8628
rect 3240 8440 3292 8492
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 3056 8347 3108 8356
rect 3056 8313 3065 8347
rect 3065 8313 3099 8347
rect 3099 8313 3108 8347
rect 4528 8372 4580 8424
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 6552 8576 6604 8628
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 8760 8576 8812 8628
rect 8852 8619 8904 8628
rect 8852 8585 8861 8619
rect 8861 8585 8895 8619
rect 8895 8585 8904 8619
rect 8852 8576 8904 8585
rect 9036 8576 9088 8628
rect 12992 8576 13044 8628
rect 13268 8576 13320 8628
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 8208 8508 8260 8560
rect 9312 8508 9364 8560
rect 11796 8551 11848 8560
rect 11796 8517 11805 8551
rect 11805 8517 11839 8551
rect 11839 8517 11848 8551
rect 11796 8508 11848 8517
rect 13084 8508 13136 8560
rect 14372 8576 14424 8628
rect 15752 8576 15804 8628
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 19248 8576 19300 8628
rect 20260 8619 20312 8628
rect 20260 8585 20269 8619
rect 20269 8585 20303 8619
rect 20303 8585 20312 8619
rect 20260 8576 20312 8585
rect 20628 8576 20680 8628
rect 22836 8576 22888 8628
rect 23848 8576 23900 8628
rect 13912 8508 13964 8560
rect 5448 8415 5500 8424
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 3056 8304 3108 8313
rect 3608 8304 3660 8356
rect 9220 8372 9272 8424
rect 12256 8440 12308 8492
rect 14096 8440 14148 8492
rect 15108 8440 15160 8492
rect 15844 8440 15896 8492
rect 18604 8508 18656 8560
rect 20352 8508 20404 8560
rect 21180 8440 21232 8492
rect 23756 8440 23808 8492
rect 24216 8483 24268 8492
rect 24216 8449 24225 8483
rect 24225 8449 24259 8483
rect 24259 8449 24268 8483
rect 24216 8440 24268 8449
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 9404 8347 9456 8356
rect 9404 8313 9413 8347
rect 9413 8313 9447 8347
rect 9447 8313 9456 8347
rect 9404 8304 9456 8313
rect 2136 8236 2188 8288
rect 2688 8279 2740 8288
rect 2688 8245 2697 8279
rect 2697 8245 2731 8279
rect 2731 8245 2740 8279
rect 2688 8236 2740 8245
rect 4252 8236 4304 8288
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 7472 8236 7524 8245
rect 7932 8279 7984 8288
rect 7932 8245 7941 8279
rect 7941 8245 7975 8279
rect 7975 8245 7984 8279
rect 7932 8236 7984 8245
rect 9036 8236 9088 8288
rect 10140 8236 10192 8288
rect 11336 8236 11388 8288
rect 12348 8236 12400 8288
rect 12532 8236 12584 8288
rect 13728 8279 13780 8288
rect 13728 8245 13737 8279
rect 13737 8245 13771 8279
rect 13771 8245 13780 8279
rect 13728 8236 13780 8245
rect 14004 8304 14056 8356
rect 25044 8372 25096 8424
rect 19340 8347 19392 8356
rect 19340 8313 19349 8347
rect 19349 8313 19383 8347
rect 19383 8313 19392 8347
rect 19340 8304 19392 8313
rect 19524 8304 19576 8356
rect 19984 8304 20036 8356
rect 23388 8347 23440 8356
rect 14188 8236 14240 8288
rect 16120 8236 16172 8288
rect 16764 8236 16816 8288
rect 18144 8236 18196 8288
rect 18788 8236 18840 8288
rect 21548 8236 21600 8288
rect 21824 8236 21876 8288
rect 23388 8313 23397 8347
rect 23397 8313 23431 8347
rect 23431 8313 23440 8347
rect 23388 8304 23440 8313
rect 22744 8279 22796 8288
rect 22744 8245 22753 8279
rect 22753 8245 22787 8279
rect 22787 8245 22796 8279
rect 22744 8236 22796 8245
rect 23848 8347 23900 8356
rect 23848 8313 23857 8347
rect 23857 8313 23891 8347
rect 23891 8313 23900 8347
rect 23848 8304 23900 8313
rect 24032 8236 24084 8288
rect 25320 8236 25372 8288
rect 25780 8279 25832 8288
rect 25780 8245 25789 8279
rect 25789 8245 25823 8279
rect 25823 8245 25832 8279
rect 25780 8236 25832 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2412 8032 2464 8084
rect 3148 8075 3200 8084
rect 3148 8041 3157 8075
rect 3157 8041 3191 8075
rect 3191 8041 3200 8075
rect 3148 8032 3200 8041
rect 3240 8032 3292 8084
rect 2320 8007 2372 8016
rect 2320 7973 2329 8007
rect 2329 7973 2363 8007
rect 2363 7973 2372 8007
rect 2320 7964 2372 7973
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 6644 8007 6696 8016
rect 6644 7973 6653 8007
rect 6653 7973 6687 8007
rect 6687 7973 6696 8007
rect 6644 7964 6696 7973
rect 7472 7964 7524 8016
rect 7932 7964 7984 8016
rect 10140 7964 10192 8016
rect 12624 8032 12676 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 16120 8075 16172 8084
rect 16120 8041 16129 8075
rect 16129 8041 16163 8075
rect 16163 8041 16172 8075
rect 16120 8032 16172 8041
rect 17040 8032 17092 8084
rect 12532 7964 12584 8016
rect 13268 7964 13320 8016
rect 16764 7964 16816 8016
rect 16948 8007 17000 8016
rect 16948 7973 16951 8007
rect 16951 7973 16985 8007
rect 16985 7973 17000 8007
rect 16948 7964 17000 7973
rect 17316 7964 17368 8016
rect 8484 7939 8536 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2044 7760 2096 7812
rect 3332 7828 3384 7880
rect 4344 7828 4396 7880
rect 5448 7828 5500 7880
rect 6276 7828 6328 7880
rect 6736 7828 6788 7880
rect 8208 7828 8260 7880
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 12440 7896 12492 7948
rect 8392 7828 8444 7880
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 11244 7828 11296 7880
rect 14740 7828 14792 7880
rect 8024 7760 8076 7812
rect 9404 7803 9456 7812
rect 9404 7769 9413 7803
rect 9413 7769 9447 7803
rect 9447 7769 9456 7803
rect 9404 7760 9456 7769
rect 13176 7760 13228 7812
rect 14280 7803 14332 7812
rect 14280 7769 14289 7803
rect 14289 7769 14323 7803
rect 14323 7769 14332 7803
rect 14280 7760 14332 7769
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 3792 7692 3844 7744
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 5448 7692 5500 7701
rect 10048 7692 10100 7744
rect 12532 7692 12584 7744
rect 12992 7692 13044 7744
rect 16212 7896 16264 7948
rect 17408 7896 17460 7948
rect 19340 8075 19392 8084
rect 19340 8041 19349 8075
rect 19349 8041 19383 8075
rect 19383 8041 19392 8075
rect 19340 8032 19392 8041
rect 21824 7964 21876 8016
rect 18236 7896 18288 7948
rect 18420 7896 18472 7948
rect 22560 7828 22612 7880
rect 21732 7760 21784 7812
rect 23848 8032 23900 8084
rect 22744 7964 22796 8016
rect 23940 7964 23992 8016
rect 25596 7896 25648 7948
rect 25044 7828 25096 7880
rect 24216 7803 24268 7812
rect 24216 7769 24225 7803
rect 24225 7769 24259 7803
rect 24259 7769 24268 7803
rect 24216 7760 24268 7769
rect 21548 7692 21600 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1584 7488 1636 7540
rect 3976 7531 4028 7540
rect 3976 7497 3985 7531
rect 3985 7497 4019 7531
rect 4019 7497 4028 7531
rect 3976 7488 4028 7497
rect 4160 7488 4212 7540
rect 4344 7531 4396 7540
rect 4344 7497 4353 7531
rect 4353 7497 4387 7531
rect 4387 7497 4396 7531
rect 4344 7488 4396 7497
rect 6644 7488 6696 7540
rect 6736 7488 6788 7540
rect 2320 7420 2372 7472
rect 2044 7284 2096 7336
rect 3056 7352 3108 7404
rect 3792 7284 3844 7336
rect 3884 7284 3936 7336
rect 8392 7420 8444 7472
rect 4896 7352 4948 7404
rect 5448 7352 5500 7404
rect 7012 7327 7064 7336
rect 7012 7293 7021 7327
rect 7021 7293 7055 7327
rect 7055 7293 7064 7327
rect 7012 7284 7064 7293
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 9588 7488 9640 7540
rect 13268 7488 13320 7540
rect 14556 7488 14608 7540
rect 16212 7531 16264 7540
rect 9496 7420 9548 7472
rect 11612 7420 11664 7472
rect 9680 7352 9732 7404
rect 11060 7284 11112 7336
rect 12900 7284 12952 7336
rect 13636 7420 13688 7472
rect 14280 7463 14332 7472
rect 13268 7352 13320 7404
rect 14280 7429 14289 7463
rect 14289 7429 14323 7463
rect 14323 7429 14332 7463
rect 14280 7420 14332 7429
rect 16212 7497 16221 7531
rect 16221 7497 16255 7531
rect 16255 7497 16264 7531
rect 16212 7488 16264 7497
rect 17684 7488 17736 7540
rect 18512 7488 18564 7540
rect 20628 7488 20680 7540
rect 22836 7531 22888 7540
rect 22836 7497 22845 7531
rect 22845 7497 22879 7531
rect 22879 7497 22888 7531
rect 22836 7488 22888 7497
rect 25044 7531 25096 7540
rect 25044 7497 25053 7531
rect 25053 7497 25087 7531
rect 25087 7497 25096 7531
rect 25044 7488 25096 7497
rect 25596 7488 25648 7540
rect 17592 7420 17644 7472
rect 17776 7420 17828 7472
rect 15384 7352 15436 7404
rect 18420 7352 18472 7404
rect 19524 7352 19576 7404
rect 20812 7420 20864 7472
rect 21088 7420 21140 7472
rect 9588 7259 9640 7268
rect 9588 7225 9597 7259
rect 9597 7225 9631 7259
rect 9631 7225 9640 7259
rect 9588 7216 9640 7225
rect 2872 7148 2924 7200
rect 3332 7148 3384 7200
rect 4528 7148 4580 7200
rect 5356 7191 5408 7200
rect 5356 7157 5365 7191
rect 5365 7157 5399 7191
rect 5399 7157 5408 7191
rect 5356 7148 5408 7157
rect 6920 7191 6972 7200
rect 6920 7157 6929 7191
rect 6929 7157 6963 7191
rect 6963 7157 6972 7191
rect 6920 7148 6972 7157
rect 10048 7216 10100 7268
rect 13728 7259 13780 7268
rect 13728 7225 13737 7259
rect 13737 7225 13771 7259
rect 13771 7225 13780 7259
rect 13728 7216 13780 7225
rect 13820 7259 13872 7268
rect 13820 7225 13829 7259
rect 13829 7225 13863 7259
rect 13863 7225 13872 7259
rect 13820 7216 13872 7225
rect 14648 7216 14700 7268
rect 16764 7284 16816 7336
rect 16948 7327 17000 7336
rect 16948 7293 16992 7327
rect 16992 7293 17000 7327
rect 16948 7284 17000 7293
rect 20628 7327 20680 7336
rect 17316 7216 17368 7268
rect 18144 7216 18196 7268
rect 18788 7259 18840 7268
rect 18788 7225 18797 7259
rect 18797 7225 18831 7259
rect 18831 7225 18840 7259
rect 18788 7216 18840 7225
rect 19156 7216 19208 7268
rect 20260 7216 20312 7268
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 24952 7352 25004 7404
rect 20628 7284 20680 7293
rect 21180 7284 21232 7336
rect 22192 7284 22244 7336
rect 22836 7284 22888 7336
rect 23388 7284 23440 7336
rect 23480 7284 23532 7336
rect 10140 7148 10192 7200
rect 12532 7148 12584 7200
rect 12624 7148 12676 7200
rect 15476 7191 15528 7200
rect 15476 7157 15485 7191
rect 15485 7157 15519 7191
rect 15519 7157 15528 7191
rect 15476 7148 15528 7157
rect 17868 7148 17920 7200
rect 18236 7148 18288 7200
rect 21180 7191 21232 7200
rect 21180 7157 21189 7191
rect 21189 7157 21223 7191
rect 21223 7157 21232 7191
rect 21180 7148 21232 7157
rect 21364 7148 21416 7200
rect 21548 7191 21600 7200
rect 21548 7157 21557 7191
rect 21557 7157 21591 7191
rect 21591 7157 21600 7191
rect 21548 7148 21600 7157
rect 21732 7148 21784 7200
rect 23112 7216 23164 7268
rect 24124 7216 24176 7268
rect 22928 7148 22980 7200
rect 23388 7191 23440 7200
rect 23388 7157 23397 7191
rect 23397 7157 23431 7191
rect 23431 7157 23440 7191
rect 23388 7148 23440 7157
rect 23756 7191 23808 7200
rect 23756 7157 23765 7191
rect 23765 7157 23799 7191
rect 23799 7157 23808 7191
rect 23756 7148 23808 7157
rect 24768 7148 24820 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 2596 6944 2648 6996
rect 3056 6944 3108 6996
rect 3424 6987 3476 6996
rect 3424 6953 3433 6987
rect 3433 6953 3467 6987
rect 3467 6953 3476 6987
rect 3424 6944 3476 6953
rect 4160 6944 4212 6996
rect 4252 6944 4304 6996
rect 2228 6876 2280 6928
rect 2872 6876 2924 6928
rect 3148 6919 3200 6928
rect 3148 6885 3157 6919
rect 3157 6885 3191 6919
rect 3191 6885 3200 6919
rect 3148 6876 3200 6885
rect 4896 6919 4948 6928
rect 4896 6885 4905 6919
rect 4905 6885 4939 6919
rect 4939 6885 4948 6919
rect 4896 6876 4948 6885
rect 6276 6944 6328 6996
rect 7288 6944 7340 6996
rect 8852 6944 8904 6996
rect 9680 6944 9732 6996
rect 9864 6944 9916 6996
rect 6000 6919 6052 6928
rect 3884 6808 3936 6860
rect 4160 6851 4212 6860
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4712 6851 4764 6860
rect 4160 6808 4212 6817
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 6000 6885 6009 6919
rect 6009 6885 6043 6919
rect 6043 6885 6052 6919
rect 6000 6876 6052 6885
rect 7656 6919 7708 6928
rect 4712 6808 4764 6817
rect 5540 6808 5592 6860
rect 7656 6885 7665 6919
rect 7665 6885 7699 6919
rect 7699 6885 7708 6919
rect 7656 6876 7708 6885
rect 9588 6876 9640 6928
rect 12716 6919 12768 6928
rect 12716 6885 12725 6919
rect 12725 6885 12759 6919
rect 12759 6885 12768 6919
rect 12716 6876 12768 6885
rect 13268 6919 13320 6928
rect 13268 6885 13277 6919
rect 13277 6885 13311 6919
rect 13311 6885 13320 6919
rect 13268 6876 13320 6885
rect 13820 6944 13872 6996
rect 17224 6944 17276 6996
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 18236 6987 18288 6996
rect 18236 6953 18245 6987
rect 18245 6953 18279 6987
rect 18279 6953 18288 6987
rect 18236 6944 18288 6953
rect 18788 6987 18840 6996
rect 18788 6953 18797 6987
rect 18797 6953 18831 6987
rect 18831 6953 18840 6987
rect 18788 6944 18840 6953
rect 19524 6944 19576 6996
rect 20260 6987 20312 6996
rect 20260 6953 20269 6987
rect 20269 6953 20303 6987
rect 20303 6953 20312 6987
rect 20260 6944 20312 6953
rect 22560 6944 22612 6996
rect 23940 6944 23992 6996
rect 24952 6987 25004 6996
rect 24952 6953 24961 6987
rect 24961 6953 24995 6987
rect 24995 6953 25004 6987
rect 24952 6944 25004 6953
rect 17868 6876 17920 6928
rect 21364 6876 21416 6928
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 2596 6740 2648 6792
rect 2872 6740 2924 6792
rect 4896 6672 4948 6724
rect 6828 6740 6880 6792
rect 7196 6740 7248 6792
rect 9956 6740 10008 6792
rect 14556 6808 14608 6860
rect 15384 6808 15436 6860
rect 16764 6851 16816 6860
rect 11520 6740 11572 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 16212 6740 16264 6792
rect 16764 6817 16773 6851
rect 16773 6817 16807 6851
rect 16807 6817 16816 6851
rect 16764 6808 16816 6817
rect 19064 6808 19116 6860
rect 19616 6851 19668 6860
rect 19616 6817 19660 6851
rect 19660 6817 19668 6851
rect 19616 6808 19668 6817
rect 18420 6740 18472 6792
rect 22284 6740 22336 6792
rect 8024 6672 8076 6724
rect 8484 6672 8536 6724
rect 11428 6672 11480 6724
rect 16948 6672 17000 6724
rect 24032 6919 24084 6928
rect 24032 6885 24041 6919
rect 24041 6885 24075 6919
rect 24075 6885 24084 6919
rect 24032 6876 24084 6885
rect 24860 6876 24912 6928
rect 25136 6851 25188 6860
rect 25136 6817 25145 6851
rect 25145 6817 25179 6851
rect 25179 6817 25188 6851
rect 25136 6808 25188 6817
rect 25412 6851 25464 6860
rect 25412 6817 25421 6851
rect 25421 6817 25455 6851
rect 25455 6817 25464 6851
rect 25412 6808 25464 6817
rect 23204 6740 23256 6792
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2412 6604 2464 6656
rect 2688 6647 2740 6656
rect 2688 6613 2697 6647
rect 2697 6613 2731 6647
rect 2731 6613 2740 6647
rect 2688 6604 2740 6613
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 11244 6604 11296 6656
rect 13820 6604 13872 6656
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 16488 6604 16540 6656
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 21548 6604 21600 6656
rect 23756 6604 23808 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2688 6400 2740 6452
rect 4160 6400 4212 6452
rect 5540 6400 5592 6452
rect 7196 6400 7248 6452
rect 7656 6400 7708 6452
rect 8576 6400 8628 6452
rect 10140 6400 10192 6452
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 12716 6400 12768 6452
rect 16212 6400 16264 6452
rect 17132 6400 17184 6452
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 23296 6400 23348 6452
rect 23572 6400 23624 6452
rect 27620 6400 27672 6452
rect 4712 6375 4764 6384
rect 4712 6341 4721 6375
rect 4721 6341 4755 6375
rect 4755 6341 4764 6375
rect 4712 6332 4764 6341
rect 5080 6332 5132 6384
rect 5356 6332 5408 6384
rect 6000 6332 6052 6384
rect 7472 6332 7524 6384
rect 9404 6375 9456 6384
rect 9404 6341 9413 6375
rect 9413 6341 9447 6375
rect 9447 6341 9456 6375
rect 9404 6332 9456 6341
rect 9864 6332 9916 6384
rect 14372 6375 14424 6384
rect 2044 6239 2096 6248
rect 2044 6205 2053 6239
rect 2053 6205 2087 6239
rect 2087 6205 2096 6239
rect 2044 6196 2096 6205
rect 3792 6307 3844 6316
rect 3792 6273 3801 6307
rect 3801 6273 3835 6307
rect 3835 6273 3844 6307
rect 4896 6307 4948 6316
rect 3792 6264 3844 6273
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 7288 6264 7340 6316
rect 4068 6196 4120 6248
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 8208 6264 8260 6316
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 9496 6239 9548 6248
rect 5540 6196 5592 6205
rect 9496 6205 9505 6239
rect 9505 6205 9539 6239
rect 9539 6205 9548 6239
rect 9496 6196 9548 6205
rect 14372 6341 14381 6375
rect 14381 6341 14415 6375
rect 14415 6341 14424 6375
rect 14372 6332 14424 6341
rect 14740 6332 14792 6384
rect 24768 6332 24820 6384
rect 25136 6332 25188 6384
rect 26608 6332 26660 6384
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 15200 6307 15252 6316
rect 13820 6264 13872 6273
rect 15200 6273 15209 6307
rect 15209 6273 15243 6307
rect 15243 6273 15252 6307
rect 15200 6264 15252 6273
rect 16488 6264 16540 6316
rect 17776 6264 17828 6316
rect 23480 6264 23532 6316
rect 24032 6264 24084 6316
rect 13176 6239 13228 6248
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 14556 6196 14608 6248
rect 17868 6196 17920 6248
rect 18236 6196 18288 6248
rect 2596 6128 2648 6180
rect 3792 6128 3844 6180
rect 3976 6128 4028 6180
rect 5172 6128 5224 6180
rect 2872 6060 2924 6112
rect 8024 6128 8076 6180
rect 11244 6128 11296 6180
rect 12992 6128 13044 6180
rect 7932 6060 7984 6112
rect 9956 6060 10008 6112
rect 13084 6060 13136 6112
rect 15752 6128 15804 6180
rect 16212 6128 16264 6180
rect 16764 6171 16816 6180
rect 16764 6137 16773 6171
rect 16773 6137 16807 6171
rect 16807 6137 16816 6171
rect 19432 6196 19484 6248
rect 19616 6239 19668 6248
rect 19616 6205 19625 6239
rect 19625 6205 19659 6239
rect 19659 6205 19668 6239
rect 19616 6196 19668 6205
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 20352 6239 20404 6248
rect 20352 6205 20361 6239
rect 20361 6205 20395 6239
rect 20395 6205 20404 6239
rect 20352 6196 20404 6205
rect 21548 6239 21600 6248
rect 21548 6205 21557 6239
rect 21557 6205 21591 6239
rect 21591 6205 21600 6239
rect 21548 6196 21600 6205
rect 23296 6196 23348 6248
rect 23572 6196 23624 6248
rect 24124 6239 24176 6248
rect 24124 6205 24133 6239
rect 24133 6205 24167 6239
rect 24167 6205 24176 6239
rect 24124 6196 24176 6205
rect 16764 6128 16816 6137
rect 17868 6103 17920 6112
rect 17868 6069 17877 6103
rect 17877 6069 17911 6103
rect 17911 6069 17920 6103
rect 17868 6060 17920 6069
rect 19064 6103 19116 6112
rect 19064 6069 19073 6103
rect 19073 6069 19107 6103
rect 19107 6069 19116 6103
rect 19064 6060 19116 6069
rect 19432 6060 19484 6112
rect 21088 6060 21140 6112
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 22468 6103 22520 6112
rect 21364 6060 21416 6069
rect 22468 6069 22477 6103
rect 22477 6069 22511 6103
rect 22511 6069 22520 6103
rect 22468 6060 22520 6069
rect 23756 6103 23808 6112
rect 23756 6069 23765 6103
rect 23765 6069 23799 6103
rect 23799 6069 23808 6103
rect 23756 6060 23808 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2964 5856 3016 5908
rect 3332 5856 3384 5908
rect 5080 5856 5132 5908
rect 5172 5856 5224 5908
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 7196 5856 7248 5908
rect 7472 5856 7524 5908
rect 7932 5899 7984 5908
rect 7932 5865 7941 5899
rect 7941 5865 7975 5899
rect 7975 5865 7984 5899
rect 7932 5856 7984 5865
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 13084 5856 13136 5908
rect 3608 5788 3660 5840
rect 4804 5788 4856 5840
rect 9956 5788 10008 5840
rect 11060 5831 11112 5840
rect 664 5720 716 5772
rect 1676 5720 1728 5772
rect 2320 5720 2372 5772
rect 3332 5720 3384 5772
rect 3884 5720 3936 5772
rect 9036 5720 9088 5772
rect 2596 5652 2648 5704
rect 2320 5627 2372 5636
rect 2320 5593 2329 5627
rect 2329 5593 2363 5627
rect 2363 5593 2372 5627
rect 2320 5584 2372 5593
rect 2044 5516 2096 5568
rect 2872 5584 2924 5636
rect 3608 5584 3660 5636
rect 2964 5516 3016 5568
rect 3332 5516 3384 5568
rect 3976 5652 4028 5704
rect 6276 5652 6328 5704
rect 8668 5652 8720 5704
rect 11060 5797 11069 5831
rect 11069 5797 11103 5831
rect 11103 5797 11112 5831
rect 11060 5788 11112 5797
rect 14004 5856 14056 5908
rect 14556 5856 14608 5908
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 18420 5899 18472 5908
rect 18420 5865 18429 5899
rect 18429 5865 18463 5899
rect 18463 5865 18472 5899
rect 18420 5856 18472 5865
rect 13820 5831 13872 5840
rect 13820 5797 13829 5831
rect 13829 5797 13863 5831
rect 13863 5797 13872 5831
rect 14372 5831 14424 5840
rect 13820 5788 13872 5797
rect 14372 5797 14381 5831
rect 14381 5797 14415 5831
rect 14415 5797 14424 5831
rect 14372 5788 14424 5797
rect 17224 5831 17276 5840
rect 17224 5797 17233 5831
rect 17233 5797 17267 5831
rect 17267 5797 17276 5831
rect 17224 5788 17276 5797
rect 12348 5763 12400 5772
rect 12348 5729 12357 5763
rect 12357 5729 12391 5763
rect 12391 5729 12400 5763
rect 12348 5720 12400 5729
rect 12532 5763 12584 5772
rect 12532 5729 12541 5763
rect 12541 5729 12575 5763
rect 12575 5729 12584 5763
rect 12532 5720 12584 5729
rect 12624 5720 12676 5772
rect 10876 5652 10928 5704
rect 9680 5584 9732 5636
rect 14832 5652 14884 5704
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 21548 5856 21600 5908
rect 19064 5831 19116 5840
rect 19064 5797 19073 5831
rect 19073 5797 19107 5831
rect 19107 5797 19116 5831
rect 19064 5788 19116 5797
rect 19616 5788 19668 5840
rect 19984 5831 20036 5840
rect 19984 5797 19993 5831
rect 19993 5797 20027 5831
rect 20027 5797 20036 5831
rect 19984 5788 20036 5797
rect 20352 5831 20404 5840
rect 20352 5797 20361 5831
rect 20361 5797 20395 5831
rect 20395 5797 20404 5831
rect 22284 5831 22336 5840
rect 20352 5788 20404 5797
rect 22284 5797 22293 5831
rect 22293 5797 22327 5831
rect 22327 5797 22336 5831
rect 22284 5788 22336 5797
rect 22468 5788 22520 5840
rect 23940 5788 23992 5840
rect 18972 5695 19024 5704
rect 14740 5627 14792 5636
rect 14740 5593 14749 5627
rect 14749 5593 14783 5627
rect 14783 5593 14792 5627
rect 18972 5661 18981 5695
rect 18981 5661 19015 5695
rect 19015 5661 19024 5695
rect 18972 5652 19024 5661
rect 17684 5627 17736 5636
rect 14740 5584 14792 5593
rect 17684 5593 17693 5627
rect 17693 5593 17727 5627
rect 17727 5593 17736 5627
rect 17684 5584 17736 5593
rect 19156 5584 19208 5636
rect 19432 5652 19484 5704
rect 20720 5652 20772 5704
rect 21272 5720 21324 5772
rect 23572 5720 23624 5772
rect 24124 5763 24176 5772
rect 24124 5729 24133 5763
rect 24133 5729 24167 5763
rect 24167 5729 24176 5763
rect 24124 5720 24176 5729
rect 22192 5652 22244 5704
rect 22652 5695 22704 5704
rect 22652 5661 22661 5695
rect 22661 5661 22695 5695
rect 22695 5661 22704 5695
rect 22652 5652 22704 5661
rect 22744 5584 22796 5636
rect 4068 5516 4120 5568
rect 5356 5516 5408 5568
rect 10508 5559 10560 5568
rect 10508 5525 10532 5559
rect 10532 5525 10560 5559
rect 10508 5516 10560 5525
rect 10692 5516 10744 5568
rect 17868 5516 17920 5568
rect 22284 5516 22336 5568
rect 23572 5516 23624 5568
rect 23756 5559 23808 5568
rect 23756 5525 23765 5559
rect 23765 5525 23799 5559
rect 23799 5525 23808 5559
rect 23756 5516 23808 5525
rect 25136 5559 25188 5568
rect 25136 5525 25145 5559
rect 25145 5525 25179 5559
rect 25179 5525 25188 5559
rect 25136 5516 25188 5525
rect 25412 5516 25464 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2044 5312 2096 5364
rect 6276 5355 6328 5364
rect 2964 5244 3016 5296
rect 3700 5244 3752 5296
rect 1308 5176 1360 5228
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 4528 5244 4580 5296
rect 5080 5244 5132 5296
rect 6276 5321 6285 5355
rect 6285 5321 6319 5355
rect 6319 5321 6328 5355
rect 6276 5312 6328 5321
rect 9680 5355 9732 5364
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 9956 5355 10008 5364
rect 9956 5321 9965 5355
rect 9965 5321 9999 5355
rect 9999 5321 10008 5355
rect 9956 5312 10008 5321
rect 10508 5312 10560 5364
rect 10692 5312 10744 5364
rect 11152 5355 11204 5364
rect 11152 5321 11161 5355
rect 11161 5321 11195 5355
rect 11195 5321 11204 5355
rect 11152 5312 11204 5321
rect 7472 5244 7524 5296
rect 9496 5244 9548 5296
rect 11060 5244 11112 5296
rect 5356 5176 5408 5228
rect 6920 5176 6972 5228
rect 2320 5108 2372 5160
rect 3056 5108 3108 5160
rect 3700 5108 3752 5160
rect 2412 5040 2464 5092
rect 2780 5040 2832 5092
rect 3976 5040 4028 5092
rect 4712 5108 4764 5160
rect 6092 5108 6144 5160
rect 2872 4972 2924 5024
rect 2964 4972 3016 5024
rect 4896 5040 4948 5092
rect 5172 5040 5224 5092
rect 5632 5040 5684 5092
rect 8852 5108 8904 5160
rect 10140 5108 10192 5160
rect 10600 5108 10652 5160
rect 10876 5219 10928 5228
rect 10876 5185 10885 5219
rect 10885 5185 10919 5219
rect 10919 5185 10928 5219
rect 10876 5176 10928 5185
rect 12348 5312 12400 5364
rect 12532 5312 12584 5364
rect 14648 5312 14700 5364
rect 15752 5312 15804 5364
rect 17224 5355 17276 5364
rect 17224 5321 17233 5355
rect 17233 5321 17267 5355
rect 17267 5321 17276 5355
rect 17224 5312 17276 5321
rect 18972 5312 19024 5364
rect 19616 5355 19668 5364
rect 19616 5321 19625 5355
rect 19625 5321 19659 5355
rect 19659 5321 19668 5355
rect 19616 5312 19668 5321
rect 21088 5355 21140 5364
rect 21088 5321 21097 5355
rect 21097 5321 21131 5355
rect 21131 5321 21140 5355
rect 21088 5312 21140 5321
rect 22192 5312 22244 5364
rect 12808 5244 12860 5296
rect 18144 5244 18196 5296
rect 14740 5176 14792 5228
rect 15476 5176 15528 5228
rect 22376 5244 22428 5296
rect 22652 5312 22704 5364
rect 23388 5355 23440 5364
rect 23388 5321 23397 5355
rect 23397 5321 23431 5355
rect 23431 5321 23440 5355
rect 23388 5312 23440 5321
rect 24124 5312 24176 5364
rect 24768 5244 24820 5296
rect 19248 5176 19300 5228
rect 10692 5040 10744 5092
rect 11520 5083 11572 5092
rect 11520 5049 11529 5083
rect 11529 5049 11563 5083
rect 11563 5049 11572 5083
rect 11520 5040 11572 5049
rect 22744 5108 22796 5160
rect 23388 5108 23440 5160
rect 23756 5108 23808 5160
rect 24124 5151 24176 5160
rect 24124 5117 24133 5151
rect 24133 5117 24167 5151
rect 24167 5117 24176 5151
rect 24124 5108 24176 5117
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 7196 5015 7248 5024
rect 7196 4981 7205 5015
rect 7205 4981 7239 5015
rect 7239 4981 7248 5015
rect 7196 4972 7248 4981
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 8024 5015 8076 5024
rect 8024 4981 8033 5015
rect 8033 4981 8067 5015
rect 8067 4981 8076 5015
rect 8024 4972 8076 4981
rect 8668 5015 8720 5024
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 13452 5015 13504 5024
rect 13452 4981 13461 5015
rect 13461 4981 13495 5015
rect 13495 4981 13504 5015
rect 13452 4972 13504 4981
rect 15660 4972 15712 5024
rect 16580 5015 16632 5024
rect 16580 4981 16589 5015
rect 16589 4981 16623 5015
rect 16623 4981 16632 5015
rect 16580 4972 16632 4981
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 19064 5040 19116 5092
rect 21088 5040 21140 5092
rect 22100 5015 22152 5024
rect 17776 4972 17828 4981
rect 22100 4981 22109 5015
rect 22109 4981 22143 5015
rect 22143 4981 22152 5015
rect 22100 4972 22152 4981
rect 23572 4972 23624 5024
rect 25412 5015 25464 5024
rect 25412 4981 25421 5015
rect 25421 4981 25455 5015
rect 25455 4981 25464 5015
rect 25412 4972 25464 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 2228 4768 2280 4820
rect 2964 4768 3016 4820
rect 3608 4768 3660 4820
rect 3700 4768 3752 4820
rect 3884 4768 3936 4820
rect 4712 4811 4764 4820
rect 4712 4777 4721 4811
rect 4721 4777 4755 4811
rect 4755 4777 4764 4811
rect 4712 4768 4764 4777
rect 6460 4811 6512 4820
rect 6460 4777 6469 4811
rect 6469 4777 6503 4811
rect 6503 4777 6512 4811
rect 6460 4768 6512 4777
rect 7196 4768 7248 4820
rect 1676 4700 1728 4752
rect 3240 4700 3292 4752
rect 4068 4700 4120 4752
rect 5080 4743 5132 4752
rect 5080 4709 5089 4743
rect 5089 4709 5123 4743
rect 5123 4709 5132 4743
rect 5080 4700 5132 4709
rect 5632 4743 5684 4752
rect 5632 4709 5641 4743
rect 5641 4709 5675 4743
rect 5675 4709 5684 4743
rect 5632 4700 5684 4709
rect 7104 4700 7156 4752
rect 8852 4768 8904 4820
rect 8944 4768 8996 4820
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 13820 4768 13872 4820
rect 14832 4768 14884 4820
rect 7748 4700 7800 4752
rect 9036 4743 9088 4752
rect 9036 4709 9045 4743
rect 9045 4709 9079 4743
rect 9079 4709 9088 4743
rect 9036 4700 9088 4709
rect 10968 4700 11020 4752
rect 11428 4700 11480 4752
rect 13636 4743 13688 4752
rect 2228 4632 2280 4684
rect 2412 4675 2464 4684
rect 2412 4641 2421 4675
rect 2421 4641 2455 4675
rect 2455 4641 2464 4675
rect 2412 4632 2464 4641
rect 3332 4632 3384 4684
rect 9864 4632 9916 4684
rect 2044 4564 2096 4616
rect 2780 4607 2832 4616
rect 2780 4573 2789 4607
rect 2789 4573 2823 4607
rect 2823 4573 2832 4607
rect 2780 4564 2832 4573
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 2688 4539 2740 4548
rect 2688 4505 2697 4539
rect 2697 4505 2731 4539
rect 2731 4505 2740 4539
rect 2688 4496 2740 4505
rect 4712 4496 4764 4548
rect 8024 4564 8076 4616
rect 9772 4564 9824 4616
rect 11612 4632 11664 4684
rect 13636 4709 13645 4743
rect 13645 4709 13679 4743
rect 13679 4709 13688 4743
rect 13636 4700 13688 4709
rect 14372 4700 14424 4752
rect 17132 4768 17184 4820
rect 18144 4811 18196 4820
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 18328 4768 18380 4820
rect 21272 4768 21324 4820
rect 16120 4700 16172 4752
rect 16580 4700 16632 4752
rect 17684 4700 17736 4752
rect 17776 4700 17828 4752
rect 20720 4700 20772 4752
rect 21088 4700 21140 4752
rect 12164 4632 12216 4684
rect 19708 4632 19760 4684
rect 20996 4632 21048 4684
rect 22468 4768 22520 4820
rect 22744 4768 22796 4820
rect 22100 4700 22152 4752
rect 22652 4700 22704 4752
rect 23940 4700 23992 4752
rect 24124 4743 24176 4752
rect 24124 4709 24133 4743
rect 24133 4709 24167 4743
rect 24167 4709 24176 4743
rect 24124 4700 24176 4709
rect 22560 4632 22612 4684
rect 23848 4632 23900 4684
rect 24676 4632 24728 4684
rect 2504 4428 2556 4480
rect 9312 4428 9364 4480
rect 10784 4428 10836 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 12256 4471 12308 4480
rect 12256 4437 12265 4471
rect 12265 4437 12299 4471
rect 12299 4437 12308 4471
rect 12256 4428 12308 4437
rect 13268 4471 13320 4480
rect 13268 4437 13277 4471
rect 13277 4437 13311 4471
rect 13311 4437 13320 4471
rect 16212 4564 16264 4616
rect 18328 4607 18380 4616
rect 18328 4573 18337 4607
rect 18337 4573 18371 4607
rect 18371 4573 18380 4607
rect 18328 4564 18380 4573
rect 18972 4607 19024 4616
rect 18972 4573 18981 4607
rect 18981 4573 19015 4607
rect 19015 4573 19024 4607
rect 18972 4564 19024 4573
rect 21088 4607 21140 4616
rect 21088 4573 21097 4607
rect 21097 4573 21131 4607
rect 21131 4573 21140 4607
rect 21088 4564 21140 4573
rect 22928 4607 22980 4616
rect 22928 4573 22937 4607
rect 22937 4573 22971 4607
rect 22971 4573 22980 4607
rect 22928 4564 22980 4573
rect 18236 4496 18288 4548
rect 20352 4496 20404 4548
rect 15660 4471 15712 4480
rect 13268 4428 13320 4437
rect 15660 4437 15669 4471
rect 15669 4437 15703 4471
rect 15703 4437 15712 4471
rect 15660 4428 15712 4437
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 20076 4428 20128 4480
rect 22008 4471 22060 4480
rect 22008 4437 22017 4471
rect 22017 4437 22051 4471
rect 22051 4437 22060 4471
rect 22008 4428 22060 4437
rect 25136 4428 25188 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2780 4156 2832 4208
rect 1952 4020 2004 4072
rect 4804 4088 4856 4140
rect 5540 4156 5592 4208
rect 6000 4088 6052 4140
rect 6460 4088 6512 4140
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 3976 4063 4028 4072
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 7748 4224 7800 4276
rect 9588 4267 9640 4276
rect 9588 4233 9597 4267
rect 9597 4233 9631 4267
rect 9631 4233 9640 4267
rect 9588 4224 9640 4233
rect 10140 4224 10192 4276
rect 10600 4224 10652 4276
rect 11612 4224 11664 4276
rect 12164 4267 12216 4276
rect 12164 4233 12173 4267
rect 12173 4233 12207 4267
rect 12207 4233 12216 4267
rect 12164 4224 12216 4233
rect 15936 4224 15988 4276
rect 16120 4267 16172 4276
rect 16120 4233 16129 4267
rect 16129 4233 16163 4267
rect 16163 4233 16172 4267
rect 16120 4224 16172 4233
rect 17776 4224 17828 4276
rect 19432 4224 19484 4276
rect 9864 4156 9916 4208
rect 11520 4199 11572 4208
rect 11520 4165 11529 4199
rect 11529 4165 11563 4199
rect 11563 4165 11572 4199
rect 11520 4156 11572 4165
rect 14372 4156 14424 4208
rect 16212 4156 16264 4208
rect 19064 4156 19116 4208
rect 19708 4199 19760 4208
rect 7840 4088 7892 4140
rect 10140 4131 10192 4140
rect 8116 4020 8168 4072
rect 9312 4020 9364 4072
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 11152 4020 11204 4072
rect 3332 3995 3384 4004
rect 3332 3961 3341 3995
rect 3341 3961 3375 3995
rect 3375 3961 3384 3995
rect 3332 3952 3384 3961
rect 4160 3995 4212 4004
rect 4160 3961 4169 3995
rect 4169 3961 4203 3995
rect 4203 3961 4212 3995
rect 4160 3952 4212 3961
rect 5172 3995 5224 4004
rect 5172 3961 5181 3995
rect 5181 3961 5215 3995
rect 5215 3961 5224 3995
rect 5172 3952 5224 3961
rect 7012 3995 7064 4004
rect 7012 3961 7021 3995
rect 7021 3961 7055 3995
rect 7055 3961 7064 3995
rect 7012 3952 7064 3961
rect 7104 3952 7156 4004
rect 7656 3952 7708 4004
rect 8944 3995 8996 4004
rect 2136 3884 2188 3936
rect 4988 3884 5040 3936
rect 5080 3884 5132 3936
rect 8300 3927 8352 3936
rect 8300 3893 8309 3927
rect 8309 3893 8343 3927
rect 8343 3893 8352 3927
rect 8944 3961 8953 3995
rect 8953 3961 8987 3995
rect 8987 3961 8996 3995
rect 8944 3952 8996 3961
rect 9496 3952 9548 4004
rect 10784 3927 10836 3936
rect 8300 3884 8352 3893
rect 10784 3893 10793 3927
rect 10793 3893 10827 3927
rect 10827 3893 10836 3927
rect 10784 3884 10836 3893
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 13636 3884 13688 3936
rect 17500 4088 17552 4140
rect 17868 4088 17920 4140
rect 19708 4165 19717 4199
rect 19717 4165 19751 4199
rect 19751 4165 19760 4199
rect 19708 4156 19760 4165
rect 16580 3995 16632 4004
rect 16580 3961 16589 3995
rect 16589 3961 16623 3995
rect 16623 3961 16632 3995
rect 16580 3952 16632 3961
rect 17960 4020 18012 4072
rect 18144 4020 18196 4072
rect 19432 4088 19484 4140
rect 20076 4088 20128 4140
rect 22008 4224 22060 4276
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 23940 4156 23992 4208
rect 24860 4156 24912 4208
rect 22468 4088 22520 4140
rect 22928 4088 22980 4140
rect 25780 4131 25832 4140
rect 23204 4020 23256 4072
rect 24124 4020 24176 4072
rect 25780 4097 25789 4131
rect 25789 4097 25823 4131
rect 25823 4097 25832 4131
rect 25780 4088 25832 4097
rect 19892 3995 19944 4004
rect 17868 3927 17920 3936
rect 17868 3893 17877 3927
rect 17877 3893 17911 3927
rect 17911 3893 17920 3927
rect 17868 3884 17920 3893
rect 18052 3884 18104 3936
rect 19892 3961 19901 3995
rect 19901 3961 19935 3995
rect 19935 3961 19944 3995
rect 19892 3952 19944 3961
rect 20076 3952 20128 4004
rect 21456 3952 21508 4004
rect 22008 3995 22060 4004
rect 22008 3961 22017 3995
rect 22017 3961 22051 3995
rect 22051 3961 22060 3995
rect 22008 3952 22060 3961
rect 22100 3995 22152 4004
rect 22100 3961 22109 3995
rect 22109 3961 22143 3995
rect 22143 3961 22152 3995
rect 22100 3952 22152 3961
rect 20720 3884 20772 3936
rect 20996 3884 21048 3936
rect 22192 3884 22244 3936
rect 23756 3927 23808 3936
rect 23756 3893 23765 3927
rect 23765 3893 23799 3927
rect 23799 3893 23808 3927
rect 23756 3884 23808 3893
rect 25504 3884 25556 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2688 3723 2740 3732
rect 2688 3689 2697 3723
rect 2697 3689 2731 3723
rect 2731 3689 2740 3723
rect 2688 3680 2740 3689
rect 3700 3680 3752 3732
rect 4620 3680 4672 3732
rect 5080 3680 5132 3732
rect 3976 3612 4028 3664
rect 4528 3612 4580 3664
rect 4988 3612 5040 3664
rect 7012 3612 7064 3664
rect 7380 3655 7432 3664
rect 7380 3621 7389 3655
rect 7389 3621 7423 3655
rect 7423 3621 7432 3655
rect 7380 3612 7432 3621
rect 8208 3612 8260 3664
rect 8852 3680 8904 3732
rect 9680 3680 9732 3732
rect 10140 3680 10192 3732
rect 16396 3680 16448 3732
rect 18236 3680 18288 3732
rect 18788 3680 18840 3732
rect 20444 3680 20496 3732
rect 21088 3680 21140 3732
rect 22652 3723 22704 3732
rect 13820 3655 13872 3664
rect 13820 3621 13829 3655
rect 13829 3621 13863 3655
rect 13863 3621 13872 3655
rect 14372 3655 14424 3664
rect 13820 3612 13872 3621
rect 14372 3621 14381 3655
rect 14381 3621 14415 3655
rect 14415 3621 14424 3655
rect 14372 3612 14424 3621
rect 15476 3655 15528 3664
rect 15476 3621 15485 3655
rect 15485 3621 15519 3655
rect 15519 3621 15528 3655
rect 15476 3612 15528 3621
rect 16212 3612 16264 3664
rect 16580 3612 16632 3664
rect 18328 3612 18380 3664
rect 18972 3655 19024 3664
rect 18972 3621 18981 3655
rect 18981 3621 19015 3655
rect 19015 3621 19024 3655
rect 18972 3612 19024 3621
rect 112 3544 164 3596
rect 1676 3544 1728 3596
rect 2228 3476 2280 3528
rect 2872 3476 2924 3528
rect 4160 3544 4212 3596
rect 6092 3544 6144 3596
rect 10600 3587 10652 3596
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 9312 3476 9364 3528
rect 12256 3544 12308 3596
rect 16948 3544 17000 3596
rect 19248 3544 19300 3596
rect 19800 3587 19852 3596
rect 19800 3553 19809 3587
rect 19809 3553 19843 3587
rect 19843 3553 19852 3587
rect 19800 3544 19852 3553
rect 19984 3612 20036 3664
rect 21732 3612 21784 3664
rect 22652 3689 22661 3723
rect 22661 3689 22695 3723
rect 22695 3689 22704 3723
rect 22652 3680 22704 3689
rect 22744 3680 22796 3732
rect 23756 3612 23808 3664
rect 21456 3587 21508 3596
rect 21456 3553 21465 3587
rect 21465 3553 21499 3587
rect 21499 3553 21508 3587
rect 21456 3544 21508 3553
rect 22468 3544 22520 3596
rect 23296 3587 23348 3596
rect 23296 3553 23305 3587
rect 23305 3553 23339 3587
rect 23339 3553 23348 3587
rect 23296 3544 23348 3553
rect 11796 3476 11848 3528
rect 14464 3476 14516 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 19340 3476 19392 3528
rect 21824 3476 21876 3528
rect 2044 3340 2096 3392
rect 4896 3408 4948 3460
rect 6460 3408 6512 3460
rect 6552 3408 6604 3460
rect 9128 3408 9180 3460
rect 10232 3408 10284 3460
rect 6736 3340 6788 3392
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 9864 3340 9916 3392
rect 10416 3340 10468 3392
rect 10692 3340 10744 3392
rect 10876 3383 10928 3392
rect 10876 3349 10885 3383
rect 10885 3349 10919 3383
rect 10919 3349 10928 3383
rect 10876 3340 10928 3349
rect 10968 3340 11020 3392
rect 11520 3340 11572 3392
rect 13360 3383 13412 3392
rect 13360 3349 13369 3383
rect 13369 3349 13403 3383
rect 13403 3349 13412 3383
rect 13360 3340 13412 3349
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 22192 3408 22244 3460
rect 22560 3476 22612 3528
rect 24768 3544 24820 3596
rect 25044 3587 25096 3596
rect 25044 3553 25053 3587
rect 25053 3553 25087 3587
rect 25087 3553 25096 3587
rect 25044 3544 25096 3553
rect 25504 3544 25556 3596
rect 23756 3519 23808 3528
rect 23756 3485 23765 3519
rect 23765 3485 23799 3519
rect 23799 3485 23808 3519
rect 23756 3476 23808 3485
rect 20444 3340 20496 3392
rect 22652 3340 22704 3392
rect 23296 3340 23348 3392
rect 24032 3340 24084 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2872 3179 2924 3188
rect 2872 3145 2881 3179
rect 2881 3145 2915 3179
rect 2915 3145 2924 3179
rect 2872 3136 2924 3145
rect 3608 3136 3660 3188
rect 6552 3136 6604 3188
rect 7196 3136 7248 3188
rect 7380 3136 7432 3188
rect 4528 3111 4580 3120
rect 4528 3077 4537 3111
rect 4537 3077 4571 3111
rect 4571 3077 4580 3111
rect 4528 3068 4580 3077
rect 5540 3111 5592 3120
rect 5540 3077 5549 3111
rect 5549 3077 5583 3111
rect 5583 3077 5592 3111
rect 5540 3068 5592 3077
rect 6736 3068 6788 3120
rect 4344 3000 4396 3052
rect 4620 3000 4672 3052
rect 8024 3000 8076 3052
rect 8300 3000 8352 3052
rect 8852 3000 8904 3052
rect 2228 2975 2280 2984
rect 2228 2941 2237 2975
rect 2237 2941 2271 2975
rect 2271 2941 2280 2975
rect 2228 2932 2280 2941
rect 3424 2975 3476 2984
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 3608 2932 3660 2984
rect 7012 2932 7064 2984
rect 9404 3000 9456 3052
rect 9956 3136 10008 3188
rect 12256 3179 12308 3188
rect 9772 3068 9824 3120
rect 10416 3068 10468 3120
rect 12256 3145 12265 3179
rect 12265 3145 12299 3179
rect 12299 3145 12308 3179
rect 12256 3136 12308 3145
rect 13820 3136 13872 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 16488 3136 16540 3188
rect 16948 3136 17000 3188
rect 19800 3179 19852 3188
rect 19800 3145 19809 3179
rect 19809 3145 19843 3179
rect 19843 3145 19852 3179
rect 19800 3136 19852 3145
rect 21272 3136 21324 3188
rect 22652 3136 22704 3188
rect 22836 3179 22888 3188
rect 22836 3145 22845 3179
rect 22845 3145 22879 3179
rect 22879 3145 22888 3179
rect 22836 3136 22888 3145
rect 18420 3068 18472 3120
rect 22284 3068 22336 3120
rect 4804 2864 4856 2916
rect 5080 2907 5132 2916
rect 5080 2873 5089 2907
rect 5089 2873 5123 2907
rect 5123 2873 5132 2907
rect 5080 2864 5132 2873
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 2504 2796 2556 2848
rect 3240 2839 3292 2848
rect 3240 2805 3249 2839
rect 3249 2805 3283 2839
rect 3283 2805 3292 2839
rect 3240 2796 3292 2805
rect 6092 2796 6144 2848
rect 7196 2796 7248 2848
rect 9128 2975 9180 2984
rect 9128 2941 9137 2975
rect 9137 2941 9171 2975
rect 9171 2941 9180 2975
rect 9128 2932 9180 2941
rect 10232 2975 10284 2984
rect 10232 2941 10241 2975
rect 10241 2941 10275 2975
rect 10275 2941 10284 2975
rect 10232 2932 10284 2941
rect 16396 3043 16448 3052
rect 16396 3009 16405 3043
rect 16405 3009 16439 3043
rect 16439 3009 16448 3043
rect 16396 3000 16448 3009
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 18972 3000 19024 3052
rect 22744 3000 22796 3052
rect 23480 3136 23532 3188
rect 23664 3068 23716 3120
rect 25044 3179 25096 3188
rect 25044 3145 25053 3179
rect 25053 3145 25087 3179
rect 25087 3145 25096 3179
rect 25044 3136 25096 3145
rect 23940 3111 23992 3120
rect 23940 3077 23949 3111
rect 23949 3077 23983 3111
rect 23983 3077 23992 3111
rect 23940 3068 23992 3077
rect 24032 3043 24084 3052
rect 10876 2932 10928 2984
rect 11704 2932 11756 2984
rect 13360 2932 13412 2984
rect 14648 2932 14700 2984
rect 24032 3009 24041 3043
rect 24041 3009 24075 3043
rect 24075 3009 24084 3043
rect 24032 3000 24084 3009
rect 24124 3043 24176 3052
rect 24124 3009 24133 3043
rect 24133 3009 24167 3043
rect 24167 3009 24176 3043
rect 24124 3000 24176 3009
rect 23112 2932 23164 2984
rect 23848 2932 23900 2984
rect 9220 2864 9272 2916
rect 9864 2796 9916 2848
rect 11796 2796 11848 2848
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 15660 2864 15712 2916
rect 16212 2864 16264 2916
rect 16488 2907 16540 2916
rect 16488 2873 16497 2907
rect 16497 2873 16531 2907
rect 16531 2873 16540 2907
rect 16488 2864 16540 2873
rect 19248 2864 19300 2916
rect 20996 2864 21048 2916
rect 21272 2864 21324 2916
rect 17776 2839 17828 2848
rect 12624 2796 12676 2805
rect 17776 2805 17785 2839
rect 17785 2805 17819 2839
rect 17819 2805 17828 2839
rect 17776 2796 17828 2805
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 21732 2839 21784 2848
rect 21732 2805 21741 2839
rect 21741 2805 21775 2839
rect 21775 2805 21784 2839
rect 21732 2796 21784 2805
rect 23296 2796 23348 2848
rect 24216 2796 24268 2848
rect 25504 2796 25556 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 3608 2592 3660 2644
rect 4528 2592 4580 2644
rect 5172 2592 5224 2644
rect 6920 2592 6972 2644
rect 848 2456 900 2508
rect 6368 2524 6420 2576
rect 8024 2592 8076 2644
rect 7196 2524 7248 2576
rect 7656 2567 7708 2576
rect 7656 2533 7665 2567
rect 7665 2533 7699 2567
rect 7699 2533 7708 2567
rect 7656 2524 7708 2533
rect 4712 2456 4764 2508
rect 4804 2456 4856 2508
rect 11152 2524 11204 2576
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 4344 2388 4396 2440
rect 2136 2252 2188 2304
rect 9588 2456 9640 2508
rect 9680 2456 9732 2508
rect 11888 2592 11940 2644
rect 13636 2635 13688 2644
rect 13636 2601 13645 2635
rect 13645 2601 13679 2635
rect 13679 2601 13688 2635
rect 13636 2592 13688 2601
rect 16212 2592 16264 2644
rect 11704 2567 11756 2576
rect 11704 2533 11713 2567
rect 11713 2533 11747 2567
rect 11747 2533 11756 2567
rect 11704 2524 11756 2533
rect 12624 2524 12676 2576
rect 17776 2592 17828 2644
rect 18328 2592 18380 2644
rect 21272 2592 21324 2644
rect 21824 2592 21876 2644
rect 17868 2524 17920 2576
rect 21732 2524 21784 2576
rect 22008 2567 22060 2576
rect 22008 2533 22017 2567
rect 22017 2533 22051 2567
rect 22051 2533 22060 2567
rect 22008 2524 22060 2533
rect 11428 2499 11480 2508
rect 11428 2465 11437 2499
rect 11437 2465 11471 2499
rect 11471 2465 11480 2499
rect 11428 2456 11480 2465
rect 11520 2456 11572 2508
rect 18420 2456 18472 2508
rect 19156 2456 19208 2508
rect 23572 2456 23624 2508
rect 12164 2388 12216 2440
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 21364 2431 21416 2440
rect 21364 2397 21373 2431
rect 21373 2397 21407 2431
rect 21407 2397 21416 2431
rect 21364 2388 21416 2397
rect 21456 2388 21508 2440
rect 23940 2592 23992 2644
rect 24124 2635 24176 2644
rect 24124 2601 24133 2635
rect 24133 2601 24167 2635
rect 24167 2601 24176 2635
rect 24124 2592 24176 2601
rect 25504 2635 25556 2644
rect 25504 2601 25513 2635
rect 25513 2601 25547 2635
rect 25547 2601 25556 2635
rect 25504 2592 25556 2601
rect 24216 2499 24268 2508
rect 24216 2465 24225 2499
rect 24225 2465 24259 2499
rect 24259 2465 24268 2499
rect 24216 2456 24268 2465
rect 25320 2456 25372 2508
rect 9772 2320 9824 2372
rect 8760 2252 8812 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 10232 2320 10284 2372
rect 12624 2320 12676 2372
rect 13452 2320 13504 2372
rect 10692 2295 10744 2304
rect 10692 2261 10701 2295
rect 10701 2261 10735 2295
rect 10735 2261 10744 2295
rect 10692 2252 10744 2261
rect 11428 2252 11480 2304
rect 14648 2295 14700 2304
rect 14648 2261 14657 2295
rect 14657 2261 14691 2295
rect 14691 2261 14700 2295
rect 14648 2252 14700 2261
rect 22008 2320 22060 2372
rect 23112 2320 23164 2372
rect 27712 2252 27764 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 15384 2048 15436 2100
rect 23112 2048 23164 2100
rect 11980 76 12032 128
rect 16304 76 16356 128
rect 16764 76 16816 128
rect 17776 76 17828 128
<< metal2 >>
rect 662 27520 718 28000
rect 768 27526 1072 27554
rect 676 27418 704 27520
rect 768 27418 796 27526
rect 676 27390 796 27418
rect 1044 22642 1072 27526
rect 2042 27520 2098 28000
rect 3422 27554 3478 28000
rect 3068 27526 3478 27554
rect 1122 26752 1178 26761
rect 1122 26687 1178 26696
rect 1136 23322 1164 26687
rect 1582 25392 1638 25401
rect 1582 25327 1638 25336
rect 1214 24032 1270 24041
rect 1214 23967 1270 23976
rect 1124 23316 1176 23322
rect 1124 23258 1176 23264
rect 1228 22778 1256 23967
rect 1596 23866 1624 25327
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1952 23656 2004 23662
rect 1952 23598 2004 23604
rect 1964 23254 1992 23598
rect 1952 23248 2004 23254
rect 1952 23190 2004 23196
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1216 22772 1268 22778
rect 1216 22714 1268 22720
rect 1032 22636 1084 22642
rect 1032 22578 1084 22584
rect 1412 22234 1440 23122
rect 1952 22568 2004 22574
rect 1582 22536 1638 22545
rect 1952 22510 2004 22516
rect 1582 22471 1638 22480
rect 1400 22228 1452 22234
rect 1400 22170 1452 22176
rect 1596 21690 1624 22471
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 664 21480 716 21486
rect 664 21422 716 21428
rect 676 5778 704 21422
rect 1122 21176 1178 21185
rect 1122 21111 1178 21120
rect 1136 15706 1164 21111
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 1216 15904 1268 15910
rect 1216 15846 1268 15852
rect 1124 15700 1176 15706
rect 1124 15642 1176 15648
rect 1030 13152 1086 13161
rect 1030 13087 1086 13096
rect 1044 8265 1072 13087
rect 1030 8256 1086 8265
rect 1030 8191 1086 8200
rect 664 5772 716 5778
rect 664 5714 716 5720
rect 112 3596 164 3602
rect 112 3538 164 3544
rect 124 3505 152 3538
rect 110 3496 166 3505
rect 110 3431 166 3440
rect 1228 2689 1256 15846
rect 1412 15570 1440 20198
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1504 18630 1532 19858
rect 1582 19816 1638 19825
rect 1582 19751 1638 19760
rect 1596 19514 1624 19751
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 15094 1440 15506
rect 1504 15337 1532 18566
rect 1582 18320 1638 18329
rect 1582 18255 1638 18264
rect 1596 17338 1624 18255
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1582 16960 1638 16969
rect 1582 16895 1638 16904
rect 1596 16250 1624 16895
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1582 15600 1638 15609
rect 1582 15535 1638 15544
rect 1490 15328 1546 15337
rect 1490 15263 1546 15272
rect 1400 15088 1452 15094
rect 1400 15030 1452 15036
rect 1596 14618 1624 15535
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1596 13190 1624 14418
rect 1688 13326 1716 19654
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1780 14074 1808 17478
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1872 13814 1900 20402
rect 1964 18834 1992 22510
rect 2056 21078 2084 27520
rect 2044 21072 2096 21078
rect 2044 21014 2096 21020
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2044 19236 2096 19242
rect 2044 19178 2096 19184
rect 2056 19145 2084 19178
rect 2042 19136 2098 19145
rect 2042 19071 2098 19080
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1964 18426 1992 18770
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1780 13786 1900 13814
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1504 11558 1532 12242
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1320 5234 1348 9522
rect 1412 9024 1440 9862
rect 1504 9382 1532 11494
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1412 8996 1532 9024
rect 1504 6225 1532 8996
rect 1596 7546 1624 13126
rect 1688 12986 1716 13262
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1688 10810 1716 11086
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9654 1716 9862
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 9178 1716 9318
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 7750 1716 8366
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1688 7449 1716 7686
rect 1674 7440 1730 7449
rect 1674 7375 1730 7384
rect 1490 6216 1546 6225
rect 1490 6151 1546 6160
rect 1674 5808 1730 5817
rect 1674 5743 1676 5752
rect 1728 5743 1730 5752
rect 1676 5714 1728 5720
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1688 4758 1716 5714
rect 1676 4752 1728 4758
rect 1676 4694 1728 4700
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1688 2854 1716 3538
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1214 2680 1270 2689
rect 1214 2615 1270 2624
rect 848 2508 900 2514
rect 848 2450 900 2456
rect 478 82 534 480
rect 860 82 888 2450
rect 1688 1873 1716 2790
rect 1674 1864 1730 1873
rect 1674 1799 1730 1808
rect 478 54 888 82
rect 1398 82 1454 480
rect 1780 82 1808 13786
rect 1964 12442 1992 18022
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2332 16998 2360 17682
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2136 16448 2188 16454
rect 2136 16390 2188 16396
rect 2042 16144 2098 16153
rect 2042 16079 2098 16088
rect 2056 16046 2084 16079
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 2148 15162 2176 16390
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 2240 15366 2268 15914
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2148 14958 2176 15098
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 2056 13530 2084 13670
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1872 9450 1900 10950
rect 1964 10146 1992 12038
rect 2056 11286 2084 12038
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 2056 10606 2084 11222
rect 2148 11121 2176 14894
rect 2240 14226 2268 15302
rect 2332 14346 2360 16934
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 2240 14198 2360 14226
rect 2226 13968 2282 13977
rect 2226 13903 2282 13912
rect 2134 11112 2190 11121
rect 2134 11047 2190 11056
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 1964 10118 2084 10146
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1872 4060 1900 9386
rect 1964 9178 1992 9998
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1950 8936 2006 8945
rect 1950 8871 2006 8880
rect 1964 7002 1992 8871
rect 2056 7818 2084 10118
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2148 9654 2176 10066
rect 2240 9722 2268 13903
rect 2332 12986 2360 14198
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2424 12850 2452 19654
rect 2516 13326 2544 20198
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2596 19168 2648 19174
rect 2700 19156 2728 19858
rect 2648 19128 2728 19156
rect 2596 19110 2648 19116
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2608 15502 2636 16594
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 11898 2360 12242
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2608 11642 2636 15438
rect 2700 14618 2728 19128
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 2976 18358 3004 18770
rect 2964 18352 3016 18358
rect 2964 18294 3016 18300
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2976 17202 3004 18022
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2792 15473 2820 16934
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2884 15706 2912 15982
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2778 15464 2834 15473
rect 2778 15399 2834 15408
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2686 14512 2742 14521
rect 2686 14447 2688 14456
rect 2740 14447 2742 14456
rect 2688 14418 2740 14424
rect 2700 13938 2728 14418
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2700 13841 2728 13874
rect 2686 13832 2742 13841
rect 2686 13767 2742 13776
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2700 12986 2728 13398
rect 2792 13297 2820 14826
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2778 13288 2834 13297
rect 2778 13223 2834 13232
rect 2780 13184 2832 13190
rect 2884 13172 2912 13806
rect 2832 13144 2912 13172
rect 2780 13126 2832 13132
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2424 11354 2452 11630
rect 2608 11614 2820 11642
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2332 10713 2360 10950
rect 2424 10810 2452 11154
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2516 10742 2544 11018
rect 2504 10736 2556 10742
rect 2318 10704 2374 10713
rect 2504 10678 2556 10684
rect 2318 10639 2374 10648
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2332 10130 2360 10542
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2148 9178 2176 9590
rect 2332 9586 2360 10066
rect 2412 9920 2464 9926
rect 2464 9880 2544 9908
rect 2412 9862 2464 9868
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2332 8956 2360 9522
rect 2516 9518 2544 9880
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2412 8968 2464 8974
rect 2332 8928 2412 8956
rect 2412 8910 2464 8916
rect 2136 8288 2188 8294
rect 2136 8230 2188 8236
rect 2044 7812 2096 7818
rect 2044 7754 2096 7760
rect 2056 7342 2084 7754
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2056 5574 2084 6190
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 5370 2084 5510
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2056 4622 2084 5170
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 1952 4072 2004 4078
rect 1872 4049 1952 4060
rect 1858 4040 1952 4049
rect 1914 4032 1952 4040
rect 1952 4014 2004 4020
rect 1858 3975 1914 3984
rect 2148 3942 2176 8230
rect 2424 8090 2452 8910
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 6934 2268 7822
rect 2332 7478 2360 7958
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2228 6928 2280 6934
rect 2228 6870 2280 6876
rect 2240 4826 2268 6870
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2332 5778 2360 6598
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2320 5636 2372 5642
rect 2424 5624 2452 6598
rect 2372 5596 2452 5624
rect 2320 5578 2372 5584
rect 2332 5166 2360 5578
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2412 5092 2464 5098
rect 2412 5034 2464 5040
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2424 4690 2452 5034
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2240 3618 2268 4626
rect 2516 4486 2544 9454
rect 2608 7002 2636 11494
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2700 10130 2728 11154
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2700 8294 2728 8978
rect 2792 8537 2820 11614
rect 2884 10713 2912 12242
rect 2870 10704 2926 10713
rect 2870 10639 2926 10648
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2884 9722 2912 10134
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2778 8528 2834 8537
rect 2778 8463 2834 8472
rect 2778 8392 2834 8401
rect 2778 8327 2834 8336
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2596 6792 2648 6798
rect 2700 6769 2728 8230
rect 2596 6734 2648 6740
rect 2686 6760 2742 6769
rect 2608 6186 2636 6734
rect 2686 6695 2742 6704
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6458 2728 6598
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2608 5710 2636 6122
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2700 4554 2728 6394
rect 2792 5098 2820 8327
rect 2884 7206 2912 9658
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 2884 6798 2912 6870
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2884 5642 2912 6054
rect 2976 5914 3004 16934
rect 3068 15162 3096 27526
rect 3422 27520 3478 27526
rect 4802 27520 4858 28000
rect 5540 27532 5592 27538
rect 3882 21448 3938 21457
rect 3882 21383 3938 21392
rect 3516 20256 3568 20262
rect 3516 20198 3568 20204
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3436 19174 3464 19246
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3160 16017 3188 16594
rect 3146 16008 3202 16017
rect 3146 15943 3202 15952
rect 3160 15910 3188 15943
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3068 14958 3096 15098
rect 3160 14958 3188 15642
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3068 13433 3096 14894
rect 3054 13424 3110 13433
rect 3054 13359 3110 13368
rect 3252 13326 3280 19110
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3068 8906 3096 12786
rect 3344 12730 3372 17614
rect 3436 16046 3464 19110
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3528 15706 3556 20198
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3436 15162 3464 15506
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3436 14890 3464 15098
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3528 14618 3556 14894
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3436 14498 3464 14554
rect 3436 14470 3556 14498
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3252 12702 3372 12730
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3160 11257 3188 12174
rect 3146 11248 3202 11257
rect 3252 11234 3280 12702
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 11354 3372 12582
rect 3436 11898 3464 14010
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3436 11694 3464 11834
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3252 11206 3372 11234
rect 3146 11183 3202 11192
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3068 7410 3096 8298
rect 3160 8090 3188 9862
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 8498 3280 9318
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3252 8090 3280 8434
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3344 7886 3372 11206
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3238 7304 3294 7313
rect 3238 7239 3294 7248
rect 3146 7032 3202 7041
rect 3056 6996 3108 7002
rect 3146 6967 3202 6976
rect 3056 6938 3108 6944
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5302 3004 5510
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2976 5030 3004 5238
rect 3068 5166 3096 6938
rect 3160 6934 3188 6967
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3146 6760 3202 6769
rect 3146 6695 3202 6704
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2780 4616 2832 4622
rect 2884 4604 2912 4966
rect 2976 4826 3004 4966
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2832 4576 2912 4604
rect 2780 4558 2832 4564
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2148 3590 2268 3618
rect 2044 3392 2096 3398
rect 2148 3380 2176 3590
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2096 3352 2176 3380
rect 2044 3334 2096 3340
rect 2056 1329 2084 3334
rect 2240 2990 2268 3470
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 1737 2176 2246
rect 2134 1728 2190 1737
rect 2134 1663 2190 1672
rect 2042 1320 2098 1329
rect 2042 1255 2098 1264
rect 1398 54 1808 82
rect 2240 82 2268 2926
rect 2516 2854 2544 4422
rect 2700 3738 2728 4490
rect 2792 4214 2820 4558
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 3160 4154 3188 6695
rect 3252 4758 3280 7239
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 5914 3372 7142
rect 3436 7002 3464 11494
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3422 6216 3478 6225
rect 3422 6151 3478 6160
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3344 5574 3372 5714
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3344 4690 3372 5510
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3068 4126 3188 4154
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2884 3194 2912 3470
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2318 82 2374 480
rect 2240 54 2374 82
rect 3068 82 3096 4126
rect 3344 4010 3372 4626
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3344 3913 3372 3946
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3436 2990 3464 6151
rect 3528 4154 3556 14470
rect 3620 9500 3648 18566
rect 3712 12986 3740 18702
rect 3804 17105 3832 20198
rect 3790 17096 3846 17105
rect 3790 17031 3846 17040
rect 3896 14906 3924 21383
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4448 20534 4476 20946
rect 4620 20800 4672 20806
rect 4620 20742 4672 20748
rect 3976 20528 4028 20534
rect 3976 20470 4028 20476
rect 4436 20528 4488 20534
rect 4436 20470 4488 20476
rect 3804 14878 3924 14906
rect 3804 13977 3832 14878
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3790 13968 3846 13977
rect 3790 13903 3846 13912
rect 3896 13841 3924 14758
rect 3882 13832 3938 13841
rect 3882 13767 3938 13776
rect 3792 13728 3844 13734
rect 3988 13682 4016 20470
rect 4632 19922 4660 20742
rect 4620 19916 4672 19922
rect 4620 19858 4672 19864
rect 4712 19848 4764 19854
rect 4816 19825 4844 27520
rect 6182 27532 6238 28000
rect 6182 27520 6184 27532
rect 5540 27474 5592 27480
rect 6236 27520 6238 27532
rect 7654 27520 7710 28000
rect 9034 27520 9090 28000
rect 10414 27554 10470 28000
rect 11794 27554 11850 28000
rect 10414 27526 10916 27554
rect 10414 27520 10470 27526
rect 6184 27474 6236 27480
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 4896 20528 4948 20534
rect 4896 20470 4948 20476
rect 4712 19790 4764 19796
rect 4802 19816 4858 19825
rect 4724 19514 4752 19790
rect 4802 19751 4858 19760
rect 4712 19508 4764 19514
rect 4764 19468 4844 19496
rect 4712 19450 4764 19456
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4080 18630 4108 19246
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4264 18970 4292 19178
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4528 18692 4580 18698
rect 4528 18634 4580 18640
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4080 18222 4108 18566
rect 4436 18352 4488 18358
rect 4436 18294 4488 18300
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4080 17882 4108 18158
rect 4448 18086 4476 18294
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4080 14958 4108 15302
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4080 14482 4108 14894
rect 4172 14822 4200 17070
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4264 16726 4292 16934
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 4264 15910 4292 16662
rect 4356 16658 4384 17002
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4264 15638 4292 15846
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4080 14074 4108 14418
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3792 13670 3844 13676
rect 3804 13462 3832 13670
rect 3896 13654 4016 13682
rect 3792 13456 3844 13462
rect 3792 13398 3844 13404
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3804 12918 3832 13262
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3712 9625 3740 12718
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3698 9616 3754 9625
rect 3698 9551 3754 9560
rect 3620 9472 3740 9500
rect 3608 9376 3660 9382
rect 3606 9344 3608 9353
rect 3660 9344 3662 9353
rect 3606 9279 3662 9288
rect 3620 9178 3648 9279
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3620 5846 3648 8298
rect 3608 5840 3660 5846
rect 3608 5782 3660 5788
rect 3606 5672 3662 5681
rect 3606 5607 3608 5616
rect 3660 5607 3662 5616
rect 3608 5578 3660 5584
rect 3620 4826 3648 5578
rect 3712 5302 3740 9472
rect 3804 9178 3832 10066
rect 3896 9625 3924 13654
rect 4172 13530 4200 14554
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4356 13530 4384 13738
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 3988 13190 4016 13466
rect 4068 13320 4120 13326
rect 4448 13297 4476 18022
rect 4540 14906 4568 18634
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4724 17338 4752 17682
rect 4816 17626 4844 19468
rect 4908 18426 4936 20470
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4816 17598 4936 17626
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4816 17066 4844 17478
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4724 16726 4752 17002
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4632 15706 4660 16526
rect 4816 16250 4844 17002
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4632 15026 4660 15642
rect 4908 15162 4936 17598
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4908 15026 4936 15098
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 4540 14878 4752 14906
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4540 13394 4568 14418
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4068 13262 4120 13268
rect 4434 13288 4490 13297
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 4080 12850 4108 13262
rect 4434 13223 4490 13232
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4080 12442 4108 12786
rect 4356 12714 4384 13126
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3882 9616 3938 9625
rect 3882 9551 3938 9560
rect 3988 9489 4016 12378
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4080 11626 4108 12242
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4080 10470 4108 11018
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 10062 4108 10406
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4172 9674 4200 12106
rect 4264 11218 4292 12310
rect 4356 12238 4384 12650
rect 4448 12306 4476 13223
rect 4540 12374 4568 13330
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4540 11801 4568 12106
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4526 11792 4582 11801
rect 4526 11727 4582 11736
rect 4632 11694 4660 12038
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4356 11286 4384 11630
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4448 10538 4476 11154
rect 4540 11082 4568 11494
rect 4632 11218 4660 11630
rect 4724 11268 4752 14878
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4816 12986 4844 13466
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4908 12170 4936 13806
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4804 11280 4856 11286
rect 4724 11240 4804 11268
rect 4804 11222 4856 11228
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4540 10606 4568 11018
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4632 10266 4660 11154
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4724 10130 4752 10406
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4724 9722 4752 10066
rect 4908 9994 4936 10406
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4080 9646 4200 9674
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 3974 9480 4030 9489
rect 3974 9415 4030 9424
rect 3882 9344 3938 9353
rect 3882 9279 3938 9288
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7342 3832 7686
rect 3896 7342 3924 9279
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3988 7546 4016 9046
rect 4080 8634 4108 9646
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4172 7546 4200 9046
rect 4448 9042 4476 9318
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4448 8294 4476 8978
rect 4724 8974 4752 9658
rect 4908 9586 4936 9930
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4816 9178 4844 9454
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4264 8022 4292 8230
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 3976 7540 4028 7546
rect 4160 7540 4212 7546
rect 4028 7500 4108 7528
rect 3976 7482 4028 7488
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3804 6322 3832 7278
rect 3896 6984 3924 7278
rect 3896 6956 4016 6984
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3712 4826 3740 5102
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3804 4154 3832 6122
rect 3896 5778 3924 6802
rect 3988 6186 4016 6956
rect 4080 6254 4108 7500
rect 4160 7482 4212 7488
rect 4264 7002 4292 7958
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4356 7546 4384 7822
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4172 6905 4200 6938
rect 4158 6896 4214 6905
rect 4158 6831 4160 6840
rect 4212 6831 4214 6840
rect 4160 6802 4212 6808
rect 4172 6458 4200 6802
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3988 5234 4016 5646
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3528 4126 3648 4154
rect 3620 3194 3648 4126
rect 3712 4126 3832 4154
rect 3712 4078 3740 4126
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3712 3738 3740 4014
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3896 3505 3924 4762
rect 3988 4078 4016 5034
rect 4080 4865 4108 5510
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4080 4758 4108 4791
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3988 3670 4016 4014
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 4172 3602 4200 3946
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3882 3496 3938 3505
rect 3882 3431 3938 3440
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3620 2990 3648 3130
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 3252 2553 3280 2790
rect 3436 2650 3464 2926
rect 3620 2650 3648 2926
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3238 2544 3294 2553
rect 3238 2479 3294 2488
rect 4356 2446 4384 2994
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 3160 2009 3188 2382
rect 3146 2000 3202 2009
rect 3146 1935 3202 1944
rect 3330 82 3386 480
rect 3068 54 3386 82
rect 478 0 534 54
rect 1398 0 1454 54
rect 2318 0 2374 54
rect 3330 0 3386 54
rect 4250 82 4306 480
rect 4448 82 4476 8230
rect 4540 7206 4568 8366
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4908 6934 4936 7346
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4724 6390 4752 6802
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4802 6352 4858 6361
rect 4528 5296 4580 5302
rect 4528 5238 4580 5244
rect 4540 3670 4568 5238
rect 4724 5166 4752 6326
rect 4908 6322 4936 6666
rect 4802 6287 4858 6296
rect 4896 6316 4948 6322
rect 4816 5846 4844 6287
rect 4896 6258 4948 6264
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4724 4826 4752 5102
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4540 3126 4568 3606
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4540 2650 4568 3062
rect 4632 3058 4660 3674
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4724 2514 4752 4490
rect 4816 4146 4844 5782
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4908 3466 4936 5034
rect 5000 4622 5028 21422
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 5092 21010 5120 21286
rect 5276 21146 5304 23462
rect 5264 21140 5316 21146
rect 5264 21082 5316 21088
rect 5080 21004 5132 21010
rect 5080 20946 5132 20952
rect 5276 20398 5304 21082
rect 5552 20602 5580 27474
rect 6196 27443 6224 27474
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 7196 23656 7248 23662
rect 7196 23598 7248 23604
rect 7208 23361 7236 23598
rect 7194 23352 7250 23361
rect 7194 23287 7250 23296
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6196 21554 6224 22034
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 6288 21486 6316 22986
rect 7208 22778 7236 23122
rect 7288 22976 7340 22982
rect 7288 22918 7340 22924
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 6460 22500 6512 22506
rect 6460 22442 6512 22448
rect 6276 21480 6328 21486
rect 6276 21422 6328 21428
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 5092 18698 5120 20334
rect 5276 19922 5304 20334
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5460 19310 5488 19858
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5080 18692 5132 18698
rect 5080 18634 5132 18640
rect 5092 15706 5120 18634
rect 5276 18630 5304 19246
rect 5460 18834 5488 19246
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5184 18222 5212 18362
rect 5276 18222 5304 18566
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5184 17814 5212 18158
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 5092 14822 5120 15506
rect 5184 14958 5212 17750
rect 5368 17746 5396 18770
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5368 16522 5396 17002
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5276 15502 5304 15914
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5184 14482 5212 14894
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5184 11218 5212 14214
rect 5276 13977 5304 14758
rect 5262 13968 5318 13977
rect 5368 13938 5396 15846
rect 5460 13938 5488 18090
rect 5552 16114 5580 20538
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6012 17134 6040 20742
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 6104 18902 6132 20334
rect 6196 20262 6224 20946
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16250 6040 16662
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5552 15570 5580 15642
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 14482 5580 15506
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6104 14482 6132 18158
rect 6196 17270 6224 20198
rect 6288 19990 6316 20742
rect 6276 19984 6328 19990
rect 6276 19926 6328 19932
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6380 19378 6408 19790
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6380 17882 6408 19110
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6380 16998 6408 17818
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 16250 6224 16526
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5552 14278 5580 14418
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5998 14104 6054 14113
rect 5998 14039 6054 14048
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5262 13903 5318 13912
rect 5356 13932 5408 13938
rect 5276 13870 5304 13903
rect 5356 13874 5408 13880
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5446 13832 5502 13841
rect 5446 13767 5502 13776
rect 5460 12306 5488 13767
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5460 11898 5488 12242
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5552 11778 5580 13942
rect 6012 13841 6040 14039
rect 5998 13832 6054 13841
rect 6104 13802 6132 14418
rect 5998 13767 6054 13776
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6104 12986 6132 13738
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12238 5948 12582
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5460 11750 5580 11778
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5460 11150 5488 11750
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5460 10810 5488 11086
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 10130 5120 10610
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5092 9518 5120 10066
rect 5552 9586 5580 11630
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10062 6040 12650
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6104 11626 6132 12242
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5276 8838 5304 9522
rect 6104 9042 6132 10406
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 5356 8900 5408 8906
rect 5408 8860 5488 8888
rect 5356 8842 5408 8848
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 5092 5914 5120 6326
rect 5184 6186 5212 6598
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5184 5914 5212 6122
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5092 5302 5120 5850
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5184 5098 5212 5850
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5092 3942 5120 4694
rect 5276 4154 5304 8774
rect 5460 8430 5488 8860
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6104 8634 6132 8978
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5460 7886 5488 8366
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7410 5488 7686
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 6390 5396 7142
rect 5552 6866 5580 8434
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5552 6458 5580 6802
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 6012 6390 6040 6870
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 5234 5396 5510
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5552 4214 5580 6190
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6104 5166 6132 8570
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5644 4758 5672 5034
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5998 4312 6054 4321
rect 5998 4247 6054 4256
rect 5540 4208 5592 4214
rect 5276 4126 5396 4154
rect 5540 4150 5592 4156
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5000 3670 5028 3878
rect 5092 3738 5120 3878
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 5092 2922 5120 3674
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 4816 2514 4844 2858
rect 5184 2650 5212 3946
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4250 54 4476 82
rect 5262 82 5318 480
rect 5368 82 5396 4126
rect 5552 3126 5580 4150
rect 6012 4146 6040 4247
rect 6196 4154 6224 15574
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6380 15026 6408 15302
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6288 14074 6316 14418
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6380 13530 6408 14350
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6380 10810 6408 11154
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9722 6408 10066
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7002 6316 7822
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6288 5370 6316 5646
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6472 4826 6500 22442
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 6828 22160 6880 22166
rect 6828 22102 6880 22108
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6564 20262 6592 21082
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6564 19990 6592 20198
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6564 19174 6592 19926
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6564 17746 6592 18022
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6564 17202 6592 17682
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6564 14113 6592 17138
rect 6550 14104 6606 14113
rect 6550 14039 6606 14048
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6564 13530 6592 13942
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6564 12850 6592 13466
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 12714 6592 12786
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6564 12442 6592 12650
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6564 11354 6592 12378
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6564 9450 6592 10066
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6564 8634 6592 8978
rect 6656 8922 6684 21966
rect 6840 21350 6868 22102
rect 7012 21616 7064 21622
rect 7012 21558 7064 21564
rect 7024 21418 7052 21558
rect 6920 21412 6972 21418
rect 6920 21354 6972 21360
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6840 20058 6868 21286
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6748 17202 6776 18090
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6748 16250 6776 17138
rect 6840 16794 6868 17614
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6748 12170 6776 16050
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6840 14006 6868 14826
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6932 13814 6960 21354
rect 7012 20324 7064 20330
rect 7012 20266 7064 20272
rect 7024 19854 7052 20266
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7024 18426 7052 18770
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 7024 15638 7052 16934
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 7116 15162 7144 22374
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7208 21146 7236 21286
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7208 18358 7236 18770
rect 7300 18408 7328 22918
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7576 22030 7604 22578
rect 7380 22024 7432 22030
rect 7564 22024 7616 22030
rect 7432 21984 7512 22012
rect 7380 21966 7432 21972
rect 7380 21412 7432 21418
rect 7380 21354 7432 21360
rect 7392 21146 7420 21354
rect 7484 21146 7512 21984
rect 7564 21966 7616 21972
rect 7576 21554 7604 21966
rect 7668 21690 7696 27520
rect 9048 23474 9076 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 8956 23446 9076 23474
rect 8576 23248 8628 23254
rect 8576 23190 8628 23196
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 22710 7788 22918
rect 8588 22778 8616 23190
rect 8852 22976 8904 22982
rect 8852 22918 8904 22924
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8576 22772 8628 22778
rect 8576 22714 8628 22720
rect 7748 22704 7800 22710
rect 7800 22664 7880 22692
rect 7748 22646 7800 22652
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7668 20398 7696 20742
rect 7760 20602 7788 22442
rect 7852 21622 7880 22664
rect 8114 21720 8170 21729
rect 8114 21655 8170 21664
rect 7840 21616 7892 21622
rect 7840 21558 7892 21564
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7760 19310 7788 19654
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7654 19136 7710 19145
rect 7654 19071 7710 19080
rect 7300 18380 7420 18408
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 6932 13786 7052 13814
rect 7300 13802 7328 14214
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6840 12374 6868 12718
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6840 9500 6868 12174
rect 6932 10742 6960 12718
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 7024 9994 7052 13786
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7300 13530 7328 13738
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7102 13288 7158 13297
rect 7102 13223 7158 13232
rect 7116 11898 7144 13223
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7116 10112 7144 11834
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 10810 7236 11086
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7196 10124 7248 10130
rect 7116 10084 7196 10112
rect 7196 10066 7248 10072
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6920 9512 6972 9518
rect 6840 9472 6920 9500
rect 6920 9454 6972 9460
rect 6656 8894 6868 8922
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6656 7546 6684 7958
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7546 6776 7822
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6840 6798 6868 8894
rect 6932 8838 6960 9454
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 7698 6960 8774
rect 7024 8634 7052 9318
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7010 7712 7066 7721
rect 6932 7670 7010 7698
rect 7010 7647 7066 7656
rect 7024 7342 7052 7647
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6932 5914 6960 7142
rect 7300 7002 7328 7278
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7208 6458 7236 6734
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7300 6322 7328 6598
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 6932 5234 6960 5850
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7208 5030 7236 5850
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4826 7236 4966
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 6000 4140 6052 4146
rect 6196 4126 6408 4154
rect 6472 4146 6500 4762
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 6000 4082 6052 4088
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 6104 2854 6132 3538
rect 6092 2848 6144 2854
rect 6092 2790 6144 2796
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5262 54 5396 82
rect 6104 82 6132 2790
rect 6380 2582 6408 4126
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 7116 4010 7144 4694
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 6458 3904 6514 3913
rect 6458 3839 6514 3848
rect 6472 3466 6500 3839
rect 7024 3670 7052 3946
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6564 3194 6592 3402
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6748 3126 6776 3334
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 7024 2990 7052 3334
rect 7208 3194 7236 4762
rect 7392 4154 7420 18380
rect 7472 18148 7524 18154
rect 7472 18090 7524 18096
rect 7484 17882 7512 18090
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7576 16114 7604 16390
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7576 15638 7604 16050
rect 7564 15632 7616 15638
rect 7564 15574 7616 15580
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7484 13530 7512 13874
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7484 12918 7512 13466
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7576 10674 7604 15030
rect 7668 12889 7696 19071
rect 7760 18290 7788 19246
rect 7932 19168 7984 19174
rect 8024 19168 8076 19174
rect 7984 19128 8024 19156
rect 7932 19110 7984 19116
rect 8024 19110 8076 19116
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7944 17338 7972 17750
rect 8036 17338 8064 18702
rect 8128 18290 8156 21655
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8128 17814 8156 18226
rect 8116 17808 8168 17814
rect 8116 17750 8168 17756
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7944 16794 7972 17274
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7840 16720 7892 16726
rect 7840 16662 7892 16668
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7760 15348 7788 16526
rect 7852 16250 7880 16662
rect 8128 16522 8156 17750
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7852 15978 7880 16186
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7852 15706 7880 15914
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 7840 15360 7892 15366
rect 7760 15320 7840 15348
rect 7840 15302 7892 15308
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14550 7788 14758
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7852 14006 7880 15302
rect 8036 15162 8064 15438
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7760 13190 7788 13670
rect 7944 13190 7972 14350
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7654 12880 7710 12889
rect 7654 12815 7710 12824
rect 7760 11830 7788 13126
rect 8036 12306 8064 14894
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8128 14074 8156 14486
rect 8220 14346 8248 22714
rect 8588 22137 8616 22714
rect 8864 22234 8892 22918
rect 8852 22228 8904 22234
rect 8852 22170 8904 22176
rect 8574 22128 8630 22137
rect 8574 22063 8630 22072
rect 8668 21956 8720 21962
rect 8668 21898 8720 21904
rect 8680 21554 8708 21898
rect 8864 21554 8892 22170
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8576 21344 8628 21350
rect 8576 21286 8628 21292
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8496 20602 8524 20946
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8588 19446 8616 21286
rect 8956 20534 8984 23446
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 9232 22710 9260 23054
rect 9220 22704 9272 22710
rect 9220 22646 9272 22652
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 9048 21418 9076 22374
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9036 21412 9088 21418
rect 9036 21354 9088 21360
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 8944 20528 8996 20534
rect 8942 20496 8944 20505
rect 8996 20496 8998 20505
rect 9048 20466 9076 20742
rect 9140 20466 9168 21490
rect 9232 21146 9260 22646
rect 9588 22636 9640 22642
rect 9588 22578 9640 22584
rect 9312 22500 9364 22506
rect 9312 22442 9364 22448
rect 9324 21894 9352 22442
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9508 21146 9536 21966
rect 9600 21962 9628 22578
rect 9588 21956 9640 21962
rect 9588 21898 9640 21904
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9494 21040 9550 21049
rect 9494 20975 9550 20984
rect 9508 20942 9536 20975
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9692 20602 9720 20878
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 8942 20431 8998 20440
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9048 20058 9076 20402
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 9140 20058 9168 20266
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9588 19984 9640 19990
rect 9588 19926 9640 19932
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8956 19242 8984 19858
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 8956 19145 8984 19178
rect 8942 19136 8998 19145
rect 8942 19071 8998 19080
rect 9416 18970 9444 19246
rect 9600 19174 9628 19926
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18086 8340 18566
rect 8680 18086 8708 18702
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 9048 18426 9076 18634
rect 9600 18630 9628 19110
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9048 18222 9076 18362
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8312 17610 8340 18022
rect 8680 17785 8708 18022
rect 8666 17776 8722 17785
rect 8666 17711 8722 17720
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 8312 16522 8340 17546
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8312 14414 8340 16458
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8496 15570 8524 15914
rect 8588 15570 8616 17002
rect 8680 16794 8708 17614
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8680 16590 8708 16730
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8680 16114 8708 16526
rect 9048 16454 9076 18158
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8588 14822 8616 15506
rect 8680 15026 8708 16050
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8588 13814 8616 14758
rect 8680 14618 8708 14826
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8772 14550 8800 14826
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8588 13786 8708 13814
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8128 12646 8156 13262
rect 8220 12986 8248 13398
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12986 8340 13126
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 8036 11626 8064 12038
rect 8312 11898 8340 12242
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7668 10810 7696 11290
rect 7760 11286 7788 11562
rect 8036 11354 8064 11562
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 8036 10538 8064 11290
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8036 10266 8064 10474
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8404 10130 8432 11154
rect 8496 10742 8524 12582
rect 8588 12306 8616 13194
rect 8680 12764 8708 13786
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8772 12918 8800 13126
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8680 12736 8800 12764
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 11558 8616 12242
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8574 11112 8630 11121
rect 8574 11047 8630 11056
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8036 9722 8064 10066
rect 8404 9722 8432 10066
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 7838 9616 7894 9625
rect 7838 9551 7894 9560
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 9042 7512 9454
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7484 8838 7512 8978
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 8022 7512 8230
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7484 6390 7512 7958
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7668 6458 7696 6870
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7484 5914 7512 6326
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7300 4126 7420 4154
rect 7300 3534 7328 4126
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7392 3194 7420 3606
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7208 2854 7236 3130
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 6932 2530 6960 2586
rect 7196 2576 7248 2582
rect 6932 2524 7196 2530
rect 6932 2518 7248 2524
rect 6932 2502 7236 2518
rect 6182 82 6238 480
rect 6104 54 6238 82
rect 4250 0 4306 54
rect 5262 0 5318 54
rect 6182 0 6238 54
rect 7194 82 7250 480
rect 7484 82 7512 5238
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4758 7788 4966
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7760 4282 7788 4694
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7852 4146 7880 9551
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7944 8294 7972 9114
rect 8392 8832 8444 8838
rect 8444 8792 8524 8820
rect 8392 8774 8444 8780
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 8022 7972 8230
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 8220 7886 8248 8502
rect 8390 7984 8446 7993
rect 8496 7954 8524 8792
rect 8390 7919 8446 7928
rect 8484 7948 8536 7954
rect 8404 7886 8432 7919
rect 8484 7890 8536 7896
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8036 6730 8064 7754
rect 8404 7478 8432 7822
rect 8392 7472 8444 7478
rect 8298 7440 8354 7449
rect 8392 7414 8444 7420
rect 8298 7375 8354 7384
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 8036 6186 8064 6666
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5914 7972 6054
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8036 5030 8064 6122
rect 8220 5914 8248 6258
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 8036 4622 8064 4966
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7668 2582 7696 3946
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8036 2650 8064 2994
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 8128 626 8156 4014
rect 8220 3670 8248 5850
rect 8312 3942 8340 7375
rect 8496 6730 8524 7890
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8588 6458 8616 11047
rect 8680 10198 8708 11154
rect 8772 10588 8800 12736
rect 8850 12472 8906 12481
rect 8850 12407 8906 12416
rect 8864 10713 8892 12407
rect 8850 10704 8906 10713
rect 8850 10639 8906 10648
rect 8772 10560 8892 10588
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8772 8838 8800 9386
rect 8864 9081 8892 10560
rect 8850 9072 8906 9081
rect 8850 9007 8906 9016
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8634 8800 8774
rect 8864 8634 8892 8910
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8680 5030 8708 5646
rect 8864 5166 8892 6938
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8864 4826 8892 5102
rect 8956 4826 8984 14214
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 9048 10849 9076 13942
rect 9140 12850 9168 17070
rect 9232 16726 9260 18566
rect 9600 17048 9628 18566
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9692 17542 9720 18158
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9680 17060 9732 17066
rect 9600 17020 9680 17048
rect 9680 17002 9732 17008
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16794 9536 16934
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9232 15706 9260 16662
rect 9508 16250 9536 16730
rect 9692 16250 9720 17002
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9692 15910 9720 16186
rect 9784 16114 9812 24006
rect 10704 23866 10732 24210
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 10692 23520 10744 23526
rect 10692 23462 10744 23468
rect 9864 23248 9916 23254
rect 9864 23190 9916 23196
rect 9876 22778 9904 23190
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9876 21078 9904 22714
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9876 20058 9904 21014
rect 9968 20602 9996 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 10060 22642 10088 23054
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10152 21350 10180 22102
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10152 20806 10180 21286
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 10152 20262 10180 20742
rect 10612 20466 10640 20810
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 10152 19514 10180 20198
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10612 19514 10640 19790
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10152 18884 10180 19314
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10232 18896 10284 18902
rect 10152 18856 10232 18884
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9876 15162 9904 15370
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9232 13734 9260 13806
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9232 12209 9260 13670
rect 9416 13394 9444 14350
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 13734 9536 14214
rect 9692 13920 9720 15030
rect 9876 14482 9904 15098
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9876 14074 9904 14418
rect 9968 14074 9996 18090
rect 10152 17882 10180 18856
rect 10232 18838 10284 18844
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10704 17678 10732 23462
rect 10888 22574 10916 27526
rect 11532 27526 11850 27554
rect 11532 24274 11560 27526
rect 11794 27520 11850 27526
rect 13174 27520 13230 28000
rect 14646 27520 14702 28000
rect 16026 27520 16082 28000
rect 17406 27520 17462 28000
rect 18786 27520 18842 28000
rect 20166 27520 20222 28000
rect 21638 27520 21694 28000
rect 23018 27554 23074 28000
rect 24398 27554 24454 28000
rect 22664 27526 23074 27554
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11244 23656 11296 23662
rect 11164 23616 11244 23644
rect 11164 23322 11192 23616
rect 11244 23598 11296 23604
rect 11348 23474 11376 24006
rect 11532 23662 11560 24210
rect 11520 23656 11572 23662
rect 11520 23598 11572 23604
rect 11716 23526 11744 24210
rect 12992 23588 13044 23594
rect 12992 23530 13044 23536
rect 11256 23446 11376 23474
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10796 22030 10824 22374
rect 11072 22234 11100 22918
rect 11060 22228 11112 22234
rect 11060 22170 11112 22176
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 11072 21554 11100 22170
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10796 20058 10824 20878
rect 11164 20602 11192 21014
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10888 18902 10916 20402
rect 11256 19258 11284 23446
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 11348 22710 11376 23122
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 11532 22098 11560 22714
rect 12176 22574 12204 23122
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11532 21690 11560 22034
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 12084 20602 12112 20946
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11336 19440 11388 19446
rect 11336 19382 11388 19388
rect 11072 19230 11284 19258
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10152 15570 10180 17478
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16794 10732 17614
rect 10796 17066 10824 17750
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10796 16250 10824 17002
rect 10888 16590 10916 17002
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 10152 15094 10180 15506
rect 10690 15464 10746 15473
rect 10690 15399 10746 15408
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9692 13892 9812 13920
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9600 12646 9628 13398
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9692 12646 9720 13262
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9218 12200 9274 12209
rect 9218 12135 9274 12144
rect 9416 11558 9444 12582
rect 9692 12374 9720 12582
rect 9680 12368 9732 12374
rect 9586 12336 9642 12345
rect 9680 12310 9732 12316
rect 9586 12271 9642 12280
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9034 10840 9090 10849
rect 9416 10810 9444 11494
rect 9034 10775 9090 10784
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9048 10062 9076 10610
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9324 10198 9352 10542
rect 9416 10538 9444 10746
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9048 8634 9076 8842
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9048 8294 9076 8570
rect 9126 8528 9182 8537
rect 9126 8463 9182 8472
rect 9036 8288 9088 8294
rect 9140 8276 9168 8463
rect 9232 8430 9260 8910
rect 9324 8566 9352 9386
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9416 8362 9444 8842
rect 9508 8838 9536 9522
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9140 8248 9260 8276
rect 9036 8230 9088 8236
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9048 4758 9076 5714
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 8850 4040 8906 4049
rect 8850 3975 8906 3984
rect 8944 4004 8996 4010
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8312 3058 8340 3878
rect 8864 3738 8892 3975
rect 8944 3946 8996 3952
rect 8956 3777 8984 3946
rect 8942 3768 8998 3777
rect 8852 3732 8904 3738
rect 8942 3703 8998 3712
rect 8852 3674 8904 3680
rect 8956 3097 8984 3703
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 8942 3088 8998 3097
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8852 3052 8904 3058
rect 8942 3023 8998 3032
rect 8852 2994 8904 3000
rect 8758 2544 8814 2553
rect 8758 2479 8814 2488
rect 8772 2310 8800 2479
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8128 598 8248 626
rect 7194 54 7512 82
rect 8114 82 8170 480
rect 8220 82 8248 598
rect 8114 54 8248 82
rect 8864 82 8892 2994
rect 9140 2990 9168 3402
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9232 2922 9260 8248
rect 9416 7818 9444 8298
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9508 7478 9536 8774
rect 9600 7546 9628 12271
rect 9784 11642 9812 13892
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9876 13530 9904 13738
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9876 12442 9904 13330
rect 9968 13326 9996 13670
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9968 12714 9996 13262
rect 10060 13258 10088 14418
rect 10152 14006 10180 15030
rect 10704 15026 10732 15399
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 14962
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10152 13326 10180 13738
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9968 12442 9996 12650
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9876 11762 9904 12378
rect 10704 11830 10732 13738
rect 10796 12238 10824 16050
rect 10888 15570 10916 16390
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10980 15162 11008 16934
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10980 12918 11008 14282
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 11898 10824 12174
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9784 11614 9996 11642
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9692 7410 9720 7822
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9600 6934 9628 7210
rect 9692 7002 9720 7346
rect 9876 7002 9904 10950
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9876 6866 9904 6938
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 6390 9904 6802
rect 9968 6798 9996 11614
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10520 10810 10548 11154
rect 10704 11082 10732 11766
rect 10888 11558 10916 12310
rect 10980 12238 11008 12650
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11286 10916 11494
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10520 10606 10548 10746
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 10198 10180 10406
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10198 10732 11018
rect 10888 10810 10916 11222
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10980 10742 11008 12174
rect 11072 11150 11100 19230
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10152 9722 10180 10134
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10152 9382 10180 9658
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10244 9489 10272 9522
rect 10230 9480 10286 9489
rect 10230 9415 10286 9424
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9178 10732 9930
rect 10980 9654 11008 10678
rect 11072 10266 11100 11086
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10060 8276 10088 9046
rect 10140 8288 10192 8294
rect 10060 8248 10140 8276
rect 10060 7750 10088 8248
rect 10140 8230 10192 8236
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 7274 10088 7686
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10152 7206 10180 7958
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10140 7200 10192 7206
rect 10060 7148 10140 7154
rect 10060 7142 10192 7148
rect 10060 7126 10180 7142
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9310 4856 9366 4865
rect 9310 4791 9366 4800
rect 9324 4486 9352 4791
rect 9312 4480 9364 4486
rect 9416 4457 9444 6326
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9508 5302 9536 6190
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5846 9996 6054
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9692 5370 9720 5578
rect 9968 5370 9996 5782
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9692 4604 9720 5306
rect 9862 4856 9918 4865
rect 9862 4791 9918 4800
rect 9876 4690 9904 4791
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9772 4616 9824 4622
rect 9600 4576 9772 4604
rect 9312 4422 9364 4428
rect 9402 4448 9458 4457
rect 9324 4357 9352 4422
rect 9402 4383 9458 4392
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9324 3534 9352 4014
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9416 3058 9444 4383
rect 9600 4282 9628 4576
rect 9772 4558 9824 4564
rect 9588 4276 9640 4282
rect 9508 4236 9588 4264
rect 9508 4010 9536 4236
rect 9640 4236 9720 4264
rect 9588 4218 9640 4224
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9508 3913 9536 3946
rect 9494 3904 9550 3913
rect 9494 3839 9550 3848
rect 9692 3738 9720 4236
rect 9876 4214 9904 4626
rect 9968 4321 9996 5306
rect 9954 4312 10010 4321
rect 9954 4247 10010 4256
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9876 3398 9904 4150
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9588 2508 9640 2514
rect 9680 2508 9732 2514
rect 9640 2468 9680 2496
rect 9588 2450 9640 2456
rect 9680 2450 9732 2456
rect 9784 2378 9812 3062
rect 9876 2854 9904 3334
rect 9968 3194 9996 4247
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9772 2372 9824 2378
rect 10060 2360 10088 7126
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10152 6458 10180 6802
rect 10322 6760 10378 6769
rect 10322 6695 10378 6704
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10336 6322 10364 6695
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10336 6225 10364 6258
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 11072 5846 11100 7278
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10876 5704 10928 5710
rect 10506 5672 10562 5681
rect 10876 5646 10928 5652
rect 10506 5607 10562 5616
rect 10520 5574 10548 5607
rect 10508 5568 10560 5574
rect 10692 5568 10744 5574
rect 10508 5510 10560 5516
rect 10612 5528 10692 5556
rect 10520 5370 10548 5510
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10612 5166 10640 5528
rect 10692 5510 10744 5516
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10152 4282 10180 5102
rect 10704 5098 10732 5306
rect 10888 5234 10916 5646
rect 11164 5370 11192 19110
rect 11348 18222 11376 19382
rect 11900 19174 11928 19858
rect 12084 19786 12112 20538
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18834 11928 19110
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 11808 18086 11836 18770
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11256 16454 11284 17138
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11256 15162 11284 16390
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11244 14476 11296 14482
rect 11348 14464 11376 18022
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 11440 16182 11468 16662
rect 11716 16590 11744 17546
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11624 15910 11652 16526
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11440 15094 11468 15506
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11296 14436 11376 14464
rect 11244 14418 11296 14424
rect 11256 13802 11284 14418
rect 11440 13870 11468 15030
rect 11532 15026 11560 15642
rect 11624 15638 11652 15846
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11808 14521 11836 18022
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11992 16998 12020 17682
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 15570 11928 16390
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11900 14958 11928 15506
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11794 14512 11850 14521
rect 11704 14476 11756 14482
rect 11794 14447 11850 14456
rect 11704 14418 11756 14424
rect 11716 14006 11744 14418
rect 12176 14414 12204 18566
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11704 14000 11756 14006
rect 11610 13968 11666 13977
rect 11704 13942 11756 13948
rect 11610 13903 11666 13912
rect 11888 13932 11940 13938
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11256 13297 11284 13738
rect 11624 13530 11652 13903
rect 11888 13874 11940 13880
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11242 13288 11298 13297
rect 11242 13223 11298 13232
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11348 8294 11376 8910
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11256 6662 11284 7822
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11256 6322 11284 6598
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4826 10732 5034
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10152 3738 10180 4082
rect 10612 3924 10640 4218
rect 10796 3942 10824 4422
rect 10784 3936 10836 3942
rect 10612 3896 10732 3924
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3754 10732 3896
rect 10784 3878 10836 3884
rect 10140 3732 10192 3738
rect 10658 3726 10732 3754
rect 10658 3720 10686 3726
rect 10140 3674 10192 3680
rect 10612 3692 10686 3720
rect 10612 3602 10640 3692
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10796 3516 10824 3878
rect 10704 3488 10824 3516
rect 10232 3460 10284 3466
rect 10232 3402 10284 3408
rect 10244 2990 10272 3402
rect 10704 3398 10732 3488
rect 10980 3398 11008 4694
rect 11072 4486 11100 5238
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10428 3126 10456 3334
rect 10888 3210 10916 3334
rect 11072 3210 11100 4422
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 10888 3182 11100 3210
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10888 2990 10916 3182
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10888 2689 10916 2926
rect 10874 2680 10930 2689
rect 10874 2615 10930 2624
rect 11164 2582 11192 4014
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 10232 2372 10284 2378
rect 10060 2332 10232 2360
rect 9772 2314 9824 2320
rect 10232 2314 10284 2320
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9126 82 9182 480
rect 9968 105 9996 2246
rect 8864 54 9182 82
rect 7194 0 7250 54
rect 8114 0 8170 54
rect 9126 0 9182 54
rect 9954 96 10010 105
rect 9954 31 10010 40
rect 10046 82 10102 480
rect 10244 82 10272 2314
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 10704 1601 10732 2246
rect 10690 1592 10746 1601
rect 10690 1527 10746 1536
rect 10046 54 10272 82
rect 11058 82 11114 480
rect 11256 82 11284 6122
rect 11348 4826 11376 8230
rect 11624 7478 11652 11698
rect 11716 10810 11744 13806
rect 11794 12744 11850 12753
rect 11794 12679 11850 12688
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11808 8566 11836 12679
rect 11900 11762 11928 13874
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12084 12646 12112 13330
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11992 11121 12020 12582
rect 11978 11112 12034 11121
rect 11978 11047 12034 11056
rect 11978 10568 12034 10577
rect 11978 10503 12034 10512
rect 11992 10130 12020 10503
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11992 9761 12020 10066
rect 11978 9752 12034 9761
rect 11978 9687 12034 9696
rect 11992 9654 12020 9687
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 12084 8401 12112 12582
rect 12176 12374 12204 13670
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12176 11626 12204 12310
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12176 10810 12204 11154
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12268 8498 12296 23462
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12452 21457 12480 22510
rect 12544 22234 12572 22918
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 12438 21448 12494 21457
rect 12438 21383 12494 21392
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12544 20602 12572 20946
rect 12532 20596 12584 20602
rect 12452 20556 12532 20584
rect 12452 19446 12480 20556
rect 12532 20538 12584 20544
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12452 18970 12480 19382
rect 12544 19310 12572 19654
rect 12532 19304 12584 19310
rect 12636 19281 12664 22374
rect 12532 19246 12584 19252
rect 12622 19272 12678 19281
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12452 18358 12480 18906
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12452 17746 12480 18294
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12452 17338 12480 17682
rect 12544 17678 12572 19246
rect 12622 19207 12678 19216
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12360 13308 12388 15438
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 14550 12664 15302
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12530 14104 12586 14113
rect 12530 14039 12586 14048
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12452 13530 12480 13874
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 13320 12492 13326
rect 12360 13280 12440 13308
rect 12440 13262 12492 13268
rect 12452 12442 12480 13262
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12544 12322 12572 14039
rect 12452 12294 12572 12322
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12360 10742 12388 11766
rect 12452 11014 12480 12294
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10810 12480 10950
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12544 10538 12572 11018
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12070 8392 12126 8401
rect 12070 8327 12126 8336
rect 12360 8294 12388 9114
rect 12544 8537 12572 10474
rect 12636 10266 12664 10474
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12530 8528 12586 8537
rect 12530 8463 12586 8472
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12452 7954 12480 8366
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12544 8022 12572 8230
rect 12636 8090 12664 10202
rect 12728 9568 12756 23462
rect 13004 23050 13032 23530
rect 13188 23322 13216 27520
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 14384 23322 14412 23598
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14660 23254 14688 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 16040 23866 16068 27520
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16028 23860 16080 23866
rect 16028 23802 16080 23808
rect 16960 23594 16988 24210
rect 17420 23866 17448 27520
rect 18328 24880 18380 24886
rect 18328 24822 18380 24828
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 18064 23866 18092 24210
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 18052 23860 18104 23866
rect 18052 23802 18104 23808
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18234 23624 18290 23633
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 16948 23588 17000 23594
rect 16948 23530 17000 23536
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 12992 23044 13044 23050
rect 12912 23004 12992 23032
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12820 21418 12848 21830
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12820 19310 12848 19790
rect 12912 19334 12940 23004
rect 12992 22986 13044 22992
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 12808 19304 12860 19310
rect 12912 19306 13032 19334
rect 12808 19246 12860 19252
rect 12820 18290 12848 19246
rect 13004 19122 13032 19306
rect 12912 19094 13032 19122
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 13190 12848 16934
rect 12912 14958 12940 19094
rect 13096 18873 13124 22714
rect 13452 22704 13504 22710
rect 13452 22646 13504 22652
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 13268 22160 13320 22166
rect 13268 22102 13320 22108
rect 13280 21690 13308 22102
rect 13268 21684 13320 21690
rect 13268 21626 13320 21632
rect 13280 21146 13308 21626
rect 13372 21622 13400 22374
rect 13464 22234 13492 22646
rect 13832 22642 13860 23122
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13728 22500 13780 22506
rect 13648 22460 13728 22488
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13360 21616 13412 21622
rect 13360 21558 13412 21564
rect 13544 21616 13596 21622
rect 13544 21558 13596 21564
rect 13556 21418 13584 21558
rect 13544 21412 13596 21418
rect 13544 21354 13596 21360
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13280 20466 13308 20878
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13188 20058 13216 20198
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13188 19242 13216 19994
rect 13358 19816 13414 19825
rect 13358 19751 13414 19760
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 13176 19236 13228 19242
rect 13176 19178 13228 19184
rect 13188 18970 13216 19178
rect 13280 19174 13308 19246
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13176 18964 13228 18970
rect 13228 18924 13308 18952
rect 13176 18906 13228 18912
rect 13082 18864 13138 18873
rect 13082 18799 13138 18808
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18154 13216 18702
rect 13280 18426 13308 18924
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13188 17882 13216 18090
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13280 17134 13308 17274
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 13004 15162 13032 15914
rect 13096 15638 13124 15982
rect 13188 15706 13216 16526
rect 13280 16454 13308 17070
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13280 15706 13308 15914
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 13004 14634 13032 15098
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 12912 14606 13032 14634
rect 12912 13814 12940 14606
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13004 14074 13032 14486
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12912 13786 13032 13814
rect 13004 13734 13032 13786
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13004 13530 13032 13670
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 11694 12848 13126
rect 13004 12986 13032 13466
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12912 12345 12940 12582
rect 12898 12336 12954 12345
rect 12898 12271 12954 12280
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12820 11354 12848 11630
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12728 9540 12848 9568
rect 12624 8084 12676 8090
rect 12676 8044 12756 8072
rect 12624 8026 12676 8032
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12544 7750 12572 7958
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 12544 7206 12572 7686
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6798 12664 7142
rect 12728 6934 12756 8044
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11440 4758 11468 6666
rect 11532 6458 11560 6734
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 12636 5778 12664 6734
rect 12728 6458 12756 6870
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12360 5681 12388 5714
rect 12346 5672 12402 5681
rect 12346 5607 12402 5616
rect 12360 5370 12388 5607
rect 12544 5370 12572 5714
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12820 5302 12848 9540
rect 12912 7732 12940 12038
rect 13004 8634 13032 12786
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13096 11354 13124 12174
rect 13188 12102 13216 14758
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13096 11257 13124 11290
rect 13082 11248 13138 11257
rect 13280 11218 13308 11562
rect 13082 11183 13138 11192
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13280 10266 13308 11154
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13188 9722 13216 10134
rect 13176 9716 13228 9722
rect 13228 9676 13308 9704
rect 13176 9658 13228 9664
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13096 9178 13124 9386
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13188 8906 13216 9386
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13280 8634 13308 9676
rect 13372 9042 13400 19751
rect 13556 18970 13584 21354
rect 13648 21060 13676 22460
rect 13728 22442 13780 22448
rect 13728 21956 13780 21962
rect 13728 21898 13780 21904
rect 13740 21554 13768 21898
rect 13832 21729 13860 22578
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 13818 21720 13874 21729
rect 13818 21655 13874 21664
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13728 21072 13780 21078
rect 13648 21032 13728 21060
rect 13728 21014 13780 21020
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 13740 20058 13768 21014
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13832 19922 13860 21014
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 17066 13584 18022
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 13740 15978 13768 16662
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13832 15026 13860 19314
rect 13924 19310 13952 21082
rect 14016 21049 14044 22510
rect 15304 22234 15332 23530
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 18052 23180 18104 23186
rect 18052 23122 18104 23128
rect 15396 22506 15424 23122
rect 15936 22976 15988 22982
rect 15936 22918 15988 22924
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15292 22228 15344 22234
rect 15344 22188 15516 22216
rect 15292 22170 15344 22176
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 14002 21040 14058 21049
rect 14002 20975 14058 20984
rect 14200 20602 14228 21286
rect 14384 21078 14412 21490
rect 14556 21344 14608 21350
rect 14476 21304 14556 21332
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14476 20262 14504 21304
rect 14556 21286 14608 21292
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14646 20496 14702 20505
rect 14646 20431 14702 20440
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14476 19922 14504 20198
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13924 18426 13952 19246
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14108 18222 14136 18566
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14002 17776 14058 17785
rect 14108 17746 14136 18158
rect 14002 17711 14058 17720
rect 14096 17740 14148 17746
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13924 17338 13952 17614
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14618 13860 14962
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 14016 14498 14044 17711
rect 14096 17682 14148 17688
rect 14108 16794 14136 17682
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17202 14412 17478
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14200 16726 14228 16934
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14108 15978 14136 16390
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14550 14136 14962
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 14200 14618 14228 14826
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 13924 14470 14044 14498
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 13924 13814 13952 14470
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 14016 14074 14044 14350
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13924 13786 14044 13814
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12850 13676 13126
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13740 12714 13768 12922
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13740 12442 13768 12650
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13556 10062 13584 10610
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13464 9382 13492 9998
rect 13556 9586 13584 9998
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13542 9072 13598 9081
rect 13360 9036 13412 9042
rect 13542 9007 13598 9016
rect 13360 8978 13412 8984
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12992 7744 13044 7750
rect 12912 7704 12992 7732
rect 12992 7686 13044 7692
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11532 4214 11560 5034
rect 11610 4856 11666 4865
rect 11610 4791 11666 4800
rect 11624 4690 11652 4791
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 11624 4282 11652 4626
rect 11886 4448 11942 4457
rect 11886 4383 11942 4392
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11624 3505 11652 4218
rect 11796 3528 11848 3534
rect 11610 3496 11666 3505
rect 11796 3470 11848 3476
rect 11610 3431 11666 3440
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11532 2514 11560 3334
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11716 2582 11744 2926
rect 11808 2854 11836 3470
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11440 2310 11468 2450
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 11808 1465 11836 2790
rect 11900 2650 11928 4383
rect 12176 4282 12204 4626
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12268 4154 12296 4422
rect 12176 4126 12296 4154
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12176 2446 12204 4126
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 3194 12296 3538
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12636 2582 12664 2790
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12636 2378 12664 2518
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 12728 2009 12756 2382
rect 12714 2000 12770 2009
rect 12714 1935 12770 1944
rect 11794 1456 11850 1465
rect 11794 1391 11850 1400
rect 11058 54 11284 82
rect 11978 128 12034 480
rect 11978 76 11980 128
rect 12032 76 12034 128
rect 10046 0 10102 54
rect 11058 0 11114 54
rect 11978 0 12034 76
rect 12912 82 12940 7278
rect 13004 6186 13032 7686
rect 13096 6236 13124 8502
rect 13280 8022 13308 8570
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13188 7392 13216 7754
rect 13280 7546 13308 7958
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13268 7404 13320 7410
rect 13188 7364 13268 7392
rect 13268 7346 13320 7352
rect 13280 6934 13308 7346
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13176 6248 13228 6254
rect 13096 6208 13176 6236
rect 13176 6190 13228 6196
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13096 5914 13124 6054
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13188 5817 13216 6190
rect 13174 5808 13230 5817
rect 13174 5743 13230 5752
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 2961 13032 3878
rect 12990 2952 13046 2961
rect 12990 2887 13046 2896
rect 13280 1737 13308 4422
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13372 2990 13400 3334
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13464 2378 13492 4966
rect 13556 3505 13584 9007
rect 13648 7478 13676 10950
rect 13740 8401 13768 12106
rect 13924 11558 13952 12582
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13820 10736 13872 10742
rect 13910 10704 13966 10713
rect 13872 10684 13910 10690
rect 13820 10678 13910 10684
rect 13832 10662 13910 10678
rect 13910 10639 13966 10648
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13726 8392 13782 8401
rect 13726 8327 13782 8336
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13636 7472 13688 7478
rect 13740 7449 13768 8230
rect 13636 7414 13688 7420
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13740 7274 13768 7375
rect 13832 7274 13860 8842
rect 13924 8566 13952 8978
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 14016 8362 14044 13786
rect 14108 12850 14136 14486
rect 14200 14074 14228 14554
rect 14278 14512 14334 14521
rect 14278 14447 14334 14456
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14200 13530 14228 14010
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14108 12238 14136 12786
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11762 14228 12038
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14200 11286 14228 11494
rect 14188 11280 14240 11286
rect 14188 11222 14240 11228
rect 14200 10470 14228 11222
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 7002 13860 7210
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6322 13860 6598
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 14016 5914 14044 8298
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13832 4826 13860 5782
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13648 3942 13676 4694
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13542 3496 13598 3505
rect 13542 3431 13598 3440
rect 13648 2650 13676 3878
rect 13832 3670 13860 4762
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13832 3194 13860 3606
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 13266 1728 13322 1737
rect 13266 1663 13322 1672
rect 12990 82 13046 480
rect 12912 54 13046 82
rect 12990 0 13046 54
rect 13910 82 13966 480
rect 14108 82 14136 8434
rect 14200 8294 14228 10406
rect 14292 8956 14320 14447
rect 14568 13814 14596 20334
rect 14660 13841 14688 20431
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14752 18630 14780 19246
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 18290 14780 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 15304 17814 15332 18702
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15304 16726 15332 16934
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16114 15332 16390
rect 15396 16114 15424 20198
rect 15488 18986 15516 22188
rect 15672 21078 15700 22374
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15764 21554 15792 22102
rect 15948 21554 15976 22918
rect 16776 22778 16804 23122
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15660 21072 15712 21078
rect 15660 21014 15712 21020
rect 15672 20602 15700 21014
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15568 20392 15620 20398
rect 15566 20360 15568 20369
rect 15620 20360 15622 20369
rect 15566 20295 15622 20304
rect 15580 20262 15608 20295
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15764 19990 15792 21490
rect 16028 21412 16080 21418
rect 16028 21354 16080 21360
rect 16396 21412 16448 21418
rect 16396 21354 16448 21360
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15856 20058 15884 21082
rect 16040 20602 16068 21354
rect 16408 20942 16436 21354
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16316 20330 16344 20742
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 16212 19984 16264 19990
rect 16212 19926 16264 19932
rect 16224 19514 16252 19926
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16210 19272 16266 19281
rect 16210 19207 16266 19216
rect 15488 18958 15608 18986
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15488 18086 15516 18838
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15488 17066 15516 18022
rect 15580 17542 15608 18958
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15936 17740 15988 17746
rect 15936 17682 15988 17688
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15488 16182 15516 16526
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 14924 15972 14976 15978
rect 14924 15914 14976 15920
rect 14936 15706 14964 15914
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 14752 15366 14780 15574
rect 15488 15502 15516 16118
rect 15580 15910 15608 17478
rect 15948 17134 15976 17682
rect 16132 17202 16160 17818
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15856 16250 15884 16662
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14752 15162 14780 15302
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14476 13786 14596 13814
rect 14646 13832 14702 13841
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14384 10266 14412 10542
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14476 9081 14504 13786
rect 14646 13767 14702 13776
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 12646 14596 13262
rect 14844 12918 14872 14554
rect 15304 14498 15332 14758
rect 15396 14618 15424 15438
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15476 14884 15528 14890
rect 15476 14826 15528 14832
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15488 14498 15516 14826
rect 15304 14470 15516 14498
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 13988 15332 14470
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15384 14000 15436 14006
rect 15304 13960 15384 13988
rect 15384 13942 15436 13948
rect 15200 13932 15252 13938
rect 15252 13892 15332 13920
rect 15200 13874 15252 13880
rect 15304 13802 15332 13892
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15212 13433 15240 13738
rect 15396 13462 15424 13942
rect 15384 13456 15436 13462
rect 15198 13424 15254 13433
rect 15384 13398 15436 13404
rect 15198 13359 15254 13368
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15396 12986 15424 13398
rect 15488 13258 15516 14282
rect 15580 13258 15608 14350
rect 15856 14006 15884 14962
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15658 13832 15714 13841
rect 15658 13767 15714 13776
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14568 9926 14596 12582
rect 15384 12368 15436 12374
rect 15304 12328 15384 12356
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14740 11688 14792 11694
rect 14646 11656 14702 11665
rect 14740 11630 14792 11636
rect 14646 11591 14702 11600
rect 14660 10849 14688 11591
rect 14646 10840 14702 10849
rect 14646 10775 14702 10784
rect 14752 10742 14780 11630
rect 14844 11286 14872 12174
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11558 15332 12328
rect 15384 12310 15436 12316
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15304 11354 15332 11494
rect 15672 11370 15700 13767
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15488 11342 15700 11370
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15382 10840 15438 10849
rect 15382 10775 15438 10784
rect 15396 10742 15424 10775
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 10266 15240 10406
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 14646 10024 14702 10033
rect 14646 9959 14702 9968
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14462 9072 14518 9081
rect 14462 9007 14518 9016
rect 14292 8928 14504 8956
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14292 7478 14320 7754
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14384 7177 14412 8570
rect 14370 7168 14426 7177
rect 14370 7103 14426 7112
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14384 5846 14412 6326
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14384 4758 14412 5782
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14384 3670 14412 4150
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14476 3534 14504 8928
rect 14554 7712 14610 7721
rect 14554 7647 14610 7656
rect 14568 7546 14596 7647
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14660 7392 14688 9959
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15396 9586 15424 10066
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14568 7364 14688 7392
rect 14568 6866 14596 7364
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14568 6254 14596 6802
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 13910 54 14136 82
rect 14568 82 14596 5850
rect 14660 5370 14688 7210
rect 14752 6390 14780 7822
rect 14844 7313 14872 9454
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15120 8090 15148 8434
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15396 7410 15424 9522
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 14830 7304 14886 7313
rect 15488 7290 15516 11342
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15580 10198 15608 11086
rect 15672 10266 15700 11222
rect 15764 10538 15792 11698
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15568 10192 15620 10198
rect 15948 10146 15976 17070
rect 16118 15328 16174 15337
rect 16118 15263 16174 15272
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16040 12850 16068 13194
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16040 11150 16068 12786
rect 16132 12374 16160 15263
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 16132 11762 16160 12310
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16132 11082 16160 11698
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 15568 10134 15620 10140
rect 15672 10118 15976 10146
rect 16224 10130 16252 19207
rect 16316 18970 16344 20266
rect 16408 19854 16436 20878
rect 16500 20874 16528 21898
rect 16868 21622 16896 22510
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 16856 21616 16908 21622
rect 16856 21558 16908 21564
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 16500 20466 16528 20810
rect 16868 20466 16896 21558
rect 16960 21350 16988 21966
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 16960 20534 16988 21286
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17420 20602 17448 21082
rect 17512 21078 17540 21286
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17512 20602 17540 21014
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16408 19514 16436 19790
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16500 18290 16528 20402
rect 16868 19990 16896 20402
rect 16856 19984 16908 19990
rect 16856 19926 16908 19932
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 18970 16620 19654
rect 17130 19408 17186 19417
rect 17130 19343 17186 19352
rect 17144 19310 17172 19343
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 16592 18358 16620 18906
rect 16670 18864 16726 18873
rect 16670 18799 16726 18808
rect 17040 18828 17092 18834
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16684 18290 16712 18799
rect 17040 18770 17092 18776
rect 17052 18426 17080 18770
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16684 16794 16712 17682
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16316 13870 16344 15846
rect 16500 15706 16528 16050
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16592 15026 16620 15914
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16212 10124 16264 10130
rect 15672 7313 15700 10118
rect 16212 10066 16264 10072
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15764 8634 15792 9386
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15856 8498 15884 9998
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15948 9382 15976 9930
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9450 16160 9862
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 14830 7239 14886 7248
rect 15396 7262 15516 7290
rect 15658 7304 15714 7313
rect 15396 6866 15424 7262
rect 15658 7239 15714 7248
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 6633 15424 6802
rect 15382 6624 15438 6633
rect 14956 6556 15252 6576
rect 15382 6559 15438 6568
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 15200 6316 15252 6322
rect 15396 6304 15424 6559
rect 15252 6276 15424 6304
rect 15200 6258 15252 6264
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14740 5636 14792 5642
rect 14740 5578 14792 5584
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14752 5234 14780 5578
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14844 4826 14872 5646
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15488 5234 15516 7142
rect 15948 6769 15976 9318
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 15934 6760 15990 6769
rect 15934 6695 15990 6704
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6186 15792 6598
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15672 5030 15700 5850
rect 15764 5370 15792 6122
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 15672 4486 15700 4966
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14660 2310 14688 2926
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 14660 1737 14688 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15396 2106 15424 3470
rect 15488 3194 15516 3606
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15672 2922 15700 4422
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15948 4185 15976 4218
rect 15934 4176 15990 4185
rect 15934 4111 15990 4120
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 14646 1728 14702 1737
rect 14646 1663 14702 1672
rect 14922 82 14978 480
rect 14568 54 14978 82
rect 13910 0 13966 54
rect 14922 0 14978 54
rect 15842 82 15898 480
rect 16040 82 16068 9114
rect 16224 9110 16252 9386
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16120 8832 16172 8838
rect 16224 8820 16252 9046
rect 16172 8792 16252 8820
rect 16120 8774 16172 8780
rect 16132 8294 16160 8774
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 8090 16160 8230
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16224 7546 16252 7890
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16210 6896 16266 6905
rect 16210 6831 16266 6840
rect 16224 6798 16252 6831
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16224 6458 16252 6734
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16132 4282 16160 4694
rect 16224 4622 16252 6122
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16224 4214 16252 4558
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 16224 3670 16252 4150
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16224 2650 16252 2858
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16316 134 16344 13806
rect 16408 13161 16436 14758
rect 16394 13152 16450 13161
rect 16394 13087 16450 13096
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16408 12442 16436 12854
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16394 10840 16450 10849
rect 16394 10775 16450 10784
rect 16408 10606 16436 10775
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16500 9178 16528 14894
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16684 11014 16712 14214
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16776 10810 16804 17614
rect 16868 17066 16896 17750
rect 17052 17678 17080 18362
rect 17144 17746 17172 18906
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17236 17542 17264 17614
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17328 17218 17356 19246
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17420 18086 17448 18770
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17814 17448 18022
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17420 17338 17448 17750
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17328 17190 17448 17218
rect 16856 17060 16908 17066
rect 16856 17002 16908 17008
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17132 15088 17184 15094
rect 17132 15030 17184 15036
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16960 12714 16988 13262
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 17052 12646 17080 13398
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 16960 11558 16988 12310
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11286 16988 11494
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16960 10470 16988 11222
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16868 9042 16896 9930
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16776 8294 16804 8910
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 8022 16804 8230
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16776 6866 16804 7278
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16500 6322 16528 6598
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16408 3058 16436 3674
rect 16500 3369 16528 6258
rect 16776 6186 16804 6802
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16592 4758 16620 4966
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 16868 4154 16896 8842
rect 16960 8022 16988 10406
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17052 8634 17080 9046
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17052 8090 17080 8570
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16960 6730 16988 7278
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16776 4126 16896 4154
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16592 3670 16620 3946
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16486 3360 16542 3369
rect 16486 3295 16542 3304
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16500 2922 16528 3130
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16500 2009 16528 2382
rect 16486 2000 16542 2009
rect 16486 1935 16542 1944
rect 16776 134 16804 4126
rect 16960 3602 16988 6666
rect 17144 6458 17172 15030
rect 17236 14618 17264 15302
rect 17328 15162 17356 15574
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17236 13326 17264 13942
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17236 12730 17264 13262
rect 17328 12850 17356 14758
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17236 12702 17356 12730
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 7002 17264 12582
rect 17328 11898 17356 12702
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17314 11248 17370 11257
rect 17314 11183 17370 11192
rect 17328 11150 17356 11183
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 10266 17356 11086
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17328 8974 17356 9386
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17420 8906 17448 17190
rect 17512 16726 17540 17478
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17512 16250 17540 16662
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17512 14346 17540 15302
rect 17604 14550 17632 22918
rect 18064 22710 18092 23122
rect 18052 22704 18104 22710
rect 18052 22646 18104 22652
rect 18156 21486 18184 23598
rect 18234 23559 18290 23568
rect 18248 23526 18276 23559
rect 18236 23520 18288 23526
rect 18236 23462 18288 23468
rect 18340 23322 18368 24822
rect 18800 24138 18828 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20180 24410 20208 27520
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 21652 23866 21680 27520
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 18524 20466 18552 23802
rect 22664 23798 22692 27526
rect 23018 27520 23074 27526
rect 24228 27526 24454 27554
rect 24228 23866 24256 27526
rect 24398 27520 24454 27526
rect 25778 27520 25834 28000
rect 27158 27520 27214 28000
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24780 23866 24808 25327
rect 24858 24032 24914 24041
rect 24858 23967 24914 23976
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 22652 23792 22704 23798
rect 22652 23734 22704 23740
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19522 20496 19578 20505
rect 18512 20460 18564 20466
rect 19522 20431 19578 20440
rect 20352 20460 20404 20466
rect 18512 20402 18564 20408
rect 19536 20398 19564 20431
rect 20352 20402 20404 20408
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17696 19242 17724 19790
rect 17788 19446 17816 19926
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17972 19514 18000 19790
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17684 19236 17736 19242
rect 17684 19178 17736 19184
rect 17696 18970 17724 19178
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17788 18698 17816 19110
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17696 15638 17724 16526
rect 17684 15632 17736 15638
rect 17684 15574 17736 15580
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17604 13530 17632 14486
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17788 11558 17816 12174
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17512 9722 17540 10134
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17512 9110 17540 9658
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17328 7274 17356 7958
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17420 7002 17448 7890
rect 17604 7478 17632 10678
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 9382 17724 9998
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 7546 17724 9318
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17788 7478 17816 11494
rect 17866 10704 17922 10713
rect 17866 10639 17922 10648
rect 17880 10606 17908 10639
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17880 6934 17908 7142
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17788 6322 17816 6598
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17880 6118 17908 6190
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17144 4826 17172 5646
rect 17236 5370 17264 5782
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17132 4820 17184 4826
rect 17052 4780 17132 4808
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16960 3194 16988 3538
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17052 3058 17080 4780
rect 17132 4762 17184 4768
rect 17696 4758 17724 5578
rect 17880 5574 17908 6054
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4758 17816 4966
rect 17684 4752 17736 4758
rect 17130 4720 17186 4729
rect 17684 4694 17736 4700
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17130 4655 17186 4664
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 15842 54 16068 82
rect 16304 128 16356 134
rect 16304 70 16356 76
rect 16764 128 16816 134
rect 16764 70 16816 76
rect 16854 82 16910 480
rect 17144 82 17172 4655
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17512 4146 17540 4422
rect 17788 4282 17816 4694
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17880 4146 17908 5510
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17880 3942 17908 4082
rect 17972 4078 18000 18090
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 18064 3942 18092 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18892 19242 18920 19858
rect 18972 19304 19024 19310
rect 19432 19304 19484 19310
rect 18972 19246 19024 19252
rect 19430 19272 19432 19281
rect 19484 19272 19486 19281
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18420 18692 18472 18698
rect 18420 18634 18472 18640
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17270 18276 17478
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 18248 17066 18276 17206
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 18156 16794 18184 17002
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18340 15706 18368 17138
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18340 15026 18368 15642
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18236 14544 18288 14550
rect 18236 14486 18288 14492
rect 18248 14074 18276 14486
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18248 13802 18276 14010
rect 18432 13814 18460 18634
rect 18524 17270 18552 18702
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18512 17264 18564 17270
rect 18512 17206 18564 17212
rect 18524 14822 18552 17206
rect 18616 16114 18644 18566
rect 18800 18426 18828 18770
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18708 16998 18736 17682
rect 18800 17066 18828 18158
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18616 15706 18644 16050
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18616 15094 18644 15438
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18708 13814 18736 16934
rect 18800 16590 18828 17002
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18800 15638 18828 15914
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18800 15026 18828 15574
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18340 13786 18460 13814
rect 18616 13786 18736 13814
rect 18156 13530 18184 13738
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18248 12442 18276 13738
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18248 9722 18276 10406
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 7274 18184 8230
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 18156 6984 18184 7210
rect 18248 7206 18276 7890
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18236 6996 18288 7002
rect 18156 6956 18236 6984
rect 18236 6938 18288 6944
rect 18248 6254 18276 6938
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 18156 4826 18184 5238
rect 18340 4826 18368 13786
rect 18512 13456 18564 13462
rect 18432 13416 18512 13444
rect 18432 12714 18460 13416
rect 18512 13398 18564 13404
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18432 11354 18460 12650
rect 18524 12442 18552 13262
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18432 10266 18460 10610
rect 18616 10538 18644 13786
rect 18694 12880 18750 12889
rect 18694 12815 18750 12824
rect 18788 12844 18840 12850
rect 18708 12714 18736 12815
rect 18788 12786 18840 12792
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18800 12374 18828 12786
rect 18788 12368 18840 12374
rect 18788 12310 18840 12316
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18432 7410 18460 7890
rect 18524 7546 18552 9454
rect 18616 9042 18644 10202
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18616 8566 18644 8978
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 18708 7993 18736 9658
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18800 8294 18828 9046
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18892 7993 18920 19178
rect 18984 18834 19012 19246
rect 19430 19207 19486 19216
rect 19444 19174 19472 19207
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 17513 19012 18022
rect 18970 17504 19026 17513
rect 18970 17439 19026 17448
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 18984 15162 19012 15574
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 18984 13326 19012 13738
rect 19076 13734 19104 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 20088 18426 20116 18770
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19260 16590 19288 17546
rect 19536 17241 19564 18362
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 19522 17232 19578 17241
rect 19522 17167 19578 17176
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 16250 19288 16526
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19248 15972 19300 15978
rect 19248 15914 19300 15920
rect 19260 14890 19288 15914
rect 19352 15910 19380 16662
rect 19444 16153 19472 17070
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19430 16144 19486 16153
rect 19536 16114 19564 16934
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19984 16720 20036 16726
rect 19984 16662 20036 16668
rect 19996 16114 20024 16662
rect 20076 16176 20128 16182
rect 20076 16118 20128 16124
rect 19430 16079 19486 16088
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19536 15706 19564 16050
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19996 15638 20024 16050
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19444 14618 19472 14894
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 19064 13524 19116 13530
rect 19168 13512 19196 14350
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 19260 14006 19288 14282
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19116 13484 19196 13512
rect 19064 13466 19116 13472
rect 19260 13462 19288 13942
rect 19444 13814 19472 14554
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19996 14074 20024 14214
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19444 13802 19564 13814
rect 19996 13802 20024 14010
rect 20088 13938 20116 16118
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20180 15434 20208 16050
rect 20168 15428 20220 15434
rect 20168 15370 20220 15376
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19444 13796 19576 13802
rect 19444 13786 19524 13796
rect 19524 13738 19576 13744
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 19154 13288 19210 13297
rect 18984 12850 19012 13262
rect 19154 13223 19210 13232
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 19062 11656 19118 11665
rect 18984 11014 19012 11630
rect 19062 11591 19118 11600
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 18984 10849 19012 10950
rect 18970 10840 19026 10849
rect 18970 10775 19026 10784
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18694 7984 18750 7993
rect 18694 7919 18750 7928
rect 18878 7984 18934 7993
rect 18878 7919 18934 7928
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 18800 7002 18828 7210
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18432 5914 18460 6734
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18340 4622 18368 4762
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17788 2650 17816 2790
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 17880 2582 17908 3878
rect 18156 3398 18184 4014
rect 18248 3738 18276 4490
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 18156 2417 18184 3334
rect 18340 2854 18368 3606
rect 18420 3120 18472 3126
rect 18420 3062 18472 3068
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18340 2650 18368 2790
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 18432 2514 18460 3062
rect 18800 3058 18828 3674
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18142 2408 18198 2417
rect 18142 2343 18198 2352
rect 16854 54 17172 82
rect 17774 128 17830 480
rect 17774 76 17776 128
rect 17828 76 17830 128
rect 15842 0 15898 54
rect 16854 0 16910 54
rect 17774 0 17830 76
rect 18786 82 18842 480
rect 18892 82 18920 7919
rect 18984 5710 19012 9998
rect 19076 6866 19104 11591
rect 19168 7392 19196 13223
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 12442 19380 12582
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19444 11830 19472 12310
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 19536 11626 19564 13738
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20088 13530 20116 13874
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11286 20024 12718
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20088 11830 20116 12174
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 20088 11354 20116 11766
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19444 10538 19472 11154
rect 19432 10532 19484 10538
rect 19432 10474 19484 10480
rect 19536 10470 19564 11154
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9586 19288 9862
rect 19352 9722 19380 10134
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19524 9988 19576 9994
rect 19524 9930 19576 9936
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19260 8634 19288 9522
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19352 8838 19380 9386
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19352 8362 19380 8774
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 8090 19380 8298
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19444 7970 19472 9522
rect 19536 9042 19564 9930
rect 19996 9518 20024 10066
rect 20180 9874 20208 14962
rect 20088 9846 20208 9874
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 19536 8362 19564 8978
rect 19982 8528 20038 8537
rect 19982 8463 20038 8472
rect 19996 8362 20024 8463
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19984 8356 20036 8362
rect 19984 8298 20036 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19352 7942 19472 7970
rect 19168 7364 19288 7392
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 19076 5846 19104 6054
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 18984 5370 19012 5646
rect 19168 5642 19196 7210
rect 19156 5636 19208 5642
rect 19156 5578 19208 5584
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18984 3670 19012 4558
rect 19076 4214 19104 5034
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18984 3058 19012 3606
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 19168 2514 19196 5578
rect 19260 5234 19288 7364
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19246 4176 19302 4185
rect 19246 4111 19302 4120
rect 19260 3602 19288 4111
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19352 3534 19380 7942
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19536 7002 19564 7346
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19628 6254 19656 6802
rect 19982 6352 20038 6361
rect 19982 6287 20038 6296
rect 19996 6254 20024 6287
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19444 6118 19472 6190
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5846 20024 6190
rect 19616 5840 19668 5846
rect 19616 5782 19668 5788
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19444 4865 19472 5646
rect 19628 5370 19656 5782
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19430 4856 19486 4865
rect 19622 4848 19918 4868
rect 19430 4791 19486 4800
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19720 4593 19748 4626
rect 19706 4584 19762 4593
rect 19706 4519 19762 4528
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19444 4146 19472 4218
rect 19720 4214 19748 4519
rect 20088 4486 20116 9846
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19708 4208 19760 4214
rect 19708 4150 19760 4156
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19248 2916 19300 2922
rect 19444 2904 19472 4082
rect 20088 4010 20116 4082
rect 19892 4004 19944 4010
rect 20076 4004 20128 4010
rect 19944 3964 20024 3992
rect 19892 3946 19944 3952
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19996 3670 20024 3964
rect 20076 3946 20128 3952
rect 19984 3664 20036 3670
rect 19984 3606 20036 3612
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 19812 3194 19840 3538
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19300 2876 19472 2904
rect 19248 2858 19300 2864
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 20180 1873 20208 9658
rect 20272 9586 20300 17478
rect 20364 17134 20392 20402
rect 20534 19408 20590 19417
rect 20534 19343 20590 19352
rect 20548 19310 20576 19343
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20364 14346 20392 17070
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20364 11354 20392 13670
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20364 10674 20392 11290
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20364 10130 20392 10610
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20456 10062 20484 18702
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20548 16266 20576 18158
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20640 16454 20668 18022
rect 20996 17740 21048 17746
rect 20996 17682 21048 17688
rect 20902 17232 20958 17241
rect 21008 17202 21036 17682
rect 20902 17167 20958 17176
rect 20996 17196 21048 17202
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20548 16238 20668 16266
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20548 14618 20576 14894
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20548 12374 20576 14418
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20534 12200 20590 12209
rect 20534 12135 20590 12144
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20272 8634 20300 9318
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20364 8566 20392 9590
rect 20548 9353 20576 12135
rect 20640 9761 20668 16238
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20732 14482 20760 14894
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20824 12442 20852 15642
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20916 12322 20944 17167
rect 20996 17138 21048 17144
rect 21100 16794 21128 23462
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21100 16250 21128 16594
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 21100 15434 21128 16186
rect 21192 15502 21220 18022
rect 21284 17785 21312 23598
rect 21928 23474 21956 23598
rect 21836 23446 21956 23474
rect 22376 23520 22428 23526
rect 22376 23462 22428 23468
rect 21454 21040 21510 21049
rect 21454 20975 21510 20984
rect 21270 17776 21326 17785
rect 21270 17711 21326 17720
rect 21364 17060 21416 17066
rect 21364 17002 21416 17008
rect 21272 15632 21324 15638
rect 21272 15574 21324 15580
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 21192 15094 21220 15438
rect 21284 15162 21312 15574
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14414 21036 14758
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 21008 13530 21036 14350
rect 21100 14074 21128 14486
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 21008 12782 21036 13126
rect 21192 12850 21220 14826
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20824 12294 20944 12322
rect 20996 12368 21048 12374
rect 20996 12310 21048 12316
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11762 20760 12038
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20732 9926 20760 10406
rect 20824 10130 20852 12294
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20916 11694 20944 12174
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20916 11354 20944 11630
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20916 10742 20944 11154
rect 20904 10736 20956 10742
rect 20904 10678 20956 10684
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20626 9752 20682 9761
rect 20626 9687 20682 9696
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20534 9344 20590 9353
rect 20534 9279 20590 9288
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20272 7002 20300 7210
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20364 5846 20392 6190
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20364 4185 20392 4490
rect 20350 4176 20406 4185
rect 20350 4111 20406 4120
rect 20456 3738 20484 8910
rect 20640 8634 20668 9454
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20640 7342 20668 7482
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20732 5710 20760 9862
rect 20824 9722 20852 10066
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20916 9654 20944 10678
rect 20904 9648 20956 9654
rect 20904 9590 20956 9596
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20720 4752 20772 4758
rect 20824 4729 20852 7414
rect 20720 4694 20772 4700
rect 20810 4720 20866 4729
rect 20732 3942 20760 4694
rect 21008 4690 21036 12310
rect 21100 7478 21128 12378
rect 21192 11558 21220 12786
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21284 12442 21312 12582
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21284 11626 21312 12378
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21192 10266 21220 10474
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 21284 10198 21312 10474
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21192 8498 21220 8774
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 21088 7472 21140 7478
rect 21088 7414 21140 7420
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 21192 7206 21220 7278
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21100 5370 21128 6054
rect 21192 5681 21220 7142
rect 21284 5896 21312 9998
rect 21376 8974 21404 17002
rect 21468 15638 21496 20975
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21640 15428 21692 15434
rect 21640 15370 21692 15376
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21468 13326 21496 14350
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21560 13938 21588 14282
rect 21652 13938 21680 15370
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21560 12986 21588 13398
rect 21652 13326 21680 13874
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21376 6934 21404 7142
rect 21364 6928 21416 6934
rect 21364 6870 21416 6876
rect 21376 6118 21404 6870
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21284 5868 21404 5896
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 21178 5672 21234 5681
rect 21178 5607 21234 5616
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 21100 5098 21128 5306
rect 21088 5092 21140 5098
rect 21088 5034 21140 5040
rect 21100 4758 21128 5034
rect 21284 4826 21312 5714
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21088 4752 21140 4758
rect 21088 4694 21140 4700
rect 20810 4655 20866 4664
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20166 1864 20222 1873
rect 20166 1799 20222 1808
rect 18786 54 18920 82
rect 19706 96 19762 480
rect 18786 0 18842 54
rect 20456 82 20484 3334
rect 21008 2922 21036 3878
rect 21100 3738 21128 4558
rect 21376 4264 21404 5868
rect 21284 4236 21404 4264
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 21284 3194 21312 4236
rect 21468 4154 21496 12718
rect 21560 11898 21588 12922
rect 21652 12306 21680 13262
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21560 10810 21588 11086
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21560 8401 21588 9454
rect 21744 9058 21772 17478
rect 21836 17202 21864 23446
rect 22388 22506 22416 23462
rect 22376 22500 22428 22506
rect 22376 22442 22428 22448
rect 22008 21480 22060 21486
rect 22008 21422 22060 21428
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 22020 16250 22048 21422
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 21914 16144 21970 16153
rect 21914 16079 21970 16088
rect 21928 15586 21956 16079
rect 22020 16046 22048 16186
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 22020 15706 22048 15982
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 21928 15558 22048 15586
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21928 14521 21956 15302
rect 21914 14512 21970 14521
rect 21914 14447 21970 14456
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21836 13802 21864 14214
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21836 12442 21864 13738
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21836 10452 21864 11494
rect 22020 11150 22048 15558
rect 22112 15502 22140 16594
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22112 15337 22140 15438
rect 22098 15328 22154 15337
rect 22098 15263 22154 15272
rect 22100 13252 22152 13258
rect 22100 13194 22152 13200
rect 22112 12442 22140 13194
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22204 11778 22232 15846
rect 22296 12782 22324 16390
rect 22388 13938 22416 22442
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23492 20369 23520 22374
rect 23938 21176 23994 21185
rect 23938 21111 23994 21120
rect 23478 20360 23534 20369
rect 23478 20295 23534 20304
rect 23112 19304 23164 19310
rect 23112 19246 23164 19252
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 15026 22508 17478
rect 22572 17134 22600 17682
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22480 14074 22508 14418
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22296 12442 22324 12582
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22296 11898 22324 12378
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22100 11756 22152 11762
rect 22204 11750 22324 11778
rect 22100 11698 22152 11704
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22112 10470 22140 11698
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22204 10606 22232 10950
rect 22192 10600 22244 10606
rect 22296 10577 22324 11750
rect 22192 10542 22244 10548
rect 22282 10568 22338 10577
rect 22100 10464 22152 10470
rect 21836 10424 21956 10452
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21836 9586 21864 10202
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21836 9110 21864 9318
rect 21652 9030 21772 9058
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21546 8392 21602 8401
rect 21546 8327 21602 8336
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21560 7750 21588 8230
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21560 7206 21588 7686
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21560 6254 21588 6598
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21560 5914 21588 6190
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21376 4126 21496 4154
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 20996 2916 21048 2922
rect 20996 2858 21048 2864
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 21284 2650 21312 2858
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21376 2446 21404 4126
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21468 3602 21496 3946
rect 21652 3754 21680 9030
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21744 7818 21772 8910
rect 21836 8294 21864 9046
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21836 8022 21864 8230
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21732 7812 21784 7818
rect 21732 7754 21784 7760
rect 21744 7206 21772 7754
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 21928 5273 21956 10424
rect 22100 10406 22152 10412
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 22020 8974 22048 9386
rect 22112 9178 22140 9998
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 22204 7342 22232 10542
rect 22282 10503 22338 10512
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22296 9382 22324 10202
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22296 5846 22324 6734
rect 22284 5840 22336 5846
rect 22284 5782 22336 5788
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22204 5370 22232 5646
rect 22296 5574 22324 5782
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22388 5386 22416 12106
rect 22480 11801 22508 14010
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22572 12374 22600 12582
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22466 11792 22522 11801
rect 22466 11727 22522 11736
rect 22572 11354 22600 12310
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22572 7002 22600 7822
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22480 5846 22508 6054
rect 22468 5840 22520 5846
rect 22468 5782 22520 5788
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22296 5358 22416 5386
rect 21914 5264 21970 5273
rect 21914 5199 21970 5208
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22112 4758 22140 4966
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22020 4282 22048 4422
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 22020 4154 22048 4218
rect 22020 4126 22140 4154
rect 22112 4010 22140 4126
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 21652 3726 21864 3754
rect 21732 3664 21784 3670
rect 21732 3606 21784 3612
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 21744 2854 21772 3606
rect 21836 3534 21864 3726
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 21744 2582 21772 2790
rect 21836 2650 21864 3470
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 22020 2582 22048 3946
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22204 3466 22232 3878
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 22296 3126 22324 5358
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 22284 3120 22336 3126
rect 22284 3062 22336 3068
rect 21732 2576 21784 2582
rect 21454 2544 21510 2553
rect 21732 2518 21784 2524
rect 22008 2576 22060 2582
rect 22008 2518 22060 2524
rect 21454 2479 21510 2488
rect 21468 2446 21496 2479
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 22008 2372 22060 2378
rect 22008 2314 22060 2320
rect 20718 82 20774 480
rect 20456 54 20774 82
rect 19706 0 19762 40
rect 20718 0 20774 54
rect 21638 82 21694 480
rect 22020 82 22048 2314
rect 21638 54 22048 82
rect 22388 82 22416 5238
rect 22480 4826 22508 5782
rect 22664 5710 22692 16526
rect 22940 16046 22968 16594
rect 22928 16040 22980 16046
rect 22926 16008 22928 16017
rect 22980 16008 22982 16017
rect 22926 15943 22982 15952
rect 22940 15910 22968 15943
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22940 15570 22968 15846
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 22940 15162 22968 15506
rect 23124 15162 23152 19246
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23124 14958 23152 15098
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22928 14340 22980 14346
rect 22928 14282 22980 14288
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22756 10130 22784 13806
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22848 12714 22876 13398
rect 22836 12708 22888 12714
rect 22836 12650 22888 12656
rect 22940 12238 22968 14282
rect 23032 13734 23060 14418
rect 23020 13728 23072 13734
rect 23020 13670 23072 13676
rect 23216 13433 23244 14758
rect 23202 13424 23258 13433
rect 23202 13359 23258 13368
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23032 12986 23060 13262
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 22940 11665 22968 11698
rect 23020 11688 23072 11694
rect 22926 11656 22982 11665
rect 23020 11630 23072 11636
rect 22926 11591 22982 11600
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22848 9450 22876 10610
rect 23032 10554 23060 11630
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 23124 10606 23152 11562
rect 22940 10526 23060 10554
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 22848 8974 22876 9386
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22744 8288 22796 8294
rect 22744 8230 22796 8236
rect 22756 8022 22784 8230
rect 22744 8016 22796 8022
rect 22744 7958 22796 7964
rect 22848 7546 22876 8570
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 22848 7342 22876 7482
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22940 7206 22968 10526
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 23032 9722 23060 10406
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23124 9042 23152 9998
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23112 7268 23164 7274
rect 23112 7210 23164 7216
rect 22928 7200 22980 7206
rect 22928 7142 22980 7148
rect 23124 6458 23152 7210
rect 23216 6798 23244 12378
rect 23308 8974 23336 17070
rect 23492 14498 23520 20295
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23584 16998 23612 17682
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23400 14470 23520 14498
rect 23400 10742 23428 14470
rect 23480 13728 23532 13734
rect 23584 13705 23612 16934
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23676 13870 23704 14214
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23756 13728 23808 13734
rect 23480 13670 23532 13676
rect 23570 13696 23626 13705
rect 23492 11626 23520 13670
rect 23756 13670 23808 13676
rect 23570 13631 23626 13640
rect 23584 13297 23612 13631
rect 23768 13530 23796 13670
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23570 13288 23626 13297
rect 23570 13223 23626 13232
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23584 11694 23612 12038
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 23480 11620 23532 11626
rect 23480 11562 23532 11568
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23492 10470 23520 11222
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23584 10282 23612 11630
rect 23676 11150 23704 12582
rect 23860 12442 23888 15642
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23952 11830 23980 21111
rect 24228 18970 24256 23666
rect 24872 23322 24900 23967
rect 25792 23633 25820 27520
rect 27172 23730 27200 27520
rect 27618 27296 27674 27305
rect 27618 27231 27674 27240
rect 27632 24886 27660 27231
rect 27620 24880 27672 24886
rect 27620 24822 27672 24828
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 25778 23624 25834 23633
rect 25778 23559 25834 23568
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22438 24716 23122
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24780 21690 24808 22471
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24766 19816 24822 19825
rect 24766 19751 24822 19760
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24780 19514 24808 19751
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 24136 18086 24164 18770
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24766 18320 24822 18329
rect 24766 18255 24822 18264
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 24136 17513 24164 18022
rect 24122 17504 24178 17513
rect 24122 17439 24178 17448
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24780 17338 24808 18255
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24582 17232 24638 17241
rect 24582 17167 24638 17176
rect 24596 17134 24624 17167
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24766 16960 24822 16969
rect 24766 16895 24822 16904
rect 24676 16516 24728 16522
rect 24676 16458 24728 16464
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 24032 14884 24084 14890
rect 24032 14826 24084 14832
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23756 11552 23808 11558
rect 23756 11494 23808 11500
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23492 10254 23612 10282
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23400 9042 23428 9590
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23400 8362 23428 8978
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23400 7857 23428 8298
rect 23386 7848 23442 7857
rect 23386 7783 23442 7792
rect 23492 7342 23520 10254
rect 23572 10192 23624 10198
rect 23676 10180 23704 11086
rect 23768 10849 23796 11494
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23754 10840 23810 10849
rect 23754 10775 23810 10784
rect 23756 10532 23808 10538
rect 23860 10520 23888 10950
rect 23808 10492 23888 10520
rect 23756 10474 23808 10480
rect 23624 10152 23704 10180
rect 23848 10192 23900 10198
rect 23572 10134 23624 10140
rect 23848 10134 23900 10140
rect 23860 9722 23888 10134
rect 23952 10062 23980 11018
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 23848 9716 23900 9722
rect 23848 9658 23900 9664
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 23584 9178 23612 9318
rect 24044 9178 24072 14826
rect 24228 14822 24256 15506
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24124 13728 24176 13734
rect 24124 13670 24176 13676
rect 24136 13161 24164 13670
rect 24122 13152 24178 13161
rect 24122 13087 24178 13096
rect 24228 10282 24256 14758
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 13870 24716 16458
rect 24780 16250 24808 16895
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24766 15600 24822 15609
rect 24766 15535 24822 15544
rect 24780 14618 24808 15535
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24872 14482 24900 16390
rect 25148 15570 25176 21422
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25240 15910 25268 16594
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25136 15564 25188 15570
rect 25136 15506 25188 15512
rect 25148 15162 25176 15506
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24872 14074 24900 14418
rect 24950 14240 25006 14249
rect 24950 14175 25006 14184
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24780 13394 24808 13874
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24780 12646 24808 13330
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24584 12300 24636 12306
rect 24636 12260 24716 12288
rect 24584 12242 24636 12248
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12260
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24400 10600 24452 10606
rect 24400 10542 24452 10548
rect 24136 10254 24256 10282
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23388 7336 23440 7342
rect 23388 7278 23440 7284
rect 23480 7336 23532 7342
rect 23480 7278 23532 7284
rect 23400 7206 23428 7278
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23400 6905 23428 7142
rect 23386 6896 23442 6905
rect 23386 6831 23442 6840
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23308 6361 23336 6394
rect 23294 6352 23350 6361
rect 23294 6287 23350 6296
rect 23308 6254 23336 6287
rect 23296 6248 23348 6254
rect 23296 6190 23348 6196
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 23202 5672 23258 5681
rect 22664 5370 22692 5646
rect 22744 5636 22796 5642
rect 23202 5607 23258 5616
rect 22744 5578 22796 5584
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 22756 5166 22784 5578
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22756 4826 22784 5102
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 22652 4752 22704 4758
rect 22652 4694 22704 4700
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22480 3602 22508 4082
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22572 3534 22600 4626
rect 22664 3738 22692 4694
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22940 4146 22968 4558
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 23216 4078 23244 5607
rect 23400 5370 23428 6831
rect 23584 6458 23612 8910
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23478 6352 23534 6361
rect 23478 6287 23480 6296
rect 23532 6287 23534 6296
rect 23480 6258 23532 6264
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23400 5166 23428 5306
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22664 3194 22692 3334
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22756 3058 22784 3674
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 23308 3398 23336 3538
rect 23296 3392 23348 3398
rect 22834 3360 22890 3369
rect 23296 3334 23348 3340
rect 22834 3295 22890 3304
rect 22848 3194 22876 3295
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 23110 3088 23166 3097
rect 22744 3052 22796 3058
rect 23110 3023 23166 3032
rect 22744 2994 22796 3000
rect 23124 2990 23152 3023
rect 23112 2984 23164 2990
rect 23112 2926 23164 2932
rect 23308 2854 23336 3334
rect 23492 3194 23520 6258
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23584 5778 23612 6190
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23584 5030 23612 5510
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23676 4154 23704 8910
rect 23860 8634 23888 8978
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23768 7206 23796 8434
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23860 8090 23888 8298
rect 24044 8294 24072 9114
rect 24136 8974 24164 10254
rect 24412 10198 24440 10542
rect 24400 10192 24452 10198
rect 24228 10152 24400 10180
rect 24228 9586 24256 10152
rect 24400 10134 24452 10140
rect 24780 10033 24808 12582
rect 24872 10130 24900 13806
rect 24964 12986 24992 14175
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 24964 12782 24992 12922
rect 24952 12776 25004 12782
rect 25148 12753 25176 15098
rect 24952 12718 25004 12724
rect 25134 12744 25190 12753
rect 25134 12679 25190 12688
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24964 11257 24992 11290
rect 24950 11248 25006 11257
rect 24950 11183 25006 11192
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24964 10470 24992 11086
rect 25148 10674 25176 11154
rect 25136 10668 25188 10674
rect 25136 10610 25188 10616
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 24766 10024 24822 10033
rect 24766 9959 24822 9968
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24124 8968 24176 8974
rect 24124 8910 24176 8916
rect 24228 8498 24256 9522
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 23940 8016 23992 8022
rect 23940 7958 23992 7964
rect 23846 7848 23902 7857
rect 23846 7783 23902 7792
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23768 6118 23796 6598
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23768 5166 23796 5510
rect 23756 5160 23808 5166
rect 23756 5102 23808 5108
rect 23860 4690 23888 7783
rect 23952 7002 23980 7958
rect 24228 7818 24256 8434
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7449 24716 9318
rect 24674 7440 24730 7449
rect 24674 7375 24730 7384
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 24044 6712 24072 6870
rect 23952 6684 24072 6712
rect 23952 5846 23980 6684
rect 24030 6624 24086 6633
rect 24030 6559 24086 6568
rect 24044 6322 24072 6559
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 24136 6254 24164 7210
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24780 6390 24808 7142
rect 24872 6934 24900 9658
rect 24964 7410 24992 10406
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 25056 8430 25084 9590
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 25056 7546 25084 7822
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24952 6996 25004 7002
rect 24952 6938 25004 6944
rect 24860 6928 24912 6934
rect 24860 6870 24912 6876
rect 24768 6384 24820 6390
rect 24768 6326 24820 6332
rect 24124 6248 24176 6254
rect 24124 6190 24176 6196
rect 23940 5840 23992 5846
rect 23940 5782 23992 5788
rect 23952 4758 23980 5782
rect 24124 5772 24176 5778
rect 24124 5714 24176 5720
rect 24136 5370 24164 5714
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24124 5364 24176 5370
rect 24124 5306 24176 5312
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24124 5160 24176 5166
rect 24124 5102 24176 5108
rect 24136 4758 24164 5102
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 24124 4752 24176 4758
rect 24124 4694 24176 4700
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23952 4214 23980 4694
rect 23584 4126 23704 4154
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 23584 2514 23612 4126
rect 24136 4078 24164 4694
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4282 24716 4626
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3670 23796 3878
rect 23756 3664 23808 3670
rect 23756 3606 23808 3612
rect 24780 3602 24808 5238
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23664 3120 23716 3126
rect 23664 3062 23716 3068
rect 23572 2508 23624 2514
rect 23572 2450 23624 2456
rect 23112 2372 23164 2378
rect 23112 2314 23164 2320
rect 23124 2106 23152 2314
rect 23112 2100 23164 2106
rect 23112 2042 23164 2048
rect 23676 1601 23704 3062
rect 23768 1737 23796 3470
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 23940 3120 23992 3126
rect 23940 3062 23992 3068
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23754 1728 23810 1737
rect 23754 1663 23810 1672
rect 23662 1592 23718 1601
rect 23662 1527 23718 1536
rect 22650 82 22706 480
rect 22388 54 22706 82
rect 21638 0 21694 54
rect 22650 0 22706 54
rect 23570 82 23626 480
rect 23860 82 23888 2926
rect 23952 2650 23980 3062
rect 24044 3058 24072 3334
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 24044 1465 24072 2994
rect 24136 2961 24164 2994
rect 24122 2952 24178 2961
rect 24122 2887 24178 2896
rect 24216 2848 24268 2854
rect 24216 2790 24268 2796
rect 24124 2644 24176 2650
rect 24124 2586 24176 2592
rect 24136 2417 24164 2586
rect 24228 2514 24256 2790
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24122 2408 24178 2417
rect 24122 2343 24178 2352
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24030 1456 24086 1465
rect 24030 1391 24086 1400
rect 23570 54 23888 82
rect 24582 82 24638 480
rect 24872 82 24900 4150
rect 24964 2009 24992 6938
rect 25148 6866 25176 10610
rect 25240 9722 25268 15846
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25700 13705 25728 13806
rect 25686 13696 25742 13705
rect 25686 13631 25742 13640
rect 25594 13016 25650 13025
rect 25594 12951 25650 12960
rect 25608 12918 25636 12951
rect 25596 12912 25648 12918
rect 25596 12854 25648 12860
rect 25412 12300 25464 12306
rect 25412 12242 25464 12248
rect 25424 11558 25452 12242
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25226 9616 25282 9625
rect 25226 9551 25282 9560
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25148 6769 25176 6802
rect 25134 6760 25190 6769
rect 25134 6695 25190 6704
rect 25148 6390 25176 6695
rect 25136 6384 25188 6390
rect 25136 6326 25188 6332
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 25148 4486 25176 5510
rect 25240 5166 25268 9551
rect 25332 9042 25360 11018
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 25332 8294 25360 8978
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 25136 4480 25188 4486
rect 25136 4422 25188 4428
rect 25044 3596 25096 3602
rect 25044 3538 25096 3544
rect 25056 3194 25084 3538
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 25332 2514 25360 8230
rect 25424 6866 25452 11494
rect 25516 10810 25544 11630
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25596 10736 25648 10742
rect 25596 10678 25648 10684
rect 25608 7954 25636 10678
rect 26056 10124 26108 10130
rect 26056 10066 26108 10072
rect 26068 9722 26096 10066
rect 27528 9920 27580 9926
rect 27528 9862 27580 9868
rect 26056 9716 26108 9722
rect 26056 9658 26108 9664
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 25700 7993 25728 9454
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25686 7984 25742 7993
rect 25596 7948 25648 7954
rect 25686 7919 25742 7928
rect 25596 7890 25648 7896
rect 25608 7546 25636 7890
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 25424 5574 25452 6802
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 24950 2000 25006 2009
rect 24950 1935 25006 1944
rect 24582 54 24900 82
rect 25424 82 25452 4966
rect 25792 4146 25820 8230
rect 26608 6384 26660 6390
rect 26608 6326 26660 6332
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25516 3602 25544 3878
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25516 2854 25544 3538
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 25516 2650 25544 2790
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 25502 82 25558 480
rect 25424 54 25558 82
rect 23570 0 23626 54
rect 24582 0 24638 54
rect 25502 0 25558 54
rect 26514 82 26570 480
rect 26620 82 26648 6326
rect 26514 54 26648 82
rect 27434 82 27490 480
rect 27540 82 27568 9862
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 27632 785 27660 6394
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27724 2145 27752 2246
rect 27710 2136 27766 2145
rect 27710 2071 27766 2080
rect 27618 776 27674 785
rect 27618 711 27674 720
rect 27434 54 27568 82
rect 26514 0 26570 54
rect 27434 0 27490 54
<< via2 >>
rect 1122 26696 1178 26752
rect 1582 25336 1638 25392
rect 1214 23976 1270 24032
rect 1582 22480 1638 22536
rect 1122 21120 1178 21176
rect 1030 13096 1086 13152
rect 1030 8200 1086 8256
rect 110 3440 166 3496
rect 1582 19760 1638 19816
rect 1582 18264 1638 18320
rect 1582 16904 1638 16960
rect 1582 15544 1638 15600
rect 1490 15272 1546 15328
rect 2042 19080 2098 19136
rect 1674 7384 1730 7440
rect 1490 6160 1546 6216
rect 1674 5772 1730 5808
rect 1674 5752 1676 5772
rect 1676 5752 1728 5772
rect 1728 5752 1730 5772
rect 1214 2624 1270 2680
rect 1674 1808 1730 1864
rect 2042 16088 2098 16144
rect 2226 13912 2282 13968
rect 2134 11056 2190 11112
rect 1950 8880 2006 8936
rect 2778 15408 2834 15464
rect 2686 14476 2742 14512
rect 2686 14456 2688 14476
rect 2688 14456 2740 14476
rect 2740 14456 2742 14476
rect 2686 13776 2742 13832
rect 2778 13232 2834 13288
rect 2318 10648 2374 10704
rect 1858 3984 1914 4040
rect 2870 10648 2926 10704
rect 2778 8472 2834 8528
rect 2778 8336 2834 8392
rect 2686 6704 2742 6760
rect 3882 21392 3938 21448
rect 3146 15952 3202 16008
rect 3054 13368 3110 13424
rect 3146 11192 3202 11248
rect 3238 7248 3294 7304
rect 3146 6976 3202 7032
rect 3146 6704 3202 6760
rect 2134 1672 2190 1728
rect 2042 1264 2098 1320
rect 3422 6160 3478 6216
rect 3330 3848 3386 3904
rect 3790 17040 3846 17096
rect 3790 13912 3846 13968
rect 3882 13776 3938 13832
rect 4802 19760 4858 19816
rect 3698 9560 3754 9616
rect 3606 9324 3608 9344
rect 3608 9324 3660 9344
rect 3660 9324 3662 9344
rect 3606 9288 3662 9324
rect 3606 5636 3662 5672
rect 3606 5616 3608 5636
rect 3608 5616 3660 5636
rect 3660 5616 3662 5636
rect 4434 13232 4490 13288
rect 3882 9560 3938 9616
rect 4526 11736 4582 11792
rect 3974 9424 4030 9480
rect 3882 9288 3938 9344
rect 4158 6860 4214 6896
rect 4158 6840 4160 6860
rect 4160 6840 4212 6860
rect 4212 6840 4214 6860
rect 4066 4800 4122 4856
rect 3882 3440 3938 3496
rect 3238 2488 3294 2544
rect 3146 1944 3202 2000
rect 4802 6296 4858 6352
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 7194 23296 7250 23352
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5262 13912 5318 13968
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5998 14048 6054 14104
rect 5446 13776 5502 13832
rect 5998 13776 6054 13832
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5998 4256 6054 4312
rect 6550 14048 6606 14104
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 8114 21664 8170 21720
rect 7654 19080 7710 19136
rect 7102 13232 7158 13288
rect 7010 7656 7066 7712
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6458 3848 6514 3904
rect 7654 12824 7710 12880
rect 8574 22072 8630 22128
rect 8942 20476 8944 20496
rect 8944 20476 8996 20496
rect 8996 20476 8998 20496
rect 8942 20440 8998 20476
rect 9494 20984 9550 21040
rect 8942 19080 8998 19136
rect 8666 17720 8722 17776
rect 8574 11056 8630 11112
rect 7838 9560 7894 9616
rect 8390 7928 8446 7984
rect 8298 7384 8354 7440
rect 8850 12416 8906 12472
rect 8850 10648 8906 10704
rect 8850 9016 8906 9072
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10690 15408 10746 15464
rect 9218 12144 9274 12200
rect 9586 12280 9642 12336
rect 9034 10784 9090 10840
rect 9126 8472 9182 8528
rect 8850 3984 8906 4040
rect 8942 3712 8998 3768
rect 8942 3032 8998 3088
rect 8758 2488 8814 2544
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10230 9424 10286 9480
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 9310 4800 9366 4856
rect 9862 4800 9918 4856
rect 9402 4392 9458 4448
rect 9494 3848 9550 3904
rect 9954 4256 10010 4312
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10322 6704 10378 6760
rect 10322 6160 10378 6216
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10506 5616 10562 5672
rect 11794 14456 11850 14512
rect 11610 13912 11666 13968
rect 11242 13232 11298 13288
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10874 2624 10930 2680
rect 9954 40 10010 96
rect 10690 1536 10746 1592
rect 11794 12688 11850 12744
rect 11978 11056 12034 11112
rect 11978 10512 12034 10568
rect 11978 9696 12034 9752
rect 12438 21392 12494 21448
rect 12622 19216 12678 19272
rect 12530 14048 12586 14104
rect 12070 8336 12126 8392
rect 12530 8472 12586 8528
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 13358 19760 13414 19816
rect 13082 18808 13138 18864
rect 12898 12280 12954 12336
rect 12346 5616 12402 5672
rect 13082 11192 13138 11248
rect 13818 21664 13874 21720
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14002 20984 14058 21040
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14646 20440 14702 20496
rect 14002 17720 14058 17776
rect 13542 9016 13598 9072
rect 11610 4800 11666 4856
rect 11886 4392 11942 4448
rect 11610 3440 11666 3496
rect 12714 1944 12770 2000
rect 11794 1400 11850 1456
rect 13174 5752 13230 5808
rect 12990 2896 13046 2952
rect 13910 10648 13966 10704
rect 13726 8336 13782 8392
rect 13726 7384 13782 7440
rect 14278 14456 14334 14512
rect 13542 3440 13598 3496
rect 13266 1672 13322 1728
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15566 20340 15568 20360
rect 15568 20340 15620 20360
rect 15620 20340 15622 20360
rect 15566 20304 15622 20340
rect 16210 19216 16266 19272
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14646 13776 14702 13832
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15198 13368 15254 13424
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15658 13776 15714 13832
rect 14646 11600 14702 11656
rect 14646 10784 14702 10840
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15382 10784 15438 10840
rect 14646 9968 14702 10024
rect 14462 9016 14518 9072
rect 14370 7112 14426 7168
rect 14554 7656 14610 7712
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14830 7248 14886 7304
rect 16118 15272 16174 15328
rect 17130 19352 17186 19408
rect 16670 18808 16726 18864
rect 15658 7248 15714 7304
rect 15382 6568 15438 6624
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15934 6704 15990 6760
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15934 4120 15990 4176
rect 14646 1672 14702 1728
rect 16210 6840 16266 6896
rect 16394 13096 16450 13152
rect 16394 10784 16450 10840
rect 16486 3304 16542 3360
rect 16486 1944 16542 2000
rect 17314 11192 17370 11248
rect 18234 23568 18290 23624
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 24766 25336 24822 25392
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24858 23976 24914 24032
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19522 20440 19578 20496
rect 17866 10648 17922 10704
rect 17130 4664 17186 4720
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19430 19252 19432 19272
rect 19432 19252 19484 19272
rect 19484 19252 19486 19272
rect 18694 12824 18750 12880
rect 19430 19216 19486 19252
rect 18970 17448 19026 17504
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19522 17176 19578 17232
rect 19430 16088 19486 16144
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19154 13232 19210 13288
rect 19062 11600 19118 11656
rect 18970 10784 19026 10840
rect 18694 7928 18750 7984
rect 18878 7928 18934 7984
rect 18142 2352 18198 2408
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19982 8472 20038 8528
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19246 4120 19302 4176
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19982 6296 20038 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19430 4800 19486 4856
rect 19706 4528 19762 4584
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20534 19352 20590 19408
rect 20902 17176 20958 17232
rect 20534 12144 20590 12200
rect 21454 20984 21510 21040
rect 21270 17720 21326 17776
rect 20626 9696 20682 9752
rect 20534 9288 20590 9344
rect 20350 4120 20406 4176
rect 20810 4664 20866 4720
rect 21178 5616 21234 5672
rect 20166 1808 20222 1864
rect 19706 40 19762 96
rect 21914 16088 21970 16144
rect 21914 14456 21970 14512
rect 22098 15272 22154 15328
rect 23938 21120 23994 21176
rect 23478 20304 23534 20360
rect 21546 8336 21602 8392
rect 22282 10512 22338 10568
rect 22466 11736 22522 11792
rect 21914 5208 21970 5264
rect 21454 2488 21510 2544
rect 22926 15988 22928 16008
rect 22928 15988 22980 16008
rect 22980 15988 22982 16008
rect 22926 15952 22982 15988
rect 23202 13368 23258 13424
rect 22926 11600 22982 11656
rect 23570 13640 23626 13696
rect 23570 13232 23626 13288
rect 27618 27240 27674 27296
rect 25778 23568 25834 23624
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 22480 24822 22536
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 19760 24822 19816
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24766 18264 24822 18320
rect 24122 17448 24178 17504
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24582 17176 24638 17232
rect 24766 16904 24822 16960
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 23386 7792 23442 7848
rect 23754 10784 23810 10840
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24122 13096 24178 13152
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 15544 24822 15600
rect 24950 14184 25006 14240
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 23386 6840 23442 6896
rect 23294 6296 23350 6352
rect 23202 5616 23258 5672
rect 23478 6316 23534 6352
rect 23478 6296 23480 6316
rect 23480 6296 23532 6316
rect 23532 6296 23534 6316
rect 22834 3304 22890 3360
rect 23110 3032 23166 3088
rect 25134 12688 25190 12744
rect 24950 11192 25006 11248
rect 24766 9968 24822 10024
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 23846 7792 23902 7848
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24674 7384 24730 7440
rect 24030 6568 24086 6624
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 23754 1672 23810 1728
rect 23662 1536 23718 1592
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24122 2896 24178 2952
rect 24122 2352 24178 2408
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24030 1400 24086 1456
rect 25686 13640 25742 13696
rect 25594 12960 25650 13016
rect 25226 9560 25282 9616
rect 25134 6704 25190 6760
rect 25686 7928 25742 7984
rect 24950 1944 25006 2000
rect 27710 2080 27766 2136
rect 27618 720 27674 776
<< metal3 >>
rect 0 27208 480 27328
rect 27520 27296 28000 27328
rect 27520 27240 27618 27296
rect 27674 27240 28000 27296
rect 27520 27208 28000 27240
rect 62 26754 122 27208
rect 1117 26754 1183 26757
rect 62 26752 1183 26754
rect 62 26696 1122 26752
rect 1178 26696 1183 26752
rect 62 26694 1183 26696
rect 1117 26691 1183 26694
rect 0 25848 480 25968
rect 27520 25848 28000 25968
rect 62 25394 122 25848
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 1577 25394 1643 25397
rect 62 25392 1643 25394
rect 62 25336 1582 25392
rect 1638 25336 1643 25392
rect 62 25334 1643 25336
rect 1577 25331 1643 25334
rect 24761 25394 24827 25397
rect 27662 25394 27722 25848
rect 24761 25392 27722 25394
rect 24761 25336 24766 25392
rect 24822 25336 27722 25392
rect 24761 25334 27722 25336
rect 24761 25331 24827 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24488 480 24608
rect 10277 24512 10597 24513
rect 62 24034 122 24488
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 27520 24488 28000 24608
rect 19610 24447 19930 24448
rect 1209 24034 1275 24037
rect 62 24032 1275 24034
rect 62 23976 1214 24032
rect 1270 23976 1275 24032
rect 62 23974 1275 23976
rect 1209 23971 1275 23974
rect 24853 24034 24919 24037
rect 27662 24034 27722 24488
rect 24853 24032 27722 24034
rect 24853 23976 24858 24032
rect 24914 23976 27722 24032
rect 24853 23974 27722 23976
rect 24853 23971 24919 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 18229 23626 18295 23629
rect 25773 23626 25839 23629
rect 18229 23624 25839 23626
rect 18229 23568 18234 23624
rect 18290 23568 25778 23624
rect 25834 23568 25839 23624
rect 18229 23566 25839 23568
rect 18229 23563 18295 23566
rect 25773 23563 25839 23566
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 2998 23292 3004 23356
rect 3068 23354 3074 23356
rect 7189 23354 7255 23357
rect 3068 23352 7255 23354
rect 3068 23296 7194 23352
rect 7250 23296 7255 23352
rect 3068 23294 7255 23296
rect 3068 23292 3074 23294
rect 7189 23291 7255 23294
rect 0 22992 480 23112
rect 27520 22992 28000 23112
rect 62 22538 122 22992
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1577 22538 1643 22541
rect 62 22536 1643 22538
rect 62 22480 1582 22536
rect 1638 22480 1643 22536
rect 62 22478 1643 22480
rect 1577 22475 1643 22478
rect 24761 22538 24827 22541
rect 27662 22538 27722 22992
rect 24761 22536 27722 22538
rect 24761 22480 24766 22536
rect 24822 22480 27722 22536
rect 24761 22478 27722 22480
rect 24761 22475 24827 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 8569 22130 8635 22133
rect 11094 22130 11100 22132
rect 8569 22128 11100 22130
rect 8569 22072 8574 22128
rect 8630 22072 11100 22128
rect 8569 22070 11100 22072
rect 8569 22067 8635 22070
rect 11094 22068 11100 22070
rect 11164 22068 11170 22132
rect 5610 21792 5930 21793
rect 0 21632 480 21752
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 8109 21722 8175 21725
rect 13813 21722 13879 21725
rect 8109 21720 13879 21722
rect 8109 21664 8114 21720
rect 8170 21664 13818 21720
rect 13874 21664 13879 21720
rect 8109 21662 13879 21664
rect 8109 21659 8175 21662
rect 13813 21659 13879 21662
rect 27520 21632 28000 21752
rect 62 21178 122 21632
rect 3877 21450 3943 21453
rect 12433 21450 12499 21453
rect 3877 21448 12499 21450
rect 3877 21392 3882 21448
rect 3938 21392 12438 21448
rect 12494 21392 12499 21448
rect 3877 21390 12499 21392
rect 3877 21387 3943 21390
rect 12433 21387 12499 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1117 21178 1183 21181
rect 62 21176 1183 21178
rect 62 21120 1122 21176
rect 1178 21120 1183 21176
rect 62 21118 1183 21120
rect 1117 21115 1183 21118
rect 23933 21178 23999 21181
rect 27662 21178 27722 21632
rect 23933 21176 27722 21178
rect 23933 21120 23938 21176
rect 23994 21120 27722 21176
rect 23933 21118 27722 21120
rect 23933 21115 23999 21118
rect 9489 21042 9555 21045
rect 13997 21042 14063 21045
rect 21449 21042 21515 21045
rect 9489 21040 21515 21042
rect 9489 20984 9494 21040
rect 9550 20984 14002 21040
rect 14058 20984 21454 21040
rect 21510 20984 21515 21040
rect 9489 20982 21515 20984
rect 9489 20979 9555 20982
rect 13997 20979 14063 20982
rect 21449 20979 21515 20982
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 8937 20498 9003 20501
rect 14641 20498 14707 20501
rect 19517 20498 19583 20501
rect 8937 20496 19583 20498
rect 8937 20440 8942 20496
rect 8998 20440 14646 20496
rect 14702 20440 19522 20496
rect 19578 20440 19583 20496
rect 8937 20438 19583 20440
rect 8937 20435 9003 20438
rect 14641 20435 14707 20438
rect 19517 20435 19583 20438
rect 0 20272 480 20392
rect 15561 20362 15627 20365
rect 23473 20362 23539 20365
rect 15561 20360 23539 20362
rect 15561 20304 15566 20360
rect 15622 20304 23478 20360
rect 23534 20304 23539 20360
rect 15561 20302 23539 20304
rect 15561 20299 15627 20302
rect 23473 20299 23539 20302
rect 27520 20272 28000 20392
rect 62 19818 122 20272
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1577 19818 1643 19821
rect 62 19816 1643 19818
rect 62 19760 1582 19816
rect 1638 19760 1643 19816
rect 62 19758 1643 19760
rect 1577 19755 1643 19758
rect 4797 19818 4863 19821
rect 13353 19818 13419 19821
rect 4797 19816 13419 19818
rect 4797 19760 4802 19816
rect 4858 19760 13358 19816
rect 13414 19760 13419 19816
rect 4797 19758 13419 19760
rect 4797 19755 4863 19758
rect 13353 19755 13419 19758
rect 24761 19818 24827 19821
rect 27662 19818 27722 20272
rect 24761 19816 27722 19818
rect 24761 19760 24766 19816
rect 24822 19760 27722 19816
rect 24761 19758 27722 19760
rect 24761 19755 24827 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 17125 19410 17191 19413
rect 20529 19410 20595 19413
rect 17125 19408 20595 19410
rect 17125 19352 17130 19408
rect 17186 19352 20534 19408
rect 20590 19352 20595 19408
rect 17125 19350 20595 19352
rect 17125 19347 17191 19350
rect 20529 19347 20595 19350
rect 12617 19274 12683 19277
rect 16205 19274 16271 19277
rect 19425 19274 19491 19277
rect 12617 19272 19491 19274
rect 12617 19216 12622 19272
rect 12678 19216 16210 19272
rect 16266 19216 19430 19272
rect 19486 19216 19491 19272
rect 12617 19214 19491 19216
rect 12617 19211 12683 19214
rect 16205 19211 16271 19214
rect 19425 19211 19491 19214
rect 2037 19138 2103 19141
rect 7649 19138 7715 19141
rect 8937 19138 9003 19141
rect 2037 19136 9003 19138
rect 2037 19080 2042 19136
rect 2098 19080 7654 19136
rect 7710 19080 8942 19136
rect 8998 19080 9003 19136
rect 2037 19078 9003 19080
rect 2037 19075 2103 19078
rect 7649 19075 7715 19078
rect 8937 19075 9003 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 0 18776 480 18896
rect 13077 18866 13143 18869
rect 16665 18866 16731 18869
rect 13077 18864 16731 18866
rect 13077 18808 13082 18864
rect 13138 18808 16670 18864
rect 16726 18808 16731 18864
rect 13077 18806 16731 18808
rect 13077 18803 13143 18806
rect 16665 18803 16731 18806
rect 27520 18776 28000 18896
rect 62 18322 122 18776
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 1577 18322 1643 18325
rect 62 18320 1643 18322
rect 62 18264 1582 18320
rect 1638 18264 1643 18320
rect 62 18262 1643 18264
rect 1577 18259 1643 18262
rect 24761 18322 24827 18325
rect 27662 18322 27722 18776
rect 24761 18320 27722 18322
rect 24761 18264 24766 18320
rect 24822 18264 27722 18320
rect 24761 18262 27722 18264
rect 24761 18259 24827 18262
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 8661 17778 8727 17781
rect 13997 17778 14063 17781
rect 21265 17778 21331 17781
rect 8661 17776 21331 17778
rect 8661 17720 8666 17776
rect 8722 17720 14002 17776
rect 14058 17720 21270 17776
rect 21326 17720 21331 17776
rect 8661 17718 21331 17720
rect 8661 17715 8727 17718
rect 13997 17715 14063 17718
rect 21265 17715 21331 17718
rect 0 17416 480 17536
rect 18965 17506 19031 17509
rect 24117 17506 24183 17509
rect 18965 17504 24183 17506
rect 18965 17448 18970 17504
rect 19026 17448 24122 17504
rect 24178 17448 24183 17504
rect 18965 17446 24183 17448
rect 18965 17443 19031 17446
rect 24117 17443 24183 17446
rect 5610 17440 5930 17441
rect 62 16962 122 17416
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17536
rect 24277 17375 24597 17376
rect 19517 17234 19583 17237
rect 20897 17234 20963 17237
rect 24577 17234 24643 17237
rect 19517 17232 24643 17234
rect 19517 17176 19522 17232
rect 19578 17176 20902 17232
rect 20958 17176 24582 17232
rect 24638 17176 24643 17232
rect 19517 17174 24643 17176
rect 19517 17171 19583 17174
rect 20897 17171 20963 17174
rect 24577 17171 24643 17174
rect 3366 17036 3372 17100
rect 3436 17098 3442 17100
rect 3785 17098 3851 17101
rect 3436 17096 3851 17098
rect 3436 17040 3790 17096
rect 3846 17040 3851 17096
rect 3436 17038 3851 17040
rect 3436 17036 3442 17038
rect 3785 17035 3851 17038
rect 1577 16962 1643 16965
rect 62 16960 1643 16962
rect 62 16904 1582 16960
rect 1638 16904 1643 16960
rect 62 16902 1643 16904
rect 1577 16899 1643 16902
rect 24761 16962 24827 16965
rect 27662 16962 27722 17416
rect 24761 16960 27722 16962
rect 24761 16904 24766 16960
rect 24822 16904 27722 16960
rect 24761 16902 27722 16904
rect 24761 16899 24827 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16056 480 16176
rect 2037 16146 2103 16149
rect 19425 16146 19491 16149
rect 21909 16146 21975 16149
rect 2037 16144 21975 16146
rect 2037 16088 2042 16144
rect 2098 16088 19430 16144
rect 19486 16088 21914 16144
rect 21970 16088 21975 16144
rect 2037 16086 21975 16088
rect 2037 16083 2103 16086
rect 19425 16083 19491 16086
rect 21909 16083 21975 16086
rect 27520 16056 28000 16176
rect 62 15602 122 16056
rect 3141 16010 3207 16013
rect 22921 16010 22987 16013
rect 3141 16008 22987 16010
rect 3141 15952 3146 16008
rect 3202 15952 22926 16008
rect 22982 15952 22987 16008
rect 3141 15950 22987 15952
rect 3141 15947 3207 15950
rect 22921 15947 22987 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 1577 15602 1643 15605
rect 62 15600 1643 15602
rect 62 15544 1582 15600
rect 1638 15544 1643 15600
rect 62 15542 1643 15544
rect 1577 15539 1643 15542
rect 24761 15602 24827 15605
rect 27662 15602 27722 16056
rect 24761 15600 27722 15602
rect 24761 15544 24766 15600
rect 24822 15544 27722 15600
rect 24761 15542 27722 15544
rect 24761 15539 24827 15542
rect 2773 15466 2839 15469
rect 10685 15466 10751 15469
rect 2773 15464 10751 15466
rect 2773 15408 2778 15464
rect 2834 15408 10690 15464
rect 10746 15408 10751 15464
rect 2773 15406 10751 15408
rect 2773 15403 2839 15406
rect 10685 15403 10751 15406
rect 1485 15330 1551 15333
rect 62 15328 1551 15330
rect 62 15272 1490 15328
rect 1546 15272 1551 15328
rect 62 15270 1551 15272
rect 62 14816 122 15270
rect 1485 15267 1551 15270
rect 16113 15330 16179 15333
rect 22093 15330 22159 15333
rect 16113 15328 22159 15330
rect 16113 15272 16118 15328
rect 16174 15272 22098 15328
rect 22154 15272 22159 15328
rect 16113 15270 22159 15272
rect 16113 15267 16179 15270
rect 22093 15267 22159 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14696 480 14816
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 27520 14696 28000 14816
rect 19610 14655 19930 14656
rect 2681 14514 2747 14517
rect 11789 14514 11855 14517
rect 2681 14512 11855 14514
rect 2681 14456 2686 14512
rect 2742 14456 11794 14512
rect 11850 14456 11855 14512
rect 2681 14454 11855 14456
rect 2681 14451 2747 14454
rect 11789 14451 11855 14454
rect 14273 14514 14339 14517
rect 21909 14514 21975 14517
rect 14273 14512 21975 14514
rect 14273 14456 14278 14512
rect 14334 14456 21914 14512
rect 21970 14456 21975 14512
rect 14273 14454 21975 14456
rect 14273 14451 14339 14454
rect 21909 14451 21975 14454
rect 24945 14242 25011 14245
rect 27662 14242 27722 14696
rect 24945 14240 27722 14242
rect 24945 14184 24950 14240
rect 25006 14184 27722 14240
rect 24945 14182 27722 14184
rect 24945 14179 25011 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 5993 14106 6059 14109
rect 6545 14106 6611 14109
rect 12525 14106 12591 14109
rect 5993 14104 12591 14106
rect 5993 14048 5998 14104
rect 6054 14048 6550 14104
rect 6606 14048 12530 14104
rect 12586 14048 12591 14104
rect 5993 14046 12591 14048
rect 5993 14043 6059 14046
rect 6545 14043 6611 14046
rect 12525 14043 12591 14046
rect 2221 13970 2287 13973
rect 3785 13970 3851 13973
rect 2221 13968 3851 13970
rect 2221 13912 2226 13968
rect 2282 13912 3790 13968
rect 3846 13912 3851 13968
rect 2221 13910 3851 13912
rect 2221 13907 2287 13910
rect 3785 13907 3851 13910
rect 5257 13970 5323 13973
rect 11605 13970 11671 13973
rect 5257 13968 11671 13970
rect 5257 13912 5262 13968
rect 5318 13912 11610 13968
rect 11666 13912 11671 13968
rect 5257 13910 11671 13912
rect 5257 13907 5323 13910
rect 11605 13907 11671 13910
rect 2446 13772 2452 13836
rect 2516 13834 2522 13836
rect 2681 13834 2747 13837
rect 2516 13832 2747 13834
rect 2516 13776 2686 13832
rect 2742 13776 2747 13832
rect 2516 13774 2747 13776
rect 2516 13772 2522 13774
rect 2681 13771 2747 13774
rect 3877 13832 3943 13837
rect 3877 13776 3882 13832
rect 3938 13776 3943 13832
rect 3877 13771 3943 13776
rect 5441 13834 5507 13837
rect 5993 13834 6059 13837
rect 5441 13832 6059 13834
rect 5441 13776 5446 13832
rect 5502 13776 5998 13832
rect 6054 13776 6059 13832
rect 5441 13774 6059 13776
rect 5441 13771 5507 13774
rect 5993 13771 6059 13774
rect 14641 13834 14707 13837
rect 15653 13834 15719 13837
rect 14641 13832 15719 13834
rect 14641 13776 14646 13832
rect 14702 13776 15658 13832
rect 15714 13776 15719 13832
rect 14641 13774 15719 13776
rect 14641 13771 14707 13774
rect 15653 13771 15719 13774
rect 3880 13700 3940 13771
rect 3880 13638 3924 13700
rect 3918 13636 3924 13638
rect 3988 13636 3994 13700
rect 23565 13698 23631 13701
rect 25681 13698 25747 13701
rect 23565 13696 25747 13698
rect 23565 13640 23570 13696
rect 23626 13640 25686 13696
rect 25742 13640 25747 13696
rect 23565 13638 25747 13640
rect 23565 13635 23631 13638
rect 25681 13635 25747 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3049 13426 3115 13429
rect 15193 13426 15259 13429
rect 23197 13426 23263 13429
rect 3049 13424 13830 13426
rect 3049 13368 3054 13424
rect 3110 13368 13830 13424
rect 3049 13366 13830 13368
rect 3049 13363 3115 13366
rect 0 13200 480 13320
rect 2773 13290 2839 13293
rect 3182 13290 3188 13292
rect 2773 13288 3188 13290
rect 2773 13232 2778 13288
rect 2834 13232 3188 13288
rect 2773 13230 3188 13232
rect 2773 13227 2839 13230
rect 3182 13228 3188 13230
rect 3252 13228 3258 13292
rect 4429 13290 4495 13293
rect 7097 13290 7163 13293
rect 11237 13290 11303 13293
rect 4429 13288 11303 13290
rect 4429 13232 4434 13288
rect 4490 13232 7102 13288
rect 7158 13232 11242 13288
rect 11298 13232 11303 13288
rect 4429 13230 11303 13232
rect 13770 13290 13830 13366
rect 15193 13424 23263 13426
rect 15193 13368 15198 13424
rect 15254 13368 23202 13424
rect 23258 13368 23263 13424
rect 15193 13366 23263 13368
rect 15193 13363 15259 13366
rect 23197 13363 23263 13366
rect 19149 13290 19215 13293
rect 23565 13290 23631 13293
rect 13770 13288 23631 13290
rect 13770 13232 19154 13288
rect 19210 13232 23570 13288
rect 23626 13232 23631 13288
rect 13770 13230 23631 13232
rect 4429 13227 4495 13230
rect 7097 13227 7163 13230
rect 11237 13227 11303 13230
rect 19149 13227 19215 13230
rect 23565 13227 23631 13230
rect 27520 13200 28000 13320
rect 62 12474 122 13200
rect 1025 13154 1091 13157
rect 3918 13154 3924 13156
rect 1025 13152 3924 13154
rect 1025 13096 1030 13152
rect 1086 13096 3924 13152
rect 1025 13094 3924 13096
rect 1025 13091 1091 13094
rect 3918 13092 3924 13094
rect 3988 13154 3994 13156
rect 16389 13154 16455 13157
rect 24117 13154 24183 13157
rect 3988 13094 4170 13154
rect 3988 13092 3994 13094
rect 4110 12746 4170 13094
rect 16389 13152 24183 13154
rect 16389 13096 16394 13152
rect 16450 13096 24122 13152
rect 24178 13096 24183 13152
rect 16389 13094 24183 13096
rect 16389 13091 16455 13094
rect 24117 13091 24183 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 25589 13018 25655 13021
rect 27662 13018 27722 13200
rect 25589 13016 27722 13018
rect 25589 12960 25594 13016
rect 25650 12960 27722 13016
rect 25589 12958 27722 12960
rect 25589 12955 25655 12958
rect 7649 12882 7715 12885
rect 18689 12882 18755 12885
rect 7649 12880 18755 12882
rect 7649 12824 7654 12880
rect 7710 12824 18694 12880
rect 18750 12824 18755 12880
rect 7649 12822 18755 12824
rect 7649 12819 7715 12822
rect 18689 12819 18755 12822
rect 11789 12746 11855 12749
rect 25129 12746 25195 12749
rect 4110 12744 25195 12746
rect 4110 12688 11794 12744
rect 11850 12688 25134 12744
rect 25190 12688 25195 12744
rect 4110 12686 25195 12688
rect 11789 12683 11855 12686
rect 25129 12683 25195 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 8845 12474 8911 12477
rect 62 12472 8911 12474
rect 62 12416 8850 12472
rect 8906 12416 8911 12472
rect 62 12414 8911 12416
rect 8845 12411 8911 12414
rect 9581 12338 9647 12341
rect 12893 12338 12959 12341
rect 62 12336 12959 12338
rect 62 12280 9586 12336
rect 9642 12280 12898 12336
rect 12954 12280 12959 12336
rect 62 12278 12959 12280
rect 62 11960 122 12278
rect 9581 12275 9647 12278
rect 12893 12275 12959 12278
rect 9213 12202 9279 12205
rect 20529 12202 20595 12205
rect 9213 12200 20595 12202
rect 9213 12144 9218 12200
rect 9274 12144 20534 12200
rect 20590 12144 20595 12200
rect 9213 12142 20595 12144
rect 9213 12139 9279 12142
rect 20529 12139 20595 12142
rect 5610 12000 5930 12001
rect 0 11840 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 27520 11840 28000 11960
rect 4521 11794 4587 11797
rect 20110 11794 20116 11796
rect 4521 11792 20116 11794
rect 4521 11736 4526 11792
rect 4582 11736 20116 11792
rect 4521 11734 20116 11736
rect 4521 11731 4587 11734
rect 20110 11732 20116 11734
rect 20180 11794 20186 11796
rect 22461 11794 22527 11797
rect 20180 11792 22527 11794
rect 20180 11736 22466 11792
rect 22522 11736 22527 11792
rect 20180 11734 22527 11736
rect 20180 11732 20186 11734
rect 22461 11731 22527 11734
rect 14641 11658 14707 11661
rect 19057 11658 19123 11661
rect 22921 11658 22987 11661
rect 14641 11656 22987 11658
rect 14641 11600 14646 11656
rect 14702 11600 19062 11656
rect 19118 11600 22926 11656
rect 22982 11600 22987 11656
rect 14641 11598 22987 11600
rect 14641 11595 14707 11598
rect 19057 11595 19123 11598
rect 22921 11595 22987 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3141 11250 3207 11253
rect 13077 11250 13143 11253
rect 3141 11248 13143 11250
rect 3141 11192 3146 11248
rect 3202 11192 13082 11248
rect 13138 11192 13143 11248
rect 3141 11190 13143 11192
rect 3141 11187 3207 11190
rect 13077 11187 13143 11190
rect 17309 11250 17375 11253
rect 24945 11250 25011 11253
rect 17309 11248 25011 11250
rect 17309 11192 17314 11248
rect 17370 11192 24950 11248
rect 25006 11192 25011 11248
rect 17309 11190 25011 11192
rect 17309 11187 17375 11190
rect 24945 11187 25011 11190
rect 2129 11114 2195 11117
rect 8569 11114 8635 11117
rect 2129 11112 8635 11114
rect 2129 11056 2134 11112
rect 2190 11056 8574 11112
rect 8630 11056 8635 11112
rect 2129 11054 8635 11056
rect 2129 11051 2195 11054
rect 8569 11051 8635 11054
rect 11973 11114 12039 11117
rect 27662 11114 27722 11840
rect 11973 11112 27722 11114
rect 11973 11056 11978 11112
rect 12034 11056 27722 11112
rect 11973 11054 27722 11056
rect 11973 11051 12039 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 9029 10842 9095 10845
rect 14641 10842 14707 10845
rect 8710 10840 9095 10842
rect 8710 10784 9034 10840
rect 9090 10784 9095 10840
rect 8710 10782 9095 10784
rect 2313 10706 2379 10709
rect 2865 10706 2931 10709
rect 8710 10706 8770 10782
rect 9029 10779 9095 10782
rect 13770 10840 14707 10842
rect 13770 10784 14646 10840
rect 14702 10784 14707 10840
rect 13770 10782 14707 10784
rect 2313 10704 8770 10706
rect 2313 10648 2318 10704
rect 2374 10648 2870 10704
rect 2926 10648 8770 10704
rect 2313 10646 8770 10648
rect 8845 10706 8911 10709
rect 13770 10706 13830 10782
rect 14641 10779 14707 10782
rect 15377 10842 15443 10845
rect 16389 10842 16455 10845
rect 15377 10840 16455 10842
rect 15377 10784 15382 10840
rect 15438 10784 16394 10840
rect 16450 10784 16455 10840
rect 15377 10782 16455 10784
rect 15377 10779 15443 10782
rect 16389 10779 16455 10782
rect 18965 10842 19031 10845
rect 23749 10842 23815 10845
rect 18965 10840 23815 10842
rect 18965 10784 18970 10840
rect 19026 10784 23754 10840
rect 23810 10784 23815 10840
rect 18965 10782 23815 10784
rect 18965 10779 19031 10782
rect 23749 10779 23815 10782
rect 8845 10704 13830 10706
rect 8845 10648 8850 10704
rect 8906 10648 13830 10704
rect 8845 10646 13830 10648
rect 13905 10706 13971 10709
rect 17861 10706 17927 10709
rect 13905 10704 17927 10706
rect 13905 10648 13910 10704
rect 13966 10648 17866 10704
rect 17922 10648 17927 10704
rect 13905 10646 17927 10648
rect 2313 10643 2379 10646
rect 2865 10643 2931 10646
rect 8845 10643 8911 10646
rect 13905 10643 13971 10646
rect 17861 10643 17927 10646
rect 0 10480 480 10600
rect 11973 10570 12039 10573
rect 22277 10570 22343 10573
rect 27520 10570 28000 10600
rect 11973 10568 28000 10570
rect 11973 10512 11978 10568
rect 12034 10512 22282 10568
rect 22338 10512 28000 10568
rect 11973 10510 28000 10512
rect 11973 10507 12039 10510
rect 22277 10507 22343 10510
rect 27520 10480 28000 10510
rect 62 10026 122 10480
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 14641 10026 14707 10029
rect 24761 10026 24827 10029
rect 62 10024 24827 10026
rect 62 9968 14646 10024
rect 14702 9968 24766 10024
rect 24822 9968 24827 10024
rect 62 9966 24827 9968
rect 14641 9963 14707 9966
rect 24761 9963 24827 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 11094 9692 11100 9756
rect 11164 9754 11170 9756
rect 11973 9754 12039 9757
rect 11164 9752 12039 9754
rect 11164 9696 11978 9752
rect 12034 9696 12039 9752
rect 11164 9694 12039 9696
rect 11164 9692 11170 9694
rect 11973 9691 12039 9694
rect 20621 9754 20687 9757
rect 20621 9752 23490 9754
rect 20621 9696 20626 9752
rect 20682 9696 23490 9752
rect 20621 9694 23490 9696
rect 20621 9691 20687 9694
rect 3693 9618 3759 9621
rect 3877 9618 3943 9621
rect 7833 9618 7899 9621
rect 3693 9616 3802 9618
rect 3693 9560 3698 9616
rect 3754 9560 3802 9616
rect 3693 9555 3802 9560
rect 3877 9616 7899 9618
rect 3877 9560 3882 9616
rect 3938 9560 7838 9616
rect 7894 9560 7899 9616
rect 3877 9558 7899 9560
rect 23430 9618 23490 9694
rect 25221 9618 25287 9621
rect 23430 9616 25287 9618
rect 23430 9560 25226 9616
rect 25282 9560 25287 9616
rect 23430 9558 25287 9560
rect 3877 9555 3943 9558
rect 7833 9555 7899 9558
rect 25221 9555 25287 9558
rect 3182 9284 3188 9348
rect 3252 9346 3258 9348
rect 3601 9346 3667 9349
rect 3252 9344 3667 9346
rect 3252 9288 3606 9344
rect 3662 9288 3667 9344
rect 3252 9286 3667 9288
rect 3742 9346 3802 9555
rect 3969 9482 4035 9485
rect 10225 9482 10291 9485
rect 3969 9480 10291 9482
rect 3969 9424 3974 9480
rect 4030 9424 10230 9480
rect 10286 9424 10291 9480
rect 3969 9422 10291 9424
rect 3969 9419 4035 9422
rect 10225 9419 10291 9422
rect 3877 9346 3943 9349
rect 3742 9344 3943 9346
rect 3742 9288 3882 9344
rect 3938 9288 3943 9344
rect 3742 9286 3943 9288
rect 3252 9284 3258 9286
rect 3601 9283 3667 9286
rect 3877 9283 3943 9286
rect 20529 9346 20595 9349
rect 20529 9344 27722 9346
rect 20529 9288 20534 9344
rect 20590 9288 27722 9344
rect 20529 9286 27722 9288
rect 20529 9283 20595 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 27662 9104 27722 9286
rect 0 9076 480 9104
rect 0 9012 60 9076
rect 124 9012 480 9076
rect 0 8984 480 9012
rect 8845 9074 8911 9077
rect 13537 9074 13603 9077
rect 14457 9074 14523 9077
rect 8845 9072 13603 9074
rect 8845 9016 8850 9072
rect 8906 9016 13542 9072
rect 13598 9016 13603 9072
rect 8845 9014 13603 9016
rect 8845 9011 8911 9014
rect 13537 9011 13603 9014
rect 13770 9072 14523 9074
rect 13770 9016 14462 9072
rect 14518 9016 14523 9072
rect 13770 9014 14523 9016
rect 1945 8938 2011 8941
rect 13770 8938 13830 9014
rect 14457 9011 14523 9014
rect 27520 8984 28000 9104
rect 614 8936 13830 8938
rect 614 8880 1950 8936
rect 2006 8880 13830 8936
rect 614 8878 13830 8880
rect 54 8740 60 8804
rect 124 8802 130 8804
rect 614 8802 674 8878
rect 1945 8875 2011 8878
rect 124 8742 674 8802
rect 124 8740 130 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 2773 8530 2839 8533
rect 9121 8530 9187 8533
rect 2773 8528 9187 8530
rect 2773 8472 2778 8528
rect 2834 8472 9126 8528
rect 9182 8472 9187 8528
rect 2773 8470 9187 8472
rect 2773 8467 2839 8470
rect 9121 8467 9187 8470
rect 12525 8530 12591 8533
rect 19977 8530 20043 8533
rect 12525 8528 20043 8530
rect 12525 8472 12530 8528
rect 12586 8472 19982 8528
rect 20038 8472 20043 8528
rect 12525 8470 20043 8472
rect 12525 8467 12591 8470
rect 19977 8467 20043 8470
rect 2773 8394 2839 8397
rect 12065 8394 12131 8397
rect 2773 8392 12131 8394
rect 2773 8336 2778 8392
rect 2834 8336 12070 8392
rect 12126 8336 12131 8392
rect 2773 8334 12131 8336
rect 2773 8331 2839 8334
rect 12065 8331 12131 8334
rect 13721 8394 13787 8397
rect 21541 8394 21607 8397
rect 13721 8392 21607 8394
rect 13721 8336 13726 8392
rect 13782 8336 21546 8392
rect 21602 8336 21607 8392
rect 13721 8334 21607 8336
rect 13721 8331 13787 8334
rect 21541 8331 21607 8334
rect 1025 8258 1091 8261
rect 62 8256 1091 8258
rect 62 8200 1030 8256
rect 1086 8200 1091 8256
rect 62 8198 1091 8200
rect 62 7744 122 8198
rect 1025 8195 1091 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 8385 7986 8451 7989
rect 18689 7986 18755 7989
rect 8385 7984 18755 7986
rect 8385 7928 8390 7984
rect 8446 7928 18694 7984
rect 18750 7928 18755 7984
rect 8385 7926 18755 7928
rect 8385 7923 8451 7926
rect 18689 7923 18755 7926
rect 18873 7986 18939 7989
rect 25681 7986 25747 7989
rect 18873 7984 25747 7986
rect 18873 7928 18878 7984
rect 18934 7928 25686 7984
rect 25742 7928 25747 7984
rect 18873 7926 25747 7928
rect 18873 7923 18939 7926
rect 25681 7923 25747 7926
rect 23381 7850 23447 7853
rect 23841 7850 23907 7853
rect 23381 7848 23907 7850
rect 23381 7792 23386 7848
rect 23442 7792 23846 7848
rect 23902 7792 23907 7848
rect 23381 7790 23907 7792
rect 23381 7787 23447 7790
rect 23841 7787 23907 7790
rect 0 7624 480 7744
rect 7005 7714 7071 7717
rect 14549 7714 14615 7717
rect 7005 7712 14615 7714
rect 7005 7656 7010 7712
rect 7066 7656 14554 7712
rect 14610 7656 14615 7712
rect 7005 7654 14615 7656
rect 7005 7651 7071 7654
rect 14549 7651 14615 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7744
rect 24277 7583 24597 7584
rect 1669 7442 1735 7445
rect 8293 7442 8359 7445
rect 1669 7440 8359 7442
rect 1669 7384 1674 7440
rect 1730 7384 8298 7440
rect 8354 7384 8359 7440
rect 1669 7382 8359 7384
rect 1669 7379 1735 7382
rect 8293 7379 8359 7382
rect 13721 7442 13787 7445
rect 24669 7442 24735 7445
rect 13721 7440 24735 7442
rect 13721 7384 13726 7440
rect 13782 7384 24674 7440
rect 24730 7384 24735 7440
rect 13721 7382 24735 7384
rect 13721 7379 13787 7382
rect 24669 7379 24735 7382
rect 3233 7306 3299 7309
rect 14825 7306 14891 7309
rect 15653 7306 15719 7309
rect 27662 7306 27722 7624
rect 3233 7304 14891 7306
rect 3233 7248 3238 7304
rect 3294 7248 14830 7304
rect 14886 7248 14891 7304
rect 3233 7246 14891 7248
rect 3233 7243 3299 7246
rect 14825 7243 14891 7246
rect 14966 7304 27722 7306
rect 14966 7248 15658 7304
rect 15714 7248 27722 7304
rect 14966 7246 27722 7248
rect 14365 7170 14431 7173
rect 14966 7170 15026 7246
rect 15653 7243 15719 7246
rect 14365 7168 15026 7170
rect 14365 7112 14370 7168
rect 14426 7112 15026 7168
rect 14365 7110 15026 7112
rect 14365 7107 14431 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 2998 6972 3004 7036
rect 3068 7034 3074 7036
rect 3141 7034 3207 7037
rect 3068 7032 3207 7034
rect 3068 6976 3146 7032
rect 3202 6976 3207 7032
rect 3068 6974 3207 6976
rect 3068 6972 3074 6974
rect 3141 6971 3207 6974
rect 4153 6898 4219 6901
rect 16205 6898 16271 6901
rect 23381 6898 23447 6901
rect 4153 6896 23447 6898
rect 4153 6840 4158 6896
rect 4214 6840 16210 6896
rect 16266 6840 23386 6896
rect 23442 6840 23447 6896
rect 4153 6838 23447 6840
rect 4153 6835 4219 6838
rect 16205 6835 16271 6838
rect 23381 6835 23447 6838
rect 2446 6762 2452 6764
rect 62 6702 2452 6762
rect 62 6384 122 6702
rect 2446 6700 2452 6702
rect 2516 6700 2522 6764
rect 2681 6762 2747 6765
rect 3141 6762 3207 6765
rect 2681 6760 3207 6762
rect 2681 6704 2686 6760
rect 2742 6704 3146 6760
rect 3202 6704 3207 6760
rect 2681 6702 3207 6704
rect 2681 6699 2747 6702
rect 3141 6699 3207 6702
rect 10317 6762 10383 6765
rect 15929 6762 15995 6765
rect 25129 6762 25195 6765
rect 10317 6760 25195 6762
rect 10317 6704 10322 6760
rect 10378 6704 15934 6760
rect 15990 6704 25134 6760
rect 25190 6704 25195 6760
rect 10317 6702 25195 6704
rect 10317 6699 10383 6702
rect 15929 6699 15995 6702
rect 25129 6699 25195 6702
rect 15377 6626 15443 6629
rect 24025 6626 24091 6629
rect 15377 6624 24091 6626
rect 15377 6568 15382 6624
rect 15438 6568 24030 6624
rect 24086 6568 24091 6624
rect 15377 6566 24091 6568
rect 15377 6563 15443 6566
rect 24025 6563 24091 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6264 480 6384
rect 3366 6292 3372 6356
rect 3436 6354 3442 6356
rect 4797 6354 4863 6357
rect 3436 6352 4863 6354
rect 3436 6296 4802 6352
rect 4858 6296 4863 6352
rect 3436 6294 4863 6296
rect 3436 6292 3442 6294
rect 4797 6291 4863 6294
rect 19977 6354 20043 6357
rect 20110 6354 20116 6356
rect 19977 6352 20116 6354
rect 19977 6296 19982 6352
rect 20038 6296 20116 6352
rect 19977 6294 20116 6296
rect 19977 6291 20043 6294
rect 20110 6292 20116 6294
rect 20180 6354 20186 6356
rect 23289 6354 23355 6357
rect 20180 6352 23355 6354
rect 20180 6296 23294 6352
rect 23350 6296 23355 6352
rect 20180 6294 23355 6296
rect 20180 6292 20186 6294
rect 23289 6291 23355 6294
rect 23473 6354 23539 6357
rect 27520 6354 28000 6384
rect 23473 6352 28000 6354
rect 23473 6296 23478 6352
rect 23534 6296 28000 6352
rect 23473 6294 28000 6296
rect 23473 6291 23539 6294
rect 27520 6264 28000 6294
rect 1485 6218 1551 6221
rect 3417 6218 3483 6221
rect 10317 6218 10383 6221
rect 1485 6216 10383 6218
rect 1485 6160 1490 6216
rect 1546 6160 3422 6216
rect 3478 6160 10322 6216
rect 10378 6160 10383 6216
rect 1485 6158 10383 6160
rect 1485 6155 1551 6158
rect 3417 6155 3483 6158
rect 10317 6155 10383 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 1669 5810 1735 5813
rect 13169 5810 13235 5813
rect 1669 5808 13235 5810
rect 1669 5752 1674 5808
rect 1730 5752 13174 5808
rect 13230 5752 13235 5808
rect 1669 5750 13235 5752
rect 1669 5747 1735 5750
rect 13169 5747 13235 5750
rect 3601 5674 3667 5677
rect 10501 5674 10567 5677
rect 3601 5672 10567 5674
rect 3601 5616 3606 5672
rect 3662 5616 10506 5672
rect 10562 5616 10567 5672
rect 3601 5614 10567 5616
rect 3601 5611 3667 5614
rect 10501 5611 10567 5614
rect 12341 5674 12407 5677
rect 21173 5674 21239 5677
rect 23197 5674 23263 5677
rect 12341 5672 23263 5674
rect 12341 5616 12346 5672
rect 12402 5616 21178 5672
rect 21234 5616 23202 5672
rect 23258 5616 23263 5672
rect 12341 5614 23263 5616
rect 12341 5611 12407 5614
rect 21173 5611 21239 5614
rect 23197 5611 23263 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 21909 5266 21975 5269
rect 21909 5264 27722 5266
rect 21909 5208 21914 5264
rect 21970 5208 27722 5264
rect 21909 5206 27722 5208
rect 21909 5203 21975 5206
rect 10277 4928 10597 4929
rect 0 4768 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27662 4888 27722 5206
rect 19610 4863 19930 4864
rect 4061 4858 4127 4861
rect 9305 4858 9371 4861
rect 9857 4858 9923 4861
rect 4061 4856 9923 4858
rect 4061 4800 4066 4856
rect 4122 4800 9310 4856
rect 9366 4800 9862 4856
rect 9918 4800 9923 4856
rect 4061 4798 9923 4800
rect 4061 4795 4127 4798
rect 9305 4795 9371 4798
rect 9857 4795 9923 4798
rect 11605 4858 11671 4861
rect 19425 4858 19491 4861
rect 11605 4856 19491 4858
rect 11605 4800 11610 4856
rect 11666 4800 19430 4856
rect 19486 4800 19491 4856
rect 11605 4798 19491 4800
rect 11605 4795 11671 4798
rect 19425 4795 19491 4798
rect 27520 4768 28000 4888
rect 62 4586 122 4768
rect 17125 4722 17191 4725
rect 20805 4722 20871 4725
rect 17125 4720 20871 4722
rect 17125 4664 17130 4720
rect 17186 4664 20810 4720
rect 20866 4664 20871 4720
rect 17125 4662 20871 4664
rect 17125 4659 17191 4662
rect 20805 4659 20871 4662
rect 19701 4586 19767 4589
rect 62 4584 19767 4586
rect 62 4528 19706 4584
rect 19762 4528 19767 4584
rect 62 4526 19767 4528
rect 19701 4523 19767 4526
rect 9397 4450 9463 4453
rect 11881 4450 11947 4453
rect 9397 4448 11947 4450
rect 9397 4392 9402 4448
rect 9458 4392 11886 4448
rect 11942 4392 11947 4448
rect 9397 4390 11947 4392
rect 9397 4387 9463 4390
rect 11881 4387 11947 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 5993 4314 6059 4317
rect 9949 4314 10015 4317
rect 5993 4312 10015 4314
rect 5993 4256 5998 4312
rect 6054 4256 9954 4312
rect 10010 4256 10015 4312
rect 5993 4254 10015 4256
rect 5993 4251 6059 4254
rect 9949 4251 10015 4254
rect 15929 4178 15995 4181
rect 19241 4178 19307 4181
rect 20345 4178 20411 4181
rect 15929 4176 20411 4178
rect 15929 4120 15934 4176
rect 15990 4120 19246 4176
rect 19302 4120 20350 4176
rect 20406 4120 20411 4176
rect 15929 4118 20411 4120
rect 15929 4115 15995 4118
rect 19241 4115 19307 4118
rect 20345 4115 20411 4118
rect 1853 4042 1919 4045
rect 8845 4042 8911 4045
rect 1853 4040 8911 4042
rect 1853 3984 1858 4040
rect 1914 3984 8850 4040
rect 8906 3984 8911 4040
rect 1853 3982 8911 3984
rect 1853 3979 1919 3982
rect 8845 3979 8911 3982
rect 3325 3906 3391 3909
rect 6453 3906 6519 3909
rect 9489 3906 9555 3909
rect 3325 3904 4170 3906
rect 3325 3848 3330 3904
rect 3386 3848 4170 3904
rect 3325 3846 4170 3848
rect 3325 3843 3391 3846
rect 4110 3770 4170 3846
rect 6453 3904 9555 3906
rect 6453 3848 6458 3904
rect 6514 3848 9494 3904
rect 9550 3848 9555 3904
rect 6453 3846 9555 3848
rect 6453 3843 6519 3846
rect 9489 3843 9555 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 8937 3770 9003 3773
rect 4110 3768 9003 3770
rect 4110 3712 8942 3768
rect 8998 3712 9003 3768
rect 4110 3710 9003 3712
rect 8937 3707 9003 3710
rect 0 3496 480 3528
rect 0 3440 110 3496
rect 166 3440 480 3496
rect 0 3408 480 3440
rect 3877 3498 3943 3501
rect 11605 3498 11671 3501
rect 3877 3496 11671 3498
rect 3877 3440 3882 3496
rect 3938 3440 11610 3496
rect 11666 3440 11671 3496
rect 3877 3438 11671 3440
rect 3877 3435 3943 3438
rect 11605 3435 11671 3438
rect 13537 3498 13603 3501
rect 27520 3500 28000 3528
rect 13537 3496 27354 3498
rect 13537 3440 13542 3496
rect 13598 3440 27354 3496
rect 13537 3438 27354 3440
rect 13537 3435 13603 3438
rect 16481 3362 16547 3365
rect 22829 3362 22895 3365
rect 16481 3360 22895 3362
rect 16481 3304 16486 3360
rect 16542 3304 22834 3360
rect 22890 3304 22895 3360
rect 16481 3302 22895 3304
rect 16481 3299 16547 3302
rect 22829 3299 22895 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 27294 3226 27354 3438
rect 27520 3436 27660 3500
rect 27724 3436 28000 3500
rect 27520 3408 28000 3436
rect 27654 3226 27660 3228
rect 27294 3166 27660 3226
rect 27654 3164 27660 3166
rect 27724 3164 27730 3228
rect 8937 3090 9003 3093
rect 23105 3090 23171 3093
rect 8937 3088 23171 3090
rect 8937 3032 8942 3088
rect 8998 3032 23110 3088
rect 23166 3032 23171 3088
rect 8937 3030 23171 3032
rect 8937 3027 9003 3030
rect 23105 3027 23171 3030
rect 12985 2954 13051 2957
rect 24117 2954 24183 2957
rect 12985 2952 24183 2954
rect 12985 2896 12990 2952
rect 13046 2896 24122 2952
rect 24178 2896 24183 2952
rect 12985 2894 24183 2896
rect 12985 2891 13051 2894
rect 24117 2891 24183 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 54 2620 60 2684
rect 124 2682 130 2684
rect 1209 2682 1275 2685
rect 124 2680 1275 2682
rect 124 2624 1214 2680
rect 1270 2624 1275 2680
rect 124 2622 1275 2624
rect 124 2620 130 2622
rect 1209 2619 1275 2622
rect 10869 2682 10935 2685
rect 10869 2680 13830 2682
rect 10869 2624 10874 2680
rect 10930 2624 13830 2680
rect 10869 2622 13830 2624
rect 10869 2619 10935 2622
rect 3233 2546 3299 2549
rect 8753 2546 8819 2549
rect 3233 2544 8819 2546
rect 3233 2488 3238 2544
rect 3294 2488 8758 2544
rect 8814 2488 8819 2544
rect 3233 2486 8819 2488
rect 13770 2546 13830 2622
rect 21449 2546 21515 2549
rect 13770 2544 21515 2546
rect 13770 2488 21454 2544
rect 21510 2488 21515 2544
rect 13770 2486 21515 2488
rect 3233 2483 3299 2486
rect 8753 2483 8819 2486
rect 21449 2483 21515 2486
rect 18137 2410 18203 2413
rect 24117 2410 24183 2413
rect 18137 2408 24183 2410
rect 18137 2352 18142 2408
rect 18198 2352 24122 2408
rect 24178 2352 24183 2408
rect 18137 2350 24183 2352
rect 18137 2347 18203 2350
rect 24117 2347 24183 2350
rect 5610 2208 5930 2209
rect 0 2140 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 0 2076 60 2140
rect 124 2076 480 2140
rect 0 2048 480 2076
rect 27520 2136 28000 2168
rect 27520 2080 27710 2136
rect 27766 2080 28000 2136
rect 27520 2048 28000 2080
rect 3141 2002 3207 2005
rect 12709 2002 12775 2005
rect 3141 2000 12775 2002
rect 3141 1944 3146 2000
rect 3202 1944 12714 2000
rect 12770 1944 12775 2000
rect 3141 1942 12775 1944
rect 3141 1939 3207 1942
rect 12709 1939 12775 1942
rect 16481 2002 16547 2005
rect 24945 2002 25011 2005
rect 16481 2000 25011 2002
rect 16481 1944 16486 2000
rect 16542 1944 24950 2000
rect 25006 1944 25011 2000
rect 16481 1942 25011 1944
rect 16481 1939 16547 1942
rect 24945 1939 25011 1942
rect 1669 1866 1735 1869
rect 20161 1866 20227 1869
rect 1669 1864 20227 1866
rect 1669 1808 1674 1864
rect 1730 1808 20166 1864
rect 20222 1808 20227 1864
rect 1669 1806 20227 1808
rect 1669 1803 1735 1806
rect 20161 1803 20227 1806
rect 2129 1730 2195 1733
rect 13261 1730 13327 1733
rect 2129 1728 13327 1730
rect 2129 1672 2134 1728
rect 2190 1672 13266 1728
rect 13322 1672 13327 1728
rect 2129 1670 13327 1672
rect 2129 1667 2195 1670
rect 13261 1667 13327 1670
rect 14641 1730 14707 1733
rect 23749 1730 23815 1733
rect 14641 1728 23815 1730
rect 14641 1672 14646 1728
rect 14702 1672 23754 1728
rect 23810 1672 23815 1728
rect 14641 1670 23815 1672
rect 14641 1667 14707 1670
rect 23749 1667 23815 1670
rect 10685 1594 10751 1597
rect 23657 1594 23723 1597
rect 10685 1592 23723 1594
rect 10685 1536 10690 1592
rect 10746 1536 23662 1592
rect 23718 1536 23723 1592
rect 10685 1534 23723 1536
rect 10685 1531 10751 1534
rect 23657 1531 23723 1534
rect 11789 1458 11855 1461
rect 24025 1458 24091 1461
rect 11789 1456 24091 1458
rect 11789 1400 11794 1456
rect 11850 1400 24030 1456
rect 24086 1400 24091 1456
rect 11789 1398 24091 1400
rect 11789 1395 11855 1398
rect 24025 1395 24091 1398
rect 2037 1322 2103 1325
rect 62 1320 2103 1322
rect 62 1264 2042 1320
rect 2098 1264 2103 1320
rect 62 1262 2103 1264
rect 62 808 122 1262
rect 2037 1259 2103 1262
rect 0 688 480 808
rect 27520 776 28000 808
rect 27520 720 27618 776
rect 27674 720 28000 776
rect 27520 688 28000 720
rect 9949 98 10015 101
rect 19701 98 19767 101
rect 9949 96 19767 98
rect 9949 40 9954 96
rect 10010 40 19706 96
rect 19762 40 19767 96
rect 9949 38 19767 40
rect 9949 35 10015 38
rect 19701 35 19767 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 3004 23292 3068 23356
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 11100 22068 11164 22132
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 3372 17036 3436 17100
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 2452 13772 2516 13836
rect 3924 13636 3988 13700
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 3188 13228 3252 13292
rect 3924 13092 3988 13156
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 20116 11732 20180 11796
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 11100 9692 11164 9756
rect 3188 9284 3252 9348
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 60 9012 124 9076
rect 60 8740 124 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 3004 6972 3068 7036
rect 2452 6700 2516 6764
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 3372 6292 3436 6356
rect 20116 6292 20180 6356
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 27660 3436 27724 3500
rect 27660 3164 27724 3228
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 60 2620 124 2684
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 60 2076 124 2140
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 3003 23356 3069 23357
rect 3003 23292 3004 23356
rect 3068 23292 3069 23356
rect 3003 23291 3069 23292
rect 2451 13836 2517 13837
rect 2451 13772 2452 13836
rect 2516 13772 2517 13836
rect 2451 13771 2517 13772
rect 59 9076 125 9077
rect 59 9012 60 9076
rect 124 9012 125 9076
rect 59 9011 125 9012
rect 62 8805 122 9011
rect 59 8804 125 8805
rect 59 8740 60 8804
rect 124 8740 125 8804
rect 59 8739 125 8740
rect 2454 6765 2514 13771
rect 3006 7037 3066 23291
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 3371 17100 3437 17101
rect 3371 17036 3372 17100
rect 3436 17036 3437 17100
rect 3371 17035 3437 17036
rect 3187 13292 3253 13293
rect 3187 13228 3188 13292
rect 3252 13228 3253 13292
rect 3187 13227 3253 13228
rect 3190 9349 3250 13227
rect 3187 9348 3253 9349
rect 3187 9284 3188 9348
rect 3252 9284 3253 9348
rect 3187 9283 3253 9284
rect 3003 7036 3069 7037
rect 3003 6972 3004 7036
rect 3068 6972 3069 7036
rect 3003 6971 3069 6972
rect 2451 6764 2517 6765
rect 2451 6700 2452 6764
rect 2516 6700 2517 6764
rect 2451 6699 2517 6700
rect 3374 6357 3434 17035
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 3923 13700 3989 13701
rect 3923 13636 3924 13700
rect 3988 13636 3989 13700
rect 3923 13635 3989 13636
rect 3926 13157 3986 13635
rect 3923 13156 3989 13157
rect 3923 13092 3924 13156
rect 3988 13092 3989 13156
rect 3923 13091 3989 13092
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 3371 6356 3437 6357
rect 3371 6292 3372 6356
rect 3436 6292 3437 6356
rect 3371 6291 3437 6292
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 59 2684 125 2685
rect 59 2620 60 2684
rect 124 2620 125 2684
rect 59 2619 125 2620
rect 62 2141 122 2619
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 59 2140 125 2141
rect 59 2076 60 2140
rect 124 2076 125 2140
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 11099 22132 11165 22133
rect 11099 22068 11100 22132
rect 11164 22068 11165 22132
rect 11099 22067 11165 22068
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 11102 9757 11162 22067
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 11099 9756 11165 9757
rect 11099 9692 11100 9756
rect 11164 9692 11165 9756
rect 11099 9691 11165 9692
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 20115 11796 20181 11797
rect 20115 11732 20116 11796
rect 20180 11732 20181 11796
rect 20115 11731 20181 11732
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 20118 6357 20178 11731
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 20115 6356 20181 6357
rect 20115 6292 20116 6356
rect 20180 6292 20181 6356
rect 20115 6291 20181 6292
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 27659 3500 27725 3501
rect 27659 3436 27660 3500
rect 27724 3436 27725 3500
rect 27659 3435 27725 3436
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 27662 3229 27722 3435
rect 27659 3228 27725 3229
rect 27659 3164 27660 3228
rect 27724 3164 27725 3228
rect 27659 3163 27725 3164
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 59 2075 125 2076
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _090_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _172_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _183_
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__C
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_16
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_20
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_35
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_33
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_39
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_50 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_54 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6900 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _119_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_80
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_78
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_91
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _278_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__C
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_or4_4  _186_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _184_
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_141
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_152
timestamp 1586364061
transform 1 0 15088 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _175_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_161
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__277__A
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_198 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_200
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_205
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_228
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _276_
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__276__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _274_
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__274__A
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_270
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_274
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _118_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_51
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_1  _089_
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_58
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_62
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_65
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_75
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_79
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_or4_4  _174_
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__D
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_112
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use scs8hd_or2_4  _185_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__186__D
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_116
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _277_
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_1  _141_
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_195
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_219
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _182_
timestamp 1586364061
transform 1 0 23184 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 23000 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_236
timestamp 1586364061
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_249
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_253
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_266
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_nand2_4  _151_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__D
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_17
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_21
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _092_
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__197__B
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__197__C
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _140_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__B
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_126
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_130
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_148
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_164
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_223
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _273_
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__273__A
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_266
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_3_270 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _120_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__D
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_79
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _197_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _193_
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__224__C
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__B
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__278__A
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_160
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_171
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_179
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_183
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_195
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21068 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_235
timestamp 1586364061
transform 1 0 22724 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_245
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_249
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_252
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_262 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_or4_4  _093_
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__B
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_37
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_49
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_or4_4  _216_
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__A
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__224__B
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__C
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use scs8hd_buf_1  _176_
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_203
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 314 592
use scs8hd_buf_2  _275_
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__275__A
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_233
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_237
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_241
timestamp 1586364061
transform 1 0 23276 0 1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _272_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__272__A
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_5_270
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_inv_8  _138_
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__C
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _190_
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 866 592
use scs8hd_or4_4  _208_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__232__C
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__D
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__B
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4324 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_50
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_49
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_54
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_75
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__B
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_79
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _088_
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__224__D
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _224_
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _195_
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__D
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_109
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_113
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13708 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_129
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_133
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_150
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_165
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_167
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 18124 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_182
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_200
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _181_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_218
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22540 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_242
timestamp 1586364061
transform 1 0 23368 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_233
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_237
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _271_
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__271__A
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 25116 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_260
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_266
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_270
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_276
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__D
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _232_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 4140 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__232__D
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_42
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_61
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__B
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _196_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__B
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_113
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_6  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_197
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_209
timestamp 1586364061
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21344 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_233
timestamp 1586364061
transform 1 0 22540 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_237
timestamp 1586364061
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_250
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_8
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__190__B
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_29
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_33
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _225_
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_126
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_145
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_166
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_189
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_216
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_233
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_237
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_265
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _194_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_164
timestamp 1586364061
transform 1 0 16192 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_179
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 21804 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21620 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_221
timestamp 1586364061
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_236
timestamp 1586364061
transform 1 0 22816 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23552 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25116 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_264
timestamp 1586364061
transform 1 0 25392 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_8  _150_
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_14
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_18
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__B
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_81
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_85
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_102
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_144
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_148
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_167
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_188
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_192
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_254
timestamp 1586364061
transform 1 0 24472 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_265
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__189__B
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__C
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _191_
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__192__B
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_66
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_12_118
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_164
timestamp 1586364061
transform 1 0 16192 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_168
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_189
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_201
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_219
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 23368 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23184 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_234
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_238
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_255
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_262
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_1  _134_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_or4_4  _152_
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_or3_4  _085_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _189_
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_14
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _112_
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 866 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_49
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 590 592
use scs8hd_or3_4  _103_
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _192_
timestamp 1586364061
transform 1 0 6900 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__C
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _206_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_72
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_74
timestamp 1586364061
transform 1 0 7912 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__B
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_112
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _121_
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_6  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_158
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_171
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_189
timestamp 1586364061
transform 1 0 18492 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_185
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_187
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__B
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_191
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_209
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_216
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_218
timestamp 1586364061
transform 1 0 21160 0 -1 10336
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_237
timestamp 1586364061
transform 1 0 22908 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_254
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _270_
timestamp 1586364061
transform 1 0 25208 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_265
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_266
timestamp 1586364061
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__270__A
timestamp 1586364061
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_or3_4  _100_
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_21
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_25
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__B
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_68
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_85
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _116_
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_140
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _227_
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__B
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_158
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _228_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_203
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_207
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_223
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_260
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_265
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_273
timestamp 1586364061
transform 1 0 26220 0 1 10336
box -38 -48 406 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__B
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_or3_4  _097_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_or3_4  _109_
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__B
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _207_
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_6  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_6  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 590 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_128
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_16_173
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_195
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_212
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_229
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_233
timestamp 1586364061
transform 1 0 22540 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_236
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_240
timestamp 1586364061
transform 1 0 23184 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_250
timestamp 1586364061
transform 1 0 24104 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_254
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 406 592
use scs8hd_buf_1  _124_
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 314 592
use scs8hd_buf_1  _130_
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _106_
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_44
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__B
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_55
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__B
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_65
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_69
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_103
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _226_
timestamp 1586364061
transform 1 0 12512 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__B
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_133
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_137
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_169
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_177
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_189
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_224
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_228
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_235
timestamp 1586364061
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_239
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _265_
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__265__A
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_17_270
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__C
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _230_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _200_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _203_
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _204_
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_101
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_139
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_143
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_186
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_194
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_226
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_230
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_18_243
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_260
timestamp 1586364061
transform 1 0 25024 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_272
timestamp 1586364061
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__260__A
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_10
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _110_
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_14
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_25
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__201__B
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_51
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_58
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_84
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__B
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_131
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_184
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_197
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_201
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_205
timestamp 1586364061
transform 1 0 19964 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_210
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_206
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_225
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_229
timestamp 1586364061
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_219
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_229
timestamp 1586364061
transform 1 0 22172 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22908 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24472 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_252
timestamp 1586364061
transform 1 0 24288 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_256
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_246
timestamp 1586364061
transform 1 0 23736 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_267
timestamp 1586364061
transform 1 0 25668 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_257
timestamp 1586364061
transform 1 0 24748 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_269
timestamp 1586364061
transform 1 0 25852 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _199_
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__B
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_85
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_89
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__214__A
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__214__B
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_105
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_109
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_148
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_165
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_169
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_212
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_217
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_21_229
timestamp 1586364061
transform 1 0 22172 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_234
timestamp 1586364061
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_238
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__269__A
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_265
timestamp 1586364061
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_buf_2  _260_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _201_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_29
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _202_
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_60
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_79
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _205_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _214_
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__213__B
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_107
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_119
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_171
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_176
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_228
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_241
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_2  _269_
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_1  _188_
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_8
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__256__A
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__B
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_90
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_94
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _213_
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__215__A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__215__B
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_134
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_146
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_201
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_222
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_226
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23092 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_233
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_237
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_241
timestamp 1586364061
transform 1 0 23276 0 1 14688
box -38 -48 314 592
use scs8hd_conb_1  _248_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_248
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_252
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_259
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_263
timestamp 1586364061
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _256_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_11
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_18
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_51
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_78
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _229_
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _215_
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_24_140
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_148
timestamp 1586364061
transform 1 0 14720 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_6  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_183
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_200
timestamp 1586364061
transform 1 0 19504 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_226
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_230
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22632 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_237
timestamp 1586364061
transform 1 0 22908 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_248
timestamp 1586364061
transform 1 0 23920 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _259_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__259__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_25
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_44
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_67
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_84
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_87
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_91
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_106
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_116
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_25_141
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_225
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_239
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_buf_2  _268_
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__268__A
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_263
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_267
timestamp 1586364061
transform 1 0 25668 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_275
timestamp 1586364061
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _187_
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _258_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__258__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_8  FILLER_26_12
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _209_
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_23
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__221__B
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _210_
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__210__B
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_120
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__219__A
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__219__B
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_146
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_155
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_170
timestamp 1586364061
transform 1 0 16744 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_176
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_178
timestamp 1586364061
transform 1 0 17480 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__212__B
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_188
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_192
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_204
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_218
timestamp 1586364061
transform 1 0 21160 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_215
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_229
timestamp 1586364061
transform 1 0 22172 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_226
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_230
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_240
timestamp 1586364061
transform 1 0 23184 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_6  FILLER_27_234
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_242
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _246_
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _267_
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__267__A
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_262
timestamp 1586364061
transform 1 0 25208 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_275
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _198_
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_8  FILLER_28_12
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _243_
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__238__B
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_29
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__B
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_45
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_49
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__231__B
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_87
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_100
timestamp 1586364061
transform 1 0 10304 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _221_
timestamp 1586364061
transform 1 0 11960 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _219_
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_148
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16008 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_160
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_164
timestamp 1586364061
transform 1 0 16192 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_28_179
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _212_
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_183
timestamp 1586364061
transform 1 0 17940 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_196
timestamp 1586364061
transform 1 0 19136 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_208
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_8  FILLER_28_218
timestamp 1586364061
transform 1 0 21160 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_226
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23184 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_232
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_243
timestamp 1586364061
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_255
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_8
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _249_
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_19
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _238_
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 866 592
use scs8hd_decap_6  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 590 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use scs8hd_fill_1  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _231_
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__222__B
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _222_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _223_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _218_
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__218__A
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_149
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_153
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__B
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_204
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _250_
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_215
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 774 592
use scs8hd_conb_1  _251_
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_226
timestamp 1586364061
transform 1 0 21896 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_238
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__279__A
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_253
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_12
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 406 592
use scs8hd_conb_1  _245_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__237__B
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_29
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_35
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _235_
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__B
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_39
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_42
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_55
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_72
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_76
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_97
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_111
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__223__B
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_118
timestamp 1586364061
transform 1 0 11960 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_122
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__218__B
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_138
timestamp 1586364061
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_165
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _211_
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_169
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_182
timestamp 1586364061
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_204
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use scs8hd_conb_1  _242_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_212
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_218
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_230
timestamp 1586364061
transform 1 0 22264 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_242
timestamp 1586364061
transform 1 0 23368 0 -1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _279_
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_254
timestamp 1586364061
transform 1 0 24472 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_259
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _257_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__257__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _237_
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _234_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_31_102
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _217_
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__217__A
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_106
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_139
timestamp 1586364061
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_165
timestamp 1586364061
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_172
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_176
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_181
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_187
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_191
timestamp 1586364061
transform 1 0 18676 0 1 19040
box -38 -48 406 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 19872 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_198
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_202
timestamp 1586364061
transform 1 0 19688 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _241_
timestamp 1586364061
transform 1 0 20056 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_233
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_241
timestamp 1586364061
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use scs8hd_buf_2  _266_
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__266__A
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_259
timestamp 1586364061
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_263
timestamp 1586364061
transform 1 0 25300 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_275
timestamp 1586364061
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 774 592
use scs8hd_nor2_4  _236_
timestamp 1586364061
transform 1 0 4784 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__234__B
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_49
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_32_53
timestamp 1586364061
transform 1 0 5980 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_115
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_151
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_171
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_188
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19136 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_199
timestamp 1586364061
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_211
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_9
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_13
timestamp 1586364061
transform 1 0 2300 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_17
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_21
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_25
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  _164_
timestamp 1586364061
transform 1 0 4416 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_32
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _239_
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__B
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_40
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_39
timestamp 1586364061
transform 1 0 4692 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_43
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_50
timestamp 1586364061
transform 1 0 5704 0 -1 21216
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_69
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_73
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_77
timestamp 1586364061
transform 1 0 8188 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_94
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_90
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_100
timestamp 1586364061
transform 1 0 10304 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_97
timestamp 1586364061
transform 1 0 10028 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_107
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_110
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _220_
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__220__B
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_127
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_118
timestamp 1586364061
transform 1 0 11960 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_128
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_134
timestamp 1586364061
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_158
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_162
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17388 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_169
timestamp 1586364061
transform 1 0 16652 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_173
timestamp 1586364061
transform 1 0 17020 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_187
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_191
timestamp 1586364061
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_186
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_198
timestamp 1586364061
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_198
timestamp 1586364061
transform 1 0 19320 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_210
timestamp 1586364061
transform 1 0 20424 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_226
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_238
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _255_
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__255__A
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_11
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_23
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_40
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_79
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_96
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_35_115
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_119
timestamp 1586364061
transform 1 0 12052 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_139
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_152
timestamp 1586364061
transform 1 0 15088 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_169
timestamp 1586364061
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_173
timestamp 1586364061
transform 1 0 17020 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_177
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_191
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_203
timestamp 1586364061
transform 1 0 19780 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_215
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_227
timestamp 1586364061
transform 1 0 21988 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_35_239
timestamp 1586364061
transform 1 0 23092 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_243
timestamp 1586364061
transform 1 0 23460 0 1 21216
box -38 -48 130 592
use scs8hd_buf_2  _264_
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__264__A
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_259
timestamp 1586364061
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_263
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_275
timestamp 1586364061
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__252__A
timestamp 1586364061
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_7
timestamp 1586364061
transform 1 0 1748 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_19
timestamp 1586364061
transform 1 0 2852 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_conb_1  _240_
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_47
timestamp 1586364061
transform 1 0 5428 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6164 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_58
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_75
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_85
timestamp 1586364061
transform 1 0 8924 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_90
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_109
timestamp 1586364061
transform 1 0 11132 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_116
timestamp 1586364061
transform 1 0 11776 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_124
timestamp 1586364061
transform 1 0 12512 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_128
timestamp 1586364061
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_36_139
timestamp 1586364061
transform 1 0 13892 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_6  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 22304
box -38 -48 866 592
use scs8hd_fill_1  FILLER_36_160
timestamp 1586364061
transform 1 0 15824 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_170
timestamp 1586364061
transform 1 0 16744 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_182
timestamp 1586364061
transform 1 0 17848 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_194
timestamp 1586364061
transform 1 0 18952 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_206
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _254_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__254__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_23
timestamp 1586364061
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_35
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_47
timestamp 1586364061
transform 1 0 5428 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_76
timestamp 1586364061
transform 1 0 8096 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_83
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_97
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_101
timestamp 1586364061
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_112
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _153_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_116
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_137
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_141
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_148
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_152
timestamp 1586364061
transform 1 0 15088 0 1 22304
box -38 -48 406 592
use scs8hd_conb_1  _247_
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_161
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_169
timestamp 1586364061
transform 1 0 16652 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__261__A
timestamp 1586364061
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_200
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_212
timestamp 1586364061
transform 1 0 20608 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_224
timestamp 1586364061
transform 1 0 21712 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__263__A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_buf_2  _252_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_70
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_74
timestamp 1586364061
transform 1 0 7912 0 -1 23392
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_113
timestamp 1586364061
transform 1 0 11500 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_124
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_132
timestamp 1586364061
transform 1 0 13248 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_138
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_150
timestamp 1586364061
transform 1 0 14904 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_159
timestamp 1586364061
transform 1 0 15732 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_167
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_173
timestamp 1586364061
transform 1 0 17020 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _261_
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_38_181
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_188
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_200
timestamp 1586364061
transform 1 0 19504 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_212
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _263_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_buf_2  _253_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__253__A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_35
timestamp 1586364061
transform 1 0 4324 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_47
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_1  _233_
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_88
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_conb_1  _244_
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_92
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_99
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_101
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10580 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_106
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_116
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_126
timestamp 1586364061
transform 1 0 12696 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_130
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _287_
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__287__A
timestamp 1586364061
transform 1 0 14904 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_148
timestamp 1586364061
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_152
timestamp 1586364061
transform 1 0 15088 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _286_
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_160
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 590 592
use scs8hd_buf_2  _285_
timestamp 1586364061
transform 1 0 16928 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__286__A
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__285__A
timestamp 1586364061
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_174
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 590 592
use scs8hd_decap_8  FILLER_40_176
timestamp 1586364061
transform 1 0 17296 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _280_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _284_
timestamp 1586364061
transform 1 0 18032 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__284__A
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__280__A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_180
timestamp 1586364061
transform 1 0 17664 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_188
timestamp 1586364061
transform 1 0 18400 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_200
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _283_
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__283__A
timestamp 1586364061
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_211
timestamp 1586364061
transform 1 0 20516 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_215
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_212
timestamp 1586364061
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _281_
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _282_
timestamp 1586364061
transform 1 0 21252 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__282__A
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__281__A
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _262_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__262__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 3330 0 3386 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 4250 0 4306 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 5262 0 5318 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 6182 0 6238 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 7194 0 7250 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 8114 0 8170 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 9126 0 9182 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 478 0 534 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal3 s 0 2048 480 2168 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 0 3408 480 3528 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 0 21632 480 21752 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal3 s 0 24488 480 24608 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal3 s 0 27208 480 27328 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 27520 2048 28000 2168 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 27520 3408 28000 3528 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 27520 6264 28000 6384 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 27520 13200 28000 13320 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 27520 16056 28000 16176 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 27520 18776 28000 18896 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 27520 21632 28000 21752 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 27520 24488 28000 24608 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 27520 27208 28000 27328 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal2 s 16854 0 16910 480 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal2 s 21638 0 21694 480 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal2 s 23570 0 23626 480 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal2 s 24582 0 24638 480 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal2 s 27434 0 27490 480 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal2 s 662 27520 718 28000 6 chany_top_in[0]
port 63 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 chany_top_in[1]
port 64 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 chany_top_in[2]
port 65 nsew default input
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[3]
port 66 nsew default input
rlabel metal2 s 6182 27520 6238 28000 6 chany_top_in[4]
port 67 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 68 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[6]
port 69 nsew default input
rlabel metal2 s 10414 27520 10470 28000 6 chany_top_in[7]
port 70 nsew default input
rlabel metal2 s 11794 27520 11850 28000 6 chany_top_in[8]
port 71 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_out[0]
port 72 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 18786 27520 18842 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 20166 27520 20222 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 21638 27520 21694 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 24398 27520 24454 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 25778 27520 25834 28000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 27158 27520 27214 28000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 10046 0 10102 480 6 data_in
port 81 nsew default input
rlabel metal2 s 2318 0 2374 480 6 enable
port 82 nsew default input
rlabel metal3 s 0 14696 480 14816 6 left_bottom_grid_pin_12_
port 83 nsew default input
rlabel metal3 s 0 688 480 808 6 left_top_grid_pin_10_
port 84 nsew default input
rlabel metal3 s 27520 14696 28000 14816 6 right_bottom_grid_pin_12_
port 85 nsew default input
rlabel metal3 s 27520 688 28000 808 6 right_top_grid_pin_10_
port 86 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 top_left_grid_pin_13_
port 87 nsew default input
rlabel metal2 s 14646 27520 14702 28000 6 top_right_grid_pin_11_
port 88 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 89 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 90 nsew default input
<< end >>
