magic
tech sky130A
magscale 1 2
timestamp 1608762952
<< checkpaint >>
rect -1260 -1260 24060 24060
<< locali >>
rect 9505 19703 9539 20009
rect 9597 19771 9631 19941
rect 10885 19771 10919 19941
rect 7389 18275 7423 18377
rect 13277 18139 13311 18377
rect 18061 18139 18095 18377
rect 18981 18071 19015 18377
rect 19257 18207 19291 18377
rect 9505 16983 9539 17085
rect 17233 14807 17267 15113
rect 13645 14331 13679 14569
rect 9505 13345 9597 13379
rect 9505 13175 9539 13345
rect 13737 12767 13771 12937
rect 5549 12087 5583 12393
rect 6377 11543 6411 11849
rect 7757 11543 7791 11713
rect 6377 10999 6411 11305
rect 6469 10999 6503 11237
rect 7389 11135 7423 11305
rect 8401 10523 8435 10693
rect 5457 9367 5491 9469
rect 12265 7803 12299 7973
rect 4629 7327 4663 7497
rect 5273 6783 5307 6953
rect 7205 6647 7239 6817
rect 7147 6613 7239 6647
rect 9689 6307 9723 6409
<< viali >>
rect 1685 20009 1719 20043
rect 5273 20009 5307 20043
rect 5733 20009 5767 20043
rect 6285 20009 6319 20043
rect 8401 20009 8435 20043
rect 9321 20009 9355 20043
rect 9505 20009 9539 20043
rect 13461 20009 13495 20043
rect 14013 20009 14047 20043
rect 15117 20009 15151 20043
rect 15669 20009 15703 20043
rect 16313 20009 16347 20043
rect 17417 20009 17451 20043
rect 18521 20009 18555 20043
rect 20085 20009 20119 20043
rect 4537 19941 4571 19975
rect 1501 19873 1535 19907
rect 2053 19873 2087 19907
rect 4445 19873 4479 19907
rect 5089 19873 5123 19907
rect 5641 19873 5675 19907
rect 2237 19805 2271 19839
rect 4721 19805 4755 19839
rect 5917 19805 5951 19839
rect 3433 19737 3467 19771
rect 3893 19737 3927 19771
rect 9597 19941 9631 19975
rect 10885 19941 10919 19975
rect 11713 19941 11747 19975
rect 20821 19941 20855 19975
rect 9781 19805 9815 19839
rect 13277 19873 13311 19907
rect 13829 19873 13863 19907
rect 16129 19873 16163 19907
rect 17233 19873 17267 19907
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 11069 19805 11103 19839
rect 14749 19805 14783 19839
rect 9597 19737 9631 19771
rect 10609 19737 10643 19771
rect 10885 19737 10919 19771
rect 17785 19737 17819 19771
rect 19073 19737 19107 19771
rect 2881 19669 2915 19703
rect 4077 19669 4111 19703
rect 6745 19669 6779 19703
rect 7113 19669 7147 19703
rect 7481 19669 7515 19703
rect 8033 19669 8067 19703
rect 8769 19669 8803 19703
rect 9505 19669 9539 19703
rect 10241 19669 10275 19703
rect 11345 19669 11379 19703
rect 12081 19669 12115 19703
rect 12817 19669 12851 19703
rect 14381 19669 14415 19703
rect 16681 19669 16715 19703
rect 17049 19669 17083 19703
rect 19809 19669 19843 19703
rect 20453 19669 20487 19703
rect 8401 19329 8435 19363
rect 8585 19329 8619 19363
rect 9413 19329 9447 19363
rect 9597 19329 9631 19363
rect 9965 19329 9999 19363
rect 12817 19329 12851 19363
rect 17233 19329 17267 19363
rect 1501 19261 1535 19295
rect 2053 19261 2087 19295
rect 3065 19261 3099 19295
rect 5089 19261 5123 19295
rect 7849 19261 7883 19295
rect 11621 19261 11655 19295
rect 12909 19261 12943 19295
rect 13645 19261 13679 19295
rect 14197 19261 14231 19295
rect 14749 19261 14783 19295
rect 15301 19261 15335 19295
rect 15853 19261 15887 19295
rect 16405 19261 16439 19295
rect 16957 19261 16991 19295
rect 18061 19261 18095 19295
rect 18797 19261 18831 19295
rect 19809 19261 19843 19295
rect 2329 19193 2363 19227
rect 3332 19193 3366 19227
rect 5356 19193 5390 19227
rect 7389 19193 7423 19227
rect 9321 19193 9355 19227
rect 10210 19193 10244 19227
rect 11897 19193 11931 19227
rect 13185 19193 13219 19227
rect 18337 19193 18371 19227
rect 19349 19193 19383 19227
rect 20453 19193 20487 19227
rect 1685 19125 1719 19159
rect 2789 19125 2823 19159
rect 4445 19125 4479 19159
rect 4905 19125 4939 19159
rect 6469 19125 6503 19159
rect 7021 19125 7055 19159
rect 7941 19125 7975 19159
rect 8309 19125 8343 19159
rect 8953 19125 8987 19159
rect 11345 19125 11379 19159
rect 13829 19125 13863 19159
rect 14381 19125 14415 19159
rect 14933 19125 14967 19159
rect 15485 19125 15519 19159
rect 16037 19125 16071 19159
rect 16589 19125 16623 19159
rect 17693 19125 17727 19159
rect 18981 19125 19015 19159
rect 20913 19125 20947 19159
rect 1593 18921 1627 18955
rect 2881 18921 2915 18955
rect 4537 18921 4571 18955
rect 6745 18921 6779 18955
rect 19533 18921 19567 18955
rect 2237 18853 2271 18887
rect 9321 18853 9355 18887
rect 10118 18853 10152 18887
rect 11529 18853 11563 18887
rect 12081 18853 12115 18887
rect 13553 18853 13587 18887
rect 15577 18853 15611 18887
rect 20269 18853 20303 18887
rect 1409 18785 1443 18819
rect 1961 18785 1995 18819
rect 3249 18785 3283 18819
rect 3341 18785 3375 18819
rect 4445 18785 4479 18819
rect 5632 18785 5666 18819
rect 7829 18785 7863 18819
rect 11805 18785 11839 18819
rect 12541 18785 12575 18819
rect 13277 18785 13311 18819
rect 15301 18785 15335 18819
rect 16037 18785 16071 18819
rect 16773 18785 16807 18819
rect 17693 18785 17727 18819
rect 17969 18785 18003 18819
rect 18429 18785 18463 18819
rect 20637 18785 20671 18819
rect 3525 18717 3559 18751
rect 4721 18717 4755 18751
rect 5365 18717 5399 18751
rect 7113 18717 7147 18751
rect 7573 18717 7607 18751
rect 9873 18717 9907 18751
rect 12817 18717 12851 18751
rect 16313 18717 16347 18751
rect 17049 18717 17083 18751
rect 18705 18717 18739 18751
rect 19165 18717 19199 18751
rect 4077 18649 4111 18683
rect 2789 18581 2823 18615
rect 5273 18581 5307 18615
rect 8953 18581 8987 18615
rect 11253 18581 11287 18615
rect 14013 18581 14047 18615
rect 14473 18581 14507 18615
rect 15117 18581 15151 18615
rect 17509 18581 17543 18615
rect 19901 18581 19935 18615
rect 21097 18581 21131 18615
rect 2605 18377 2639 18411
rect 4077 18377 4111 18411
rect 4997 18377 5031 18411
rect 5549 18377 5583 18411
rect 7389 18377 7423 18411
rect 7573 18377 7607 18411
rect 11161 18377 11195 18411
rect 12449 18377 12483 18411
rect 13277 18377 13311 18411
rect 14841 18377 14875 18411
rect 18061 18377 18095 18411
rect 18337 18377 18371 18411
rect 18981 18377 19015 18411
rect 5365 18309 5399 18343
rect 8769 18309 8803 18343
rect 4445 18241 4479 18275
rect 6193 18241 6227 18275
rect 7389 18241 7423 18275
rect 8217 18241 8251 18275
rect 9321 18241 9355 18275
rect 12173 18241 12207 18275
rect 12909 18241 12943 18275
rect 13093 18241 13127 18275
rect 1777 18173 1811 18207
rect 2697 18173 2731 18207
rect 6009 18173 6043 18207
rect 6837 18173 6871 18207
rect 8585 18173 8619 18207
rect 9137 18173 9171 18207
rect 9781 18173 9815 18207
rect 14013 18241 14047 18275
rect 15485 18241 15519 18275
rect 15669 18241 15703 18275
rect 16681 18241 16715 18275
rect 17141 18173 17175 18207
rect 18705 18309 18739 18343
rect 18153 18173 18187 18207
rect 1685 18105 1719 18139
rect 2964 18105 2998 18139
rect 6561 18105 6595 18139
rect 7113 18105 7147 18139
rect 7941 18105 7975 18139
rect 8033 18105 8067 18139
rect 9229 18105 9263 18139
rect 10048 18105 10082 18139
rect 11897 18105 11931 18139
rect 13277 18105 13311 18139
rect 13829 18105 13863 18139
rect 16497 18105 16531 18139
rect 17417 18105 17451 18139
rect 18061 18105 18095 18139
rect 19257 18377 19291 18411
rect 19441 18377 19475 18411
rect 20545 18309 20579 18343
rect 21005 18241 21039 18275
rect 19073 18173 19107 18207
rect 19257 18173 19291 18207
rect 1961 18037 1995 18071
rect 5917 18037 5951 18071
rect 11437 18037 11471 18071
rect 12817 18037 12851 18071
rect 13461 18037 13495 18071
rect 13921 18037 13955 18071
rect 14473 18037 14507 18071
rect 15025 18037 15059 18071
rect 15393 18037 15427 18071
rect 16037 18037 16071 18071
rect 16405 18037 16439 18071
rect 18981 18037 19015 18071
rect 19809 18037 19843 18071
rect 20177 18037 20211 18071
rect 2513 17833 2547 17867
rect 3433 17833 3467 17867
rect 4261 17833 4295 17867
rect 7665 17833 7699 17867
rect 8033 17833 8067 17867
rect 8401 17833 8435 17867
rect 9229 17833 9263 17867
rect 10149 17833 10183 17867
rect 10701 17833 10735 17867
rect 13645 17833 13679 17867
rect 14197 17833 14231 17867
rect 21097 17833 21131 17867
rect 5540 17765 5574 17799
rect 17877 17765 17911 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 2881 17697 2915 17731
rect 7297 17697 7331 17731
rect 8493 17697 8527 17731
rect 10057 17697 10091 17731
rect 12245 17697 12279 17731
rect 14565 17697 14599 17731
rect 14657 17697 14691 17731
rect 15568 17697 15602 17731
rect 17785 17697 17819 17731
rect 18429 17697 18463 17731
rect 20361 17697 20395 17731
rect 4813 17629 4847 17663
rect 5273 17629 5307 17663
rect 8769 17629 8803 17663
rect 10333 17629 10367 17663
rect 11989 17629 12023 17663
rect 14841 17629 14875 17663
rect 15301 17629 15335 17663
rect 16957 17629 16991 17663
rect 17969 17629 18003 17663
rect 18889 17629 18923 17663
rect 3065 17561 3099 17595
rect 9689 17561 9723 17595
rect 13369 17561 13403 17595
rect 17417 17561 17451 17595
rect 19993 17561 20027 17595
rect 1685 17493 1719 17527
rect 1961 17493 1995 17527
rect 4721 17493 4755 17527
rect 6653 17493 6687 17527
rect 11161 17493 11195 17527
rect 11437 17493 11471 17527
rect 11897 17493 11931 17527
rect 16681 17493 16715 17527
rect 19257 17493 19291 17527
rect 19625 17493 19659 17527
rect 2881 17289 2915 17323
rect 10977 17289 11011 17323
rect 11897 17289 11931 17323
rect 20453 17289 20487 17323
rect 4721 17221 4755 17255
rect 14105 17221 14139 17255
rect 16037 17221 16071 17255
rect 16497 17221 16531 17255
rect 16957 17221 16991 17255
rect 2329 17153 2363 17187
rect 2973 17153 3007 17187
rect 5089 17153 5123 17187
rect 5825 17153 5859 17187
rect 9597 17153 9631 17187
rect 11253 17153 11287 17187
rect 12265 17153 12299 17187
rect 17417 17153 17451 17187
rect 17601 17153 17635 17187
rect 18061 17153 18095 17187
rect 21189 17153 21223 17187
rect 1501 17085 1535 17119
rect 2053 17085 2087 17119
rect 3240 17085 3274 17119
rect 5549 17085 5583 17119
rect 6193 17085 6227 17119
rect 7297 17085 7331 17119
rect 7564 17085 7598 17119
rect 9505 17085 9539 17119
rect 9864 17085 9898 17119
rect 12725 17085 12759 17119
rect 12992 17085 13026 17119
rect 14657 17085 14691 17119
rect 20085 17085 20119 17119
rect 9045 17017 9079 17051
rect 14902 17017 14936 17051
rect 18306 17017 18340 17051
rect 19717 17017 19751 17051
rect 1685 16949 1719 16983
rect 4353 16949 4387 16983
rect 5181 16949 5215 16983
rect 5641 16949 5675 16983
rect 6561 16949 6595 16983
rect 7205 16949 7239 16983
rect 8677 16949 8711 16983
rect 9137 16949 9171 16983
rect 9505 16949 9539 16983
rect 14565 16949 14599 16983
rect 16773 16949 16807 16983
rect 17325 16949 17359 16983
rect 19441 16949 19475 16983
rect 20821 16949 20855 16983
rect 1777 16745 1811 16779
rect 4537 16745 4571 16779
rect 7849 16745 7883 16779
rect 7941 16745 7975 16779
rect 9413 16745 9447 16779
rect 10057 16745 10091 16779
rect 10149 16745 10183 16779
rect 11069 16745 11103 16779
rect 11437 16745 11471 16779
rect 11897 16745 11931 16779
rect 12909 16745 12943 16779
rect 13461 16745 13495 16779
rect 13829 16745 13863 16779
rect 13921 16745 13955 16779
rect 15669 16745 15703 16779
rect 16313 16745 16347 16779
rect 17785 16745 17819 16779
rect 19441 16745 19475 16779
rect 20453 16745 20487 16779
rect 21097 16745 21131 16779
rect 19717 16677 19751 16711
rect 1593 16609 1627 16643
rect 2145 16609 2179 16643
rect 3249 16609 3283 16643
rect 3341 16609 3375 16643
rect 4445 16609 4479 16643
rect 5181 16609 5215 16643
rect 5917 16609 5951 16643
rect 6377 16609 6411 16643
rect 6653 16609 6687 16643
rect 8677 16609 8711 16643
rect 11805 16609 11839 16643
rect 12817 16609 12851 16643
rect 14473 16609 14507 16643
rect 16672 16609 16706 16643
rect 18328 16609 18362 16643
rect 20085 16609 20119 16643
rect 2421 16541 2455 16575
rect 3525 16541 3559 16575
rect 4629 16541 4663 16575
rect 5273 16541 5307 16575
rect 7389 16541 7423 16575
rect 8125 16541 8159 16575
rect 10333 16541 10367 16575
rect 11989 16541 12023 16575
rect 13093 16541 13127 16575
rect 14105 16541 14139 16575
rect 16412 16541 16446 16575
rect 18061 16541 18095 16575
rect 12449 16473 12483 16507
rect 2881 16405 2915 16439
rect 4077 16405 4111 16439
rect 5733 16405 5767 16439
rect 6193 16405 6227 16439
rect 7481 16405 7515 16439
rect 8493 16405 8527 16439
rect 9137 16405 9171 16439
rect 9689 16405 9723 16439
rect 10701 16405 10735 16439
rect 14933 16405 14967 16439
rect 1593 16201 1627 16235
rect 4077 16201 4111 16235
rect 4537 16201 4571 16235
rect 6285 16201 6319 16235
rect 8769 16201 8803 16235
rect 10333 16201 10367 16235
rect 12081 16201 12115 16235
rect 17877 16201 17911 16235
rect 18061 16201 18095 16235
rect 19441 16201 19475 16235
rect 14933 16133 14967 16167
rect 15945 16133 15979 16167
rect 20545 16133 20579 16167
rect 2145 16065 2179 16099
rect 6653 16065 6687 16099
rect 12633 16065 12667 16099
rect 18705 16065 18739 16099
rect 1409 15997 1443 16031
rect 1961 15997 1995 16031
rect 2697 15997 2731 16031
rect 2964 15997 2998 16031
rect 4905 15997 4939 16031
rect 7113 15997 7147 16031
rect 7380 15997 7414 16031
rect 8953 15997 8987 16031
rect 10701 15997 10735 16031
rect 10968 15997 11002 16031
rect 13277 15997 13311 16031
rect 15117 15997 15151 16031
rect 16129 15997 16163 16031
rect 18521 15997 18555 16031
rect 20913 15997 20947 16031
rect 5172 15929 5206 15963
rect 9198 15929 9232 15963
rect 13544 15929 13578 15963
rect 18429 15929 18463 15963
rect 19073 15929 19107 15963
rect 19809 15929 19843 15963
rect 8493 15861 8527 15895
rect 12817 15861 12851 15895
rect 14657 15861 14691 15895
rect 15393 15861 15427 15895
rect 15761 15861 15795 15895
rect 16405 15861 16439 15895
rect 16865 15861 16899 15895
rect 17141 15861 17175 15895
rect 20177 15861 20211 15895
rect 2053 15657 2087 15691
rect 2421 15657 2455 15691
rect 3249 15657 3283 15691
rect 3709 15657 3743 15691
rect 4997 15657 5031 15691
rect 6101 15657 6135 15691
rect 6929 15657 6963 15691
rect 9045 15657 9079 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 12909 15657 12943 15691
rect 13921 15657 13955 15691
rect 15853 15657 15887 15691
rect 16221 15657 16255 15691
rect 16865 15657 16899 15691
rect 17877 15657 17911 15691
rect 18889 15657 18923 15691
rect 19441 15657 19475 15691
rect 20085 15657 20119 15691
rect 14013 15589 14047 15623
rect 14933 15589 14967 15623
rect 20453 15589 20487 15623
rect 2789 15521 2823 15555
rect 3157 15521 3191 15555
rect 4537 15521 4571 15555
rect 6009 15521 6043 15555
rect 6653 15521 6687 15555
rect 7297 15521 7331 15555
rect 7941 15521 7975 15555
rect 8953 15521 8987 15555
rect 10057 15521 10091 15555
rect 11060 15521 11094 15555
rect 15485 15521 15519 15555
rect 18245 15521 18279 15555
rect 21097 15521 21131 15555
rect 5089 15453 5123 15487
rect 5273 15453 5307 15487
rect 6285 15453 6319 15487
rect 7389 15453 7423 15487
rect 7481 15453 7515 15487
rect 9137 15453 9171 15487
rect 10241 15453 10275 15487
rect 10793 15453 10827 15487
rect 13001 15453 13035 15487
rect 13185 15453 13219 15487
rect 14197 15453 14231 15487
rect 16313 15453 16347 15487
rect 16497 15453 16531 15487
rect 18337 15453 18371 15487
rect 18521 15453 18555 15487
rect 8585 15385 8619 15419
rect 14565 15385 14599 15419
rect 19717 15385 19751 15419
rect 1593 15317 1627 15351
rect 4629 15317 4663 15351
rect 5641 15317 5675 15351
rect 8401 15317 8435 15351
rect 12173 15317 12207 15351
rect 12541 15317 12575 15351
rect 13553 15317 13587 15351
rect 17417 15317 17451 15351
rect 17785 15317 17819 15351
rect 4721 15113 4755 15147
rect 6193 15113 6227 15147
rect 6561 15113 6595 15147
rect 7941 15113 7975 15147
rect 8585 15113 8619 15147
rect 10333 15113 10367 15147
rect 10701 15113 10735 15147
rect 11161 15113 11195 15147
rect 14013 15113 14047 15147
rect 17141 15113 17175 15147
rect 17233 15113 17267 15147
rect 20269 15113 20303 15147
rect 1593 15045 1627 15079
rect 7113 15045 7147 15079
rect 2237 14977 2271 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 13185 14977 13219 15011
rect 14841 14977 14875 15011
rect 15025 14977 15059 15011
rect 15761 14977 15795 15011
rect 1409 14909 1443 14943
rect 1961 14909 1995 14943
rect 2881 14909 2915 14943
rect 3148 14909 3182 14943
rect 4813 14909 4847 14943
rect 5080 14909 5114 14943
rect 7297 14909 7331 14943
rect 8677 14909 8711 14943
rect 13001 14909 13035 14943
rect 13093 14909 13127 14943
rect 14197 14909 14231 14943
rect 14749 14909 14783 14943
rect 15393 14909 15427 14943
rect 2697 14841 2731 14875
rect 8922 14841 8956 14875
rect 16028 14841 16062 14875
rect 19625 15045 19659 15079
rect 17417 14977 17451 15011
rect 19901 14977 19935 15011
rect 18245 14909 18279 14943
rect 18512 14909 18546 14943
rect 21005 14909 21039 14943
rect 17785 14841 17819 14875
rect 20637 14841 20671 14875
rect 4261 14773 4295 14807
rect 7573 14773 7607 14807
rect 10057 14773 10091 14807
rect 11345 14773 11379 14807
rect 11713 14773 11747 14807
rect 12633 14773 12667 14807
rect 13645 14773 13679 14807
rect 14381 14773 14415 14807
rect 17233 14773 17267 14807
rect 1593 14569 1627 14603
rect 4537 14569 4571 14603
rect 5089 14569 5123 14603
rect 6561 14569 6595 14603
rect 9045 14569 9079 14603
rect 10149 14569 10183 14603
rect 10609 14569 10643 14603
rect 13185 14569 13219 14603
rect 13645 14569 13679 14603
rect 15945 14569 15979 14603
rect 16589 14569 16623 14603
rect 21097 14569 21131 14603
rect 8401 14501 8435 14535
rect 1409 14433 1443 14467
rect 1961 14433 1995 14467
rect 3341 14433 3375 14467
rect 3433 14433 3467 14467
rect 4445 14433 4479 14467
rect 6920 14433 6954 14467
rect 11253 14433 11287 14467
rect 11805 14433 11839 14467
rect 2145 14365 2179 14399
rect 3525 14365 3559 14399
rect 4629 14365 4663 14399
rect 6653 14365 6687 14399
rect 10977 14365 11011 14399
rect 11897 14365 11931 14399
rect 12081 14365 12115 14399
rect 12449 14365 12483 14399
rect 13277 14365 13311 14399
rect 13461 14365 13495 14399
rect 14197 14501 14231 14535
rect 18337 14501 18371 14535
rect 18696 14501 18730 14535
rect 20453 14501 20487 14535
rect 16037 14433 16071 14467
rect 16957 14433 16991 14467
rect 20085 14433 20119 14467
rect 14289 14365 14323 14399
rect 14473 14365 14507 14399
rect 16221 14365 16255 14399
rect 17049 14365 17083 14399
rect 17233 14365 17267 14399
rect 17601 14365 17635 14399
rect 18429 14365 18463 14399
rect 2973 14297 3007 14331
rect 5825 14297 5859 14331
rect 11437 14297 11471 14331
rect 12817 14297 12851 14331
rect 13645 14297 13679 14331
rect 15577 14297 15611 14331
rect 2881 14229 2915 14263
rect 4077 14229 4111 14263
rect 6101 14229 6135 14263
rect 8033 14229 8067 14263
rect 8677 14229 8711 14263
rect 13829 14229 13863 14263
rect 14841 14229 14875 14263
rect 19809 14229 19843 14263
rect 1777 14025 1811 14059
rect 3157 14025 3191 14059
rect 3801 14025 3835 14059
rect 5733 14025 5767 14059
rect 9781 14025 9815 14059
rect 10425 14025 10459 14059
rect 20177 14025 20211 14059
rect 5273 13957 5307 13991
rect 5641 13957 5675 13991
rect 6837 13957 6871 13991
rect 15945 13957 15979 13991
rect 19441 13957 19475 13991
rect 19809 13957 19843 13991
rect 2329 13889 2363 13923
rect 3249 13889 3283 13923
rect 6285 13889 6319 13923
rect 7389 13889 7423 13923
rect 13461 13889 13495 13923
rect 13645 13889 13679 13923
rect 18705 13889 18739 13923
rect 20545 13889 20579 13923
rect 1593 13821 1627 13855
rect 2145 13821 2179 13855
rect 3893 13821 3927 13855
rect 4160 13821 4194 13855
rect 6193 13821 6227 13855
rect 7205 13821 7239 13855
rect 8401 13821 8435 13855
rect 8668 13821 8702 13855
rect 10609 13821 10643 13855
rect 10876 13821 10910 13855
rect 14013 13821 14047 13855
rect 16313 13821 16347 13855
rect 16580 13821 16614 13855
rect 18429 13821 18463 13855
rect 19073 13821 19107 13855
rect 20913 13821 20947 13855
rect 6101 13753 6135 13787
rect 7849 13753 7883 13787
rect 14280 13753 14314 13787
rect 18521 13753 18555 13787
rect 7297 13685 7331 13719
rect 10057 13685 10091 13719
rect 11989 13685 12023 13719
rect 12909 13685 12943 13719
rect 13001 13685 13035 13719
rect 13369 13685 13403 13719
rect 15393 13685 15427 13719
rect 17693 13685 17727 13719
rect 18061 13685 18095 13719
rect 2789 13481 2823 13515
rect 4445 13481 4479 13515
rect 8309 13481 8343 13515
rect 9045 13481 9079 13515
rect 14657 13481 14691 13515
rect 16313 13481 16347 13515
rect 16957 13481 16991 13515
rect 18797 13481 18831 13515
rect 20545 13481 20579 13515
rect 2237 13413 2271 13447
rect 9965 13413 9999 13447
rect 10517 13413 10551 13447
rect 13544 13413 13578 13447
rect 15945 13413 15979 13447
rect 17316 13413 17350 13447
rect 20177 13413 20211 13447
rect 1409 13345 1443 13379
rect 1961 13345 1995 13379
rect 3525 13345 3559 13379
rect 5172 13345 5206 13379
rect 6909 13345 6943 13379
rect 8493 13345 8527 13379
rect 8953 13345 8987 13379
rect 9597 13345 9631 13379
rect 12725 13345 12759 13379
rect 19441 13345 19475 13379
rect 4905 13277 4939 13311
rect 6653 13277 6687 13311
rect 9229 13277 9263 13311
rect 1593 13209 1627 13243
rect 3157 13209 3191 13243
rect 6285 13209 6319 13243
rect 10057 13277 10091 13311
rect 12817 13277 12851 13311
rect 13001 13277 13035 13311
rect 13277 13277 13311 13311
rect 14933 13277 14967 13311
rect 17049 13277 17083 13311
rect 21097 13277 21131 13311
rect 11805 13209 11839 13243
rect 19809 13209 19843 13243
rect 3893 13141 3927 13175
rect 8033 13141 8067 13175
rect 8585 13141 8619 13175
rect 9505 13141 9539 13175
rect 12357 13141 12391 13175
rect 15485 13141 15519 13175
rect 18429 13141 18463 13175
rect 19073 13141 19107 13175
rect 1685 12937 1719 12971
rect 5917 12937 5951 12971
rect 9597 12937 9631 12971
rect 13737 12937 13771 12971
rect 13829 12937 13863 12971
rect 16773 12937 16807 12971
rect 17141 12937 17175 12971
rect 18061 12937 18095 12971
rect 19073 12937 19107 12971
rect 9873 12869 9907 12903
rect 13461 12869 13495 12903
rect 2237 12801 2271 12835
rect 3065 12801 3099 12835
rect 4169 12801 4203 12835
rect 4537 12801 4571 12835
rect 7665 12801 7699 12835
rect 10609 12801 10643 12835
rect 13093 12801 13127 12835
rect 20177 12869 20211 12903
rect 14289 12801 14323 12835
rect 14381 12801 14415 12835
rect 14841 12801 14875 12835
rect 18705 12801 18739 12835
rect 19441 12801 19475 12835
rect 1501 12733 1535 12767
rect 2053 12733 2087 12767
rect 3433 12733 3467 12767
rect 6193 12733 6227 12767
rect 8217 12733 8251 12767
rect 8473 12733 8507 12767
rect 10701 12733 10735 12767
rect 12817 12733 12851 12767
rect 13645 12733 13679 12767
rect 13737 12733 13771 12767
rect 14197 12733 14231 12767
rect 15393 12733 15427 12767
rect 15761 12733 15795 12767
rect 18429 12733 18463 12767
rect 20913 12733 20947 12767
rect 3893 12665 3927 12699
rect 4804 12665 4838 12699
rect 10968 12665 11002 12699
rect 18521 12665 18555 12699
rect 20545 12665 20579 12699
rect 3525 12597 3559 12631
rect 3985 12597 4019 12631
rect 7205 12597 7239 12631
rect 7757 12597 7791 12631
rect 12081 12597 12115 12631
rect 12449 12597 12483 12631
rect 12909 12597 12943 12631
rect 16129 12597 16163 12631
rect 16497 12597 16531 12631
rect 17601 12597 17635 12631
rect 19809 12597 19843 12631
rect 1777 12393 1811 12427
rect 3065 12393 3099 12427
rect 5549 12393 5583 12427
rect 5825 12393 5859 12427
rect 9321 12393 9355 12427
rect 13737 12393 13771 12427
rect 16865 12393 16899 12427
rect 17509 12393 17543 12427
rect 20545 12393 20579 12427
rect 21189 12393 21223 12427
rect 1593 12257 1627 12291
rect 2145 12257 2179 12291
rect 2881 12257 2915 12291
rect 4333 12257 4367 12291
rect 2329 12189 2363 12223
rect 4077 12189 4111 12223
rect 5457 12121 5491 12155
rect 14197 12325 14231 12359
rect 5917 12257 5951 12291
rect 6184 12257 6218 12291
rect 7757 12257 7791 12291
rect 8585 12257 8619 12291
rect 10609 12257 10643 12291
rect 11621 12257 11655 12291
rect 11888 12257 11922 12291
rect 14105 12257 14139 12291
rect 14933 12257 14967 12291
rect 15485 12257 15519 12291
rect 15752 12257 15786 12291
rect 17877 12257 17911 12291
rect 19432 12257 19466 12291
rect 8677 12189 8711 12223
rect 8861 12189 8895 12223
rect 10701 12189 10735 12223
rect 10885 12189 10919 12223
rect 13553 12189 13587 12223
rect 14289 12189 14323 12223
rect 17969 12189 18003 12223
rect 18153 12189 18187 12223
rect 18521 12189 18555 12223
rect 19165 12189 19199 12223
rect 8217 12121 8251 12155
rect 11253 12121 11287 12155
rect 18981 12121 19015 12155
rect 3525 12053 3559 12087
rect 3801 12053 3835 12087
rect 5549 12053 5583 12087
rect 7297 12053 7331 12087
rect 7573 12053 7607 12087
rect 8033 12053 8067 12087
rect 9873 12053 9907 12087
rect 10241 12053 10275 12087
rect 13001 12053 13035 12087
rect 14749 12053 14783 12087
rect 17417 12053 17451 12087
rect 6377 11849 6411 11883
rect 6561 11849 6595 11883
rect 9229 11849 9263 11883
rect 10149 11849 10183 11883
rect 12081 11849 12115 11883
rect 12449 11849 12483 11883
rect 19441 11849 19475 11883
rect 4169 11781 4203 11815
rect 4997 11713 5031 11747
rect 5917 11713 5951 11747
rect 6101 11713 6135 11747
rect 1961 11645 1995 11679
rect 2789 11645 2823 11679
rect 2237 11577 2271 11611
rect 3056 11577 3090 11611
rect 9505 11781 9539 11815
rect 11897 11781 11931 11815
rect 16313 11781 16347 11815
rect 17785 11781 17819 11815
rect 20821 11781 20855 11815
rect 7389 11713 7423 11747
rect 7757 11713 7791 11747
rect 7849 11713 7883 11747
rect 13001 11713 13035 11747
rect 13829 11713 13863 11747
rect 17141 11713 17175 11747
rect 7297 11645 7331 11679
rect 10241 11645 10275 11679
rect 10508 11645 10542 11679
rect 12265 11645 12299 11679
rect 12817 11645 12851 11679
rect 14105 11645 14139 11679
rect 14933 11645 14967 11679
rect 18061 11645 18095 11679
rect 20453 11645 20487 11679
rect 8116 11577 8150 11611
rect 13645 11577 13679 11611
rect 13737 11577 13771 11611
rect 14381 11577 14415 11611
rect 15200 11577 15234 11611
rect 18328 11577 18362 11611
rect 20085 11577 20119 11611
rect 1685 11509 1719 11543
rect 4445 11509 4479 11543
rect 4813 11509 4847 11543
rect 4905 11509 4939 11543
rect 5457 11509 5491 11543
rect 5825 11509 5859 11543
rect 6377 11509 6411 11543
rect 6837 11509 6871 11543
rect 7205 11509 7239 11543
rect 7757 11509 7791 11543
rect 11621 11509 11655 11543
rect 12909 11509 12943 11543
rect 13277 11509 13311 11543
rect 16589 11509 16623 11543
rect 16957 11509 16991 11543
rect 17049 11509 17083 11543
rect 19809 11509 19843 11543
rect 21189 11509 21223 11543
rect 2697 11305 2731 11339
rect 4261 11305 4295 11339
rect 4629 11305 4663 11339
rect 5273 11305 5307 11339
rect 5733 11305 5767 11339
rect 6377 11305 6411 11339
rect 2053 11237 2087 11271
rect 1777 11169 1811 11203
rect 2513 11169 2547 11203
rect 4721 11169 4755 11203
rect 5917 11169 5951 11203
rect 6285 11169 6319 11203
rect 3157 11101 3191 11135
rect 3525 11101 3559 11135
rect 4905 11101 4939 11135
rect 7389 11305 7423 11339
rect 8953 11305 8987 11339
rect 9321 11305 9355 11339
rect 10517 11305 10551 11339
rect 11529 11305 11563 11339
rect 11989 11305 12023 11339
rect 13645 11305 13679 11339
rect 14197 11305 14231 11339
rect 15301 11305 15335 11339
rect 16313 11305 16347 11339
rect 17233 11305 17267 11339
rect 17509 11305 17543 11339
rect 18981 11305 19015 11339
rect 19625 11305 19659 11339
rect 20453 11305 20487 11339
rect 1685 10965 1719 10999
rect 3893 10965 3927 10999
rect 6377 10965 6411 10999
rect 6469 11237 6503 11271
rect 6929 11169 6963 11203
rect 10241 11237 10275 11271
rect 12357 11237 12391 11271
rect 12449 11237 12483 11271
rect 17877 11237 17911 11271
rect 19257 11237 19291 11271
rect 7573 11169 7607 11203
rect 7840 11169 7874 11203
rect 11161 11169 11195 11203
rect 13093 11169 13127 11203
rect 13553 11169 13587 11203
rect 14565 11169 14599 11203
rect 14657 11169 14691 11203
rect 15669 11169 15703 11203
rect 16957 11169 16991 11203
rect 18613 11169 18647 11203
rect 7021 11101 7055 11135
rect 7205 11101 7239 11135
rect 7389 11101 7423 11135
rect 12541 11101 12575 11135
rect 13737 11101 13771 11135
rect 14841 11101 14875 11135
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 17969 11101 18003 11135
rect 18153 11101 18187 11135
rect 13185 11033 13219 11067
rect 19993 11033 20027 11067
rect 21097 11033 21131 11067
rect 6469 10965 6503 10999
rect 6561 10965 6595 10999
rect 9873 10965 9907 10999
rect 16773 10965 16807 10999
rect 5181 10761 5215 10795
rect 6193 10761 6227 10795
rect 9505 10761 9539 10795
rect 10793 10761 10827 10795
rect 15485 10761 15519 10795
rect 20545 10761 20579 10795
rect 4445 10693 4479 10727
rect 6653 10693 6687 10727
rect 8217 10693 8251 10727
rect 8401 10693 8435 10727
rect 8493 10693 8527 10727
rect 19809 10693 19843 10727
rect 20177 10693 20211 10727
rect 1685 10625 1719 10659
rect 2789 10625 2823 10659
rect 3893 10625 3927 10659
rect 4077 10625 4111 10659
rect 6837 10625 6871 10659
rect 1409 10557 1443 10591
rect 9045 10625 9079 10659
rect 10057 10625 10091 10659
rect 11437 10625 11471 10659
rect 14105 10625 14139 10659
rect 18061 10625 18095 10659
rect 8861 10557 8895 10591
rect 8953 10557 8987 10591
rect 11161 10557 11195 10591
rect 12449 10557 12483 10591
rect 15761 10557 15795 10591
rect 18328 10557 18362 10591
rect 2513 10489 2547 10523
rect 4905 10489 4939 10523
rect 7104 10489 7138 10523
rect 8401 10489 8435 10523
rect 9965 10489 9999 10523
rect 10517 10489 10551 10523
rect 11253 10489 11287 10523
rect 12716 10489 12750 10523
rect 14372 10489 14406 10523
rect 16028 10489 16062 10523
rect 2145 10421 2179 10455
rect 2605 10421 2639 10455
rect 3249 10421 3283 10455
rect 3433 10421 3467 10455
rect 3801 10421 3835 10455
rect 5641 10421 5675 10455
rect 9873 10421 9907 10455
rect 11897 10421 11931 10455
rect 13829 10421 13863 10455
rect 17141 10421 17175 10455
rect 17417 10421 17451 10455
rect 19441 10421 19475 10455
rect 2329 10217 2363 10251
rect 8033 10217 8067 10251
rect 8493 10217 8527 10251
rect 13093 10217 13127 10251
rect 17785 10217 17819 10251
rect 18153 10217 18187 10251
rect 18797 10217 18831 10251
rect 19257 10217 19291 10251
rect 19625 10217 19659 10251
rect 19993 10217 20027 10251
rect 1777 10149 1811 10183
rect 4344 10149 4378 10183
rect 13636 10149 13670 10183
rect 15117 10149 15151 10183
rect 15853 10149 15887 10183
rect 16672 10149 16706 10183
rect 2237 10081 2271 10115
rect 3249 10081 3283 10115
rect 4077 10081 4111 10115
rect 6000 10081 6034 10115
rect 7941 10081 7975 10115
rect 8401 10081 8435 10115
rect 9045 10081 9079 10115
rect 10057 10081 10091 10115
rect 10324 10081 10358 10115
rect 11713 10081 11747 10115
rect 11980 10081 12014 10115
rect 13369 10081 13403 10115
rect 15761 10081 15795 10115
rect 16405 10081 16439 10115
rect 18521 10081 18555 10115
rect 2513 10013 2547 10047
rect 3341 10013 3375 10047
rect 3433 10013 3467 10047
rect 5733 10013 5767 10047
rect 8585 10013 8619 10047
rect 16037 10013 16071 10047
rect 1869 9945 1903 9979
rect 7113 9945 7147 9979
rect 9413 9945 9447 9979
rect 14749 9945 14783 9979
rect 2881 9877 2915 9911
rect 5457 9877 5491 9911
rect 7389 9877 7423 9911
rect 7757 9877 7791 9911
rect 9965 9877 9999 9911
rect 11437 9877 11471 9911
rect 15393 9877 15427 9911
rect 1777 9673 1811 9707
rect 16405 9673 16439 9707
rect 17601 9673 17635 9707
rect 18705 9673 18739 9707
rect 4537 9605 4571 9639
rect 5549 9605 5583 9639
rect 11437 9605 11471 9639
rect 13645 9605 13679 9639
rect 14841 9605 14875 9639
rect 16589 9605 16623 9639
rect 4169 9537 4203 9571
rect 5181 9537 5215 9571
rect 6377 9537 6411 9571
rect 7389 9537 7423 9571
rect 8677 9537 8711 9571
rect 10793 9537 10827 9571
rect 10977 9537 11011 9571
rect 12909 9537 12943 9571
rect 13093 9537 13127 9571
rect 14381 9537 14415 9571
rect 15669 9537 15703 9571
rect 17141 9537 17175 9571
rect 18245 9537 18279 9571
rect 19073 9537 19107 9571
rect 1869 9469 1903 9503
rect 2125 9469 2159 9503
rect 3893 9469 3927 9503
rect 5457 9469 5491 9503
rect 6101 9469 6135 9503
rect 7205 9469 7239 9503
rect 11713 9469 11747 9503
rect 12081 9469 12115 9503
rect 12817 9469 12851 9503
rect 14197 9469 14231 9503
rect 16957 9469 16991 9503
rect 8944 9401 8978 9435
rect 17049 9401 17083 9435
rect 3249 9333 3283 9367
rect 3525 9333 3559 9367
rect 3985 9333 4019 9367
rect 4905 9333 4939 9367
rect 4997 9333 5031 9367
rect 5457 9333 5491 9367
rect 5733 9333 5767 9367
rect 6193 9333 6227 9367
rect 6837 9333 6871 9367
rect 7297 9333 7331 9367
rect 7849 9333 7883 9367
rect 8125 9333 8159 9367
rect 10057 9333 10091 9367
rect 10333 9333 10367 9367
rect 10701 9333 10735 9367
rect 12449 9333 12483 9367
rect 15209 9333 15243 9367
rect 16037 9333 16071 9367
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 3525 9129 3559 9163
rect 5733 9129 5767 9163
rect 6009 9129 6043 9163
rect 6377 9129 6411 9163
rect 6561 9129 6595 9163
rect 7297 9129 7331 9163
rect 9873 9129 9907 9163
rect 10241 9129 10275 9163
rect 11069 9129 11103 9163
rect 11529 9129 11563 9163
rect 12817 9129 12851 9163
rect 13185 9129 13219 9163
rect 13553 9129 13587 9163
rect 14473 9129 14507 9163
rect 15669 9129 15703 9163
rect 16037 9129 16071 9163
rect 17049 9129 17083 9163
rect 17325 9129 17359 9163
rect 18153 9129 18187 9163
rect 1685 9061 1719 9095
rect 14841 9061 14875 9095
rect 1777 8993 1811 9027
rect 8861 8993 8895 9027
rect 16405 8993 16439 9027
rect 17693 8993 17727 9027
rect 7665 8925 7699 8959
rect 8309 8925 8343 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 12449 8925 12483 8959
rect 4353 8857 4387 8891
rect 10793 8857 10827 8891
rect 1961 8789 1995 8823
rect 3893 8789 3927 8823
rect 4905 8789 4939 8823
rect 5365 8789 5399 8823
rect 8493 8789 8527 8823
rect 11897 8789 11931 8823
rect 13921 8789 13955 8823
rect 1777 8585 1811 8619
rect 3893 8585 3927 8619
rect 6929 8585 6963 8619
rect 9321 8585 9355 8619
rect 10425 8585 10459 8619
rect 11161 8585 11195 8619
rect 11989 8585 12023 8619
rect 13185 8585 13219 8619
rect 13737 8585 13771 8619
rect 14473 8585 14507 8619
rect 16037 8585 16071 8619
rect 16405 8585 16439 8619
rect 16865 8585 16899 8619
rect 17233 8585 17267 8619
rect 3617 8517 3651 8551
rect 10057 8517 10091 8551
rect 10701 8517 10735 8551
rect 11713 8517 11747 8551
rect 12817 8517 12851 8551
rect 14749 8517 14783 8551
rect 5365 8449 5399 8483
rect 6101 8449 6135 8483
rect 6561 8449 6595 8483
rect 7573 8449 7607 8483
rect 15117 8449 15151 8483
rect 2237 8381 2271 8415
rect 7297 8381 7331 8415
rect 7941 8381 7975 8415
rect 15485 8381 15519 8415
rect 2145 8313 2179 8347
rect 2482 8313 2516 8347
rect 5089 8313 5123 8347
rect 5181 8313 5215 8347
rect 5825 8313 5859 8347
rect 7389 8313 7423 8347
rect 8208 8313 8242 8347
rect 14013 8313 14047 8347
rect 4261 8245 4295 8279
rect 4721 8245 4755 8279
rect 9597 8245 9631 8279
rect 1685 8041 1719 8075
rect 3341 8041 3375 8075
rect 8493 8041 8527 8075
rect 9873 8041 9907 8075
rect 11713 8041 11747 8075
rect 12081 8041 12115 8075
rect 12541 8041 12575 8075
rect 13277 8041 13311 8075
rect 13553 8041 13587 8075
rect 13921 8041 13955 8075
rect 14657 8041 14691 8075
rect 15577 8041 15611 8075
rect 15945 8041 15979 8075
rect 12265 7973 12299 8007
rect 1501 7905 1535 7939
rect 2053 7905 2087 7939
rect 3433 7905 3467 7939
rect 4445 7905 4479 7939
rect 4537 7905 4571 7939
rect 5356 7905 5390 7939
rect 7113 7905 7147 7939
rect 7380 7905 7414 7939
rect 2329 7837 2363 7871
rect 2881 7837 2915 7871
rect 3525 7837 3559 7871
rect 4629 7837 4663 7871
rect 5089 7837 5123 7871
rect 10701 7837 10735 7871
rect 11345 7837 11379 7871
rect 12817 7905 12851 7939
rect 14289 7837 14323 7871
rect 8953 7769 8987 7803
rect 11069 7769 11103 7803
rect 12265 7769 12299 7803
rect 2973 7701 3007 7735
rect 4077 7701 4111 7735
rect 6469 7701 6503 7735
rect 6929 7701 6963 7735
rect 9229 7701 9263 7735
rect 10241 7701 10275 7735
rect 15025 7701 15059 7735
rect 1777 7497 1811 7531
rect 4445 7497 4479 7531
rect 4629 7497 4663 7531
rect 9505 7497 9539 7531
rect 11253 7497 11287 7531
rect 11805 7497 11839 7531
rect 12265 7497 12299 7531
rect 12725 7497 12759 7531
rect 13185 7497 13219 7531
rect 13461 7497 13495 7531
rect 18705 7497 18739 7531
rect 3065 7361 3099 7395
rect 8493 7429 8527 7463
rect 19073 7429 19107 7463
rect 6837 7361 6871 7395
rect 9045 7361 9079 7395
rect 9965 7361 9999 7395
rect 10149 7361 10183 7395
rect 10517 7361 10551 7395
rect 13829 7361 13863 7395
rect 14197 7361 14231 7395
rect 14565 7361 14599 7395
rect 1869 7293 1903 7327
rect 3332 7293 3366 7327
rect 4629 7293 4663 7327
rect 4721 7293 4755 7327
rect 4977 7293 5011 7327
rect 6377 7293 6411 7327
rect 18521 7293 18555 7327
rect 2145 7225 2179 7259
rect 7104 7225 7138 7259
rect 10885 7225 10919 7259
rect 2881 7157 2915 7191
rect 6101 7157 6135 7191
rect 8217 7157 8251 7191
rect 8861 7157 8895 7191
rect 8953 7157 8987 7191
rect 9873 7157 9907 7191
rect 3433 6953 3467 6987
rect 5273 6953 5307 6987
rect 5733 6953 5767 6987
rect 3709 6885 3743 6919
rect 4721 6885 4755 6919
rect 4813 6885 4847 6919
rect 1593 6817 1627 6851
rect 2053 6817 2087 6851
rect 2513 6817 2547 6851
rect 2973 6817 3007 6851
rect 6837 6885 6871 6919
rect 6101 6817 6135 6851
rect 6745 6817 6779 6851
rect 7205 6817 7239 6851
rect 7665 6817 7699 6851
rect 8677 6817 8711 6851
rect 9321 6817 9355 6851
rect 10333 6817 10367 6851
rect 12449 6817 12483 6851
rect 13185 6817 13219 6851
rect 19073 6817 19107 6851
rect 19625 6817 19659 6851
rect 4905 6749 4939 6783
rect 5273 6749 5307 6783
rect 4353 6681 4387 6715
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 8769 6749 8803 6783
rect 8861 6749 8895 6783
rect 12725 6749 12759 6783
rect 8309 6681 8343 6715
rect 9873 6681 9907 6715
rect 19809 6681 19843 6715
rect 5365 6613 5399 6647
rect 7113 6613 7147 6647
rect 7297 6613 7331 6647
rect 10609 6613 10643 6647
rect 11069 6613 11103 6647
rect 11345 6613 11379 6647
rect 11713 6613 11747 6647
rect 13553 6613 13587 6647
rect 13829 6613 13863 6647
rect 19257 6613 19291 6647
rect 1685 6409 1719 6443
rect 2513 6409 2547 6443
rect 3525 6409 3559 6443
rect 5549 6409 5583 6443
rect 6101 6409 6135 6443
rect 6653 6409 6687 6443
rect 8309 6409 8343 6443
rect 9045 6409 9079 6443
rect 9413 6409 9447 6443
rect 9689 6409 9723 6443
rect 9873 6409 9907 6443
rect 10241 6409 10275 6443
rect 10609 6409 10643 6443
rect 12725 6409 12759 6443
rect 19625 6409 19659 6443
rect 20085 6409 20119 6443
rect 2145 6341 2179 6375
rect 3433 6341 3467 6375
rect 7113 6341 7147 6375
rect 7297 6341 7331 6375
rect 11345 6341 11379 6375
rect 11805 6341 11839 6375
rect 12173 6341 12207 6375
rect 3065 6273 3099 6307
rect 3985 6273 4019 6307
rect 4077 6273 4111 6307
rect 7849 6273 7883 6307
rect 9689 6273 9723 6307
rect 3893 6205 3927 6239
rect 7665 6205 7699 6239
rect 10885 6205 10919 6239
rect 19901 6205 19935 6239
rect 20453 6205 20487 6239
rect 8677 6137 8711 6171
rect 4721 6069 4755 6103
rect 5089 6069 5123 6103
rect 7757 6069 7791 6103
rect 19073 6069 19107 6103
rect 1593 5865 1627 5899
rect 2329 5865 2363 5899
rect 2789 5865 2823 5899
rect 3433 5865 3467 5899
rect 3893 5865 3927 5899
rect 5181 5865 5215 5899
rect 5641 5865 5675 5899
rect 6193 5865 6227 5899
rect 6561 5865 6595 5899
rect 7297 5865 7331 5899
rect 8125 5865 8159 5899
rect 8769 5865 8803 5899
rect 10701 5865 10735 5899
rect 11069 5865 11103 5899
rect 11437 5865 11471 5899
rect 20453 5865 20487 5899
rect 1961 5797 1995 5831
rect 3157 5797 3191 5831
rect 4353 5729 4387 5763
rect 7021 5729 7055 5763
rect 8401 5729 8435 5763
rect 20269 5729 20303 5763
rect 4905 5661 4939 5695
rect 9137 5661 9171 5695
rect 7665 5525 7699 5559
rect 9873 5525 9907 5559
rect 10241 5525 10275 5559
rect 2237 5321 2271 5355
rect 2605 5321 2639 5355
rect 2973 5321 3007 5355
rect 4537 5321 4571 5355
rect 6009 5321 6043 5355
rect 7113 5321 7147 5355
rect 7941 5321 7975 5355
rect 8309 5321 8343 5355
rect 8585 5321 8619 5355
rect 8953 5321 8987 5355
rect 9321 5321 9355 5355
rect 20729 5321 20763 5355
rect 3341 5253 3375 5287
rect 6377 5253 6411 5287
rect 1685 5185 1719 5219
rect 3617 5185 3651 5219
rect 4169 5185 4203 5219
rect 4813 5185 4847 5219
rect 5181 5185 5215 5219
rect 5549 5185 5583 5219
rect 7481 5185 7515 5219
rect 20545 5117 20579 5151
rect 21097 5117 21131 5151
rect 20269 5049 20303 5083
rect 1869 4777 1903 4811
rect 2237 4777 2271 4811
rect 2605 4777 2639 4811
rect 2973 4777 3007 4811
rect 3249 4777 3283 4811
rect 4905 4777 4939 4811
rect 5273 4777 5307 4811
rect 5641 4777 5675 4811
rect 6561 4777 6595 4811
rect 6929 4777 6963 4811
rect 7297 4777 7331 4811
rect 7665 4777 7699 4811
rect 8033 4777 8067 4811
rect 6101 4709 6135 4743
rect 3709 4437 3743 4471
rect 4537 4437 4571 4471
rect 7481 4233 7515 4267
rect 7849 4233 7883 4267
rect 2789 4165 2823 4199
rect 3157 4165 3191 4199
rect 1593 4097 1627 4131
rect 2329 4097 2363 4131
rect 3525 4097 3559 4131
rect 3985 4097 4019 4131
rect 4997 4097 5031 4131
rect 5365 4097 5399 4131
rect 5733 4097 5767 4131
rect 7021 4097 7055 4131
rect 2973 3689 3007 3723
rect 5089 3689 5123 3723
<< metal1 >>
rect 4062 20340 4068 20392
rect 4120 20380 4126 20392
rect 20070 20380 20076 20392
rect 4120 20352 20076 20380
rect 4120 20340 4126 20352
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 8202 20272 8208 20324
rect 8260 20312 8266 20324
rect 15286 20312 15292 20324
rect 8260 20284 15292 20312
rect 8260 20272 8266 20284
rect 15286 20272 15292 20284
rect 15344 20272 15350 20324
rect 7190 20204 7196 20256
rect 7248 20244 7254 20256
rect 15102 20244 15108 20256
rect 7248 20216 15108 20244
rect 7248 20204 7254 20216
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1670 20040 1676 20052
rect 1631 20012 1676 20040
rect 1670 20000 1676 20012
rect 1728 20000 1734 20052
rect 5261 20043 5319 20049
rect 5261 20009 5273 20043
rect 5307 20009 5319 20043
rect 5261 20003 5319 20009
rect 2314 19972 2320 19984
rect 1504 19944 2320 19972
rect 1504 19913 1532 19944
rect 2314 19932 2320 19944
rect 2372 19932 2378 19984
rect 4525 19975 4583 19981
rect 4525 19941 4537 19975
rect 4571 19972 4583 19975
rect 5276 19972 5304 20003
rect 5626 20000 5632 20052
rect 5684 20040 5690 20052
rect 5721 20043 5779 20049
rect 5721 20040 5733 20043
rect 5684 20012 5733 20040
rect 5684 20000 5690 20012
rect 5721 20009 5733 20012
rect 5767 20040 5779 20043
rect 6273 20043 6331 20049
rect 6273 20040 6285 20043
rect 5767 20012 6285 20040
rect 5767 20009 5779 20012
rect 5721 20003 5779 20009
rect 6273 20009 6285 20012
rect 6319 20009 6331 20043
rect 8386 20040 8392 20052
rect 8299 20012 8392 20040
rect 6273 20003 6331 20009
rect 8386 20000 8392 20012
rect 8444 20040 8450 20052
rect 8846 20040 8852 20052
rect 8444 20012 8852 20040
rect 8444 20000 8450 20012
rect 8846 20000 8852 20012
rect 8904 20000 8910 20052
rect 9306 20040 9312 20052
rect 9267 20012 9312 20040
rect 9306 20000 9312 20012
rect 9364 20000 9370 20052
rect 9493 20043 9551 20049
rect 9493 20009 9505 20043
rect 9539 20040 9551 20043
rect 9674 20040 9680 20052
rect 9539 20012 9680 20040
rect 9539 20009 9551 20012
rect 9493 20003 9551 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 13354 20000 13360 20052
rect 13412 20040 13418 20052
rect 13449 20043 13507 20049
rect 13449 20040 13461 20043
rect 13412 20012 13461 20040
rect 13412 20000 13418 20012
rect 13449 20009 13461 20012
rect 13495 20009 13507 20043
rect 13449 20003 13507 20009
rect 14001 20043 14059 20049
rect 14001 20009 14013 20043
rect 14047 20040 14059 20043
rect 14274 20040 14280 20052
rect 14047 20012 14280 20040
rect 14047 20009 14059 20012
rect 14001 20003 14059 20009
rect 14274 20000 14280 20012
rect 14332 20000 14338 20052
rect 15102 20040 15108 20052
rect 15063 20012 15108 20040
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15286 20000 15292 20052
rect 15344 20040 15350 20052
rect 15657 20043 15715 20049
rect 15657 20040 15669 20043
rect 15344 20012 15669 20040
rect 15344 20000 15350 20012
rect 15657 20009 15669 20012
rect 15703 20009 15715 20043
rect 15657 20003 15715 20009
rect 16301 20043 16359 20049
rect 16301 20009 16313 20043
rect 16347 20040 16359 20043
rect 16574 20040 16580 20052
rect 16347 20012 16580 20040
rect 16347 20009 16359 20012
rect 16301 20003 16359 20009
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 17034 20000 17040 20052
rect 17092 20040 17098 20052
rect 17405 20043 17463 20049
rect 17405 20040 17417 20043
rect 17092 20012 17417 20040
rect 17092 20000 17098 20012
rect 17405 20009 17417 20012
rect 17451 20009 17463 20043
rect 17405 20003 17463 20009
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18012 20012 18521 20040
rect 18012 20000 18018 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 20070 20040 20076 20052
rect 20031 20012 20076 20040
rect 18509 20003 18567 20009
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 9585 19975 9643 19981
rect 4571 19944 6868 19972
rect 4571 19941 4583 19944
rect 4525 19935 4583 19941
rect 1489 19907 1547 19913
rect 1489 19873 1501 19907
rect 1535 19873 1547 19907
rect 1489 19867 1547 19873
rect 2041 19907 2099 19913
rect 2041 19873 2053 19907
rect 2087 19904 2099 19907
rect 2866 19904 2872 19916
rect 2087 19876 2872 19904
rect 2087 19873 2099 19876
rect 2041 19867 2099 19873
rect 2866 19864 2872 19876
rect 2924 19904 2930 19916
rect 4062 19904 4068 19916
rect 2924 19876 4068 19904
rect 2924 19864 2930 19876
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 4246 19864 4252 19916
rect 4304 19904 4310 19916
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 4304 19876 4445 19904
rect 4304 19864 4310 19876
rect 4433 19873 4445 19876
rect 4479 19904 4491 19907
rect 5077 19907 5135 19913
rect 5077 19904 5089 19907
rect 4479 19876 5089 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 5077 19873 5089 19876
rect 5123 19873 5135 19907
rect 5077 19867 5135 19873
rect 5629 19907 5687 19913
rect 5629 19873 5641 19907
rect 5675 19873 5687 19907
rect 5629 19867 5687 19873
rect 1394 19796 1400 19848
rect 1452 19836 1458 19848
rect 2225 19839 2283 19845
rect 2225 19836 2237 19839
rect 1452 19808 2237 19836
rect 1452 19796 1458 19808
rect 2225 19805 2237 19808
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 4982 19836 4988 19848
rect 4755 19808 4988 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 3421 19771 3479 19777
rect 3421 19737 3433 19771
rect 3467 19768 3479 19771
rect 3881 19771 3939 19777
rect 3881 19768 3893 19771
rect 3467 19740 3893 19768
rect 3467 19737 3479 19740
rect 3421 19731 3479 19737
rect 3881 19737 3893 19740
rect 3927 19768 3939 19771
rect 4724 19768 4752 19799
rect 4982 19796 4988 19808
rect 5040 19796 5046 19848
rect 3927 19740 4752 19768
rect 3927 19737 3939 19740
rect 3881 19731 3939 19737
rect 4890 19728 4896 19780
rect 4948 19768 4954 19780
rect 5644 19768 5672 19867
rect 5905 19839 5963 19845
rect 5905 19805 5917 19839
rect 5951 19836 5963 19839
rect 5951 19808 6776 19836
rect 5951 19805 5963 19808
rect 5905 19799 5963 19805
rect 4948 19740 5672 19768
rect 4948 19728 4954 19740
rect 6748 19712 6776 19808
rect 6840 19768 6868 19944
rect 9585 19941 9597 19975
rect 9631 19972 9643 19975
rect 10873 19975 10931 19981
rect 10873 19972 10885 19975
rect 9631 19944 10885 19972
rect 9631 19941 9643 19944
rect 9585 19935 9643 19941
rect 10873 19941 10885 19944
rect 10919 19941 10931 19975
rect 10873 19935 10931 19941
rect 11054 19932 11060 19984
rect 11112 19972 11118 19984
rect 11701 19975 11759 19981
rect 11701 19972 11713 19975
rect 11112 19944 11713 19972
rect 11112 19932 11118 19944
rect 11701 19941 11713 19944
rect 11747 19941 11759 19975
rect 17310 19972 17316 19984
rect 17223 19944 17316 19972
rect 11701 19935 11759 19941
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 13265 19907 13323 19913
rect 9732 19876 12756 19904
rect 9732 19864 9738 19876
rect 9122 19796 9128 19848
rect 9180 19836 9186 19848
rect 9769 19839 9827 19845
rect 9769 19836 9781 19839
rect 9180 19808 9781 19836
rect 9180 19796 9186 19808
rect 9769 19805 9781 19808
rect 9815 19805 9827 19839
rect 9769 19799 9827 19805
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19836 11115 19839
rect 12618 19836 12624 19848
rect 11103 19808 12624 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 12728 19836 12756 19876
rect 13265 19873 13277 19907
rect 13311 19904 13323 19907
rect 13354 19904 13360 19916
rect 13311 19876 13360 19904
rect 13311 19873 13323 19876
rect 13265 19867 13323 19873
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 13817 19907 13875 19913
rect 13817 19873 13829 19907
rect 13863 19904 13875 19907
rect 14458 19904 14464 19916
rect 13863 19876 14464 19904
rect 13863 19873 13875 19876
rect 13817 19867 13875 19873
rect 14458 19864 14464 19876
rect 14516 19904 14522 19916
rect 15102 19904 15108 19916
rect 14516 19876 15108 19904
rect 14516 19864 14522 19876
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 16117 19907 16175 19913
rect 16117 19873 16129 19907
rect 16163 19904 16175 19907
rect 16574 19904 16580 19916
rect 16163 19876 16580 19904
rect 16163 19873 16175 19876
rect 16117 19867 16175 19873
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 17236 19913 17264 19944
rect 17310 19932 17316 19944
rect 17368 19972 17374 19984
rect 20809 19975 20867 19981
rect 20809 19972 20821 19975
rect 17368 19944 20821 19972
rect 17368 19932 17374 19944
rect 20809 19941 20821 19944
rect 20855 19941 20867 19975
rect 20809 19935 20867 19941
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19873 17279 19907
rect 17221 19867 17279 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18690 19904 18696 19916
rect 18371 19876 18696 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18690 19864 18696 19876
rect 18748 19864 18754 19916
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19904 18935 19907
rect 18966 19904 18972 19916
rect 18923 19876 18972 19904
rect 18923 19873 18935 19876
rect 18877 19867 18935 19873
rect 18966 19864 18972 19876
rect 19024 19864 19030 19916
rect 14737 19839 14795 19845
rect 14737 19836 14749 19839
rect 12728 19808 14749 19836
rect 14737 19805 14749 19808
rect 14783 19805 14795 19839
rect 14737 19799 14795 19805
rect 9585 19771 9643 19777
rect 9585 19768 9597 19771
rect 6840 19740 9597 19768
rect 9585 19737 9597 19740
rect 9631 19737 9643 19771
rect 9585 19731 9643 19737
rect 9858 19728 9864 19780
rect 9916 19768 9922 19780
rect 10597 19771 10655 19777
rect 10597 19768 10609 19771
rect 9916 19740 10609 19768
rect 9916 19728 9922 19740
rect 10597 19737 10609 19740
rect 10643 19737 10655 19771
rect 10597 19731 10655 19737
rect 10873 19771 10931 19777
rect 10873 19737 10885 19771
rect 10919 19768 10931 19771
rect 17773 19771 17831 19777
rect 17773 19768 17785 19771
rect 10919 19740 17785 19768
rect 10919 19737 10931 19740
rect 10873 19731 10931 19737
rect 17773 19737 17785 19740
rect 17819 19737 17831 19771
rect 17773 19731 17831 19737
rect 18414 19728 18420 19780
rect 18472 19768 18478 19780
rect 19061 19771 19119 19777
rect 19061 19768 19073 19771
rect 18472 19740 19073 19768
rect 18472 19728 18478 19740
rect 19061 19737 19073 19740
rect 19107 19737 19119 19771
rect 19061 19731 19119 19737
rect 2869 19703 2927 19709
rect 2869 19669 2881 19703
rect 2915 19700 2927 19703
rect 3602 19700 3608 19712
rect 2915 19672 3608 19700
rect 2915 19669 2927 19672
rect 2869 19663 2927 19669
rect 3602 19660 3608 19672
rect 3660 19660 3666 19712
rect 4062 19700 4068 19712
rect 4023 19672 4068 19700
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 6730 19700 6736 19712
rect 6691 19672 6736 19700
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 7098 19700 7104 19712
rect 7059 19672 7104 19700
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 7469 19703 7527 19709
rect 7469 19700 7481 19703
rect 7340 19672 7481 19700
rect 7340 19660 7346 19672
rect 7469 19669 7481 19672
rect 7515 19669 7527 19703
rect 7469 19663 7527 19669
rect 8021 19703 8079 19709
rect 8021 19669 8033 19703
rect 8067 19700 8079 19703
rect 8570 19700 8576 19712
rect 8067 19672 8576 19700
rect 8067 19669 8079 19672
rect 8021 19663 8079 19669
rect 8570 19660 8576 19672
rect 8628 19660 8634 19712
rect 8754 19700 8760 19712
rect 8715 19672 8760 19700
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 9398 19660 9404 19712
rect 9456 19700 9462 19712
rect 9493 19703 9551 19709
rect 9493 19700 9505 19703
rect 9456 19672 9505 19700
rect 9456 19660 9462 19672
rect 9493 19669 9505 19672
rect 9539 19669 9551 19703
rect 9493 19663 9551 19669
rect 10134 19660 10140 19712
rect 10192 19700 10198 19712
rect 10229 19703 10287 19709
rect 10229 19700 10241 19703
rect 10192 19672 10241 19700
rect 10192 19660 10198 19672
rect 10229 19669 10241 19672
rect 10275 19669 10287 19703
rect 10229 19663 10287 19669
rect 10410 19660 10416 19712
rect 10468 19700 10474 19712
rect 11333 19703 11391 19709
rect 11333 19700 11345 19703
rect 10468 19672 11345 19700
rect 10468 19660 10474 19672
rect 11333 19669 11345 19672
rect 11379 19669 11391 19703
rect 11333 19663 11391 19669
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 12069 19703 12127 19709
rect 12069 19700 12081 19703
rect 11848 19672 12081 19700
rect 11848 19660 11854 19672
rect 12069 19669 12081 19672
rect 12115 19669 12127 19703
rect 12069 19663 12127 19669
rect 12618 19660 12624 19712
rect 12676 19700 12682 19712
rect 12805 19703 12863 19709
rect 12805 19700 12817 19703
rect 12676 19672 12817 19700
rect 12676 19660 12682 19672
rect 12805 19669 12817 19672
rect 12851 19669 12863 19703
rect 14366 19700 14372 19712
rect 14327 19672 14372 19700
rect 12805 19663 12863 19669
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 16666 19700 16672 19712
rect 16627 19672 16672 19700
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 17034 19700 17040 19712
rect 16995 19672 17040 19700
rect 17034 19660 17040 19672
rect 17092 19660 17098 19712
rect 19794 19700 19800 19712
rect 19755 19672 19800 19700
rect 19794 19660 19800 19672
rect 19852 19660 19858 19712
rect 20438 19700 20444 19712
rect 20399 19672 20444 19700
rect 20438 19660 20444 19672
rect 20496 19660 20502 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 2222 19456 2228 19508
rect 2280 19496 2286 19508
rect 17034 19496 17040 19508
rect 2280 19468 17040 19496
rect 2280 19456 2286 19468
rect 17034 19456 17040 19468
rect 17092 19456 17098 19508
rect 19058 19496 19064 19508
rect 17144 19468 19064 19496
rect 9674 19388 9680 19440
rect 9732 19428 9738 19440
rect 17144 19428 17172 19468
rect 19058 19456 19064 19468
rect 19116 19456 19122 19508
rect 18690 19428 18696 19440
rect 9732 19400 9996 19428
rect 9732 19388 9738 19400
rect 2222 19360 2228 19372
rect 1504 19332 2228 19360
rect 1504 19301 1532 19332
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 4890 19320 4896 19372
rect 4948 19360 4954 19372
rect 8386 19360 8392 19372
rect 4948 19332 5212 19360
rect 8347 19332 8392 19360
rect 4948 19320 4954 19332
rect 1489 19295 1547 19301
rect 1489 19261 1501 19295
rect 1535 19261 1547 19295
rect 1489 19255 1547 19261
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19292 2099 19295
rect 2087 19264 2452 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 2314 19224 2320 19236
rect 2275 19196 2320 19224
rect 2314 19184 2320 19196
rect 2372 19184 2378 19236
rect 2424 19224 2452 19264
rect 2590 19252 2596 19304
rect 2648 19292 2654 19304
rect 3053 19295 3111 19301
rect 3053 19292 3065 19295
rect 2648 19264 3065 19292
rect 2648 19252 2654 19264
rect 3053 19261 3065 19264
rect 3099 19261 3111 19295
rect 4062 19292 4068 19304
rect 3053 19255 3111 19261
rect 3252 19264 4068 19292
rect 3252 19224 3280 19264
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 5074 19292 5080 19304
rect 5035 19264 5080 19292
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5184 19292 5212 19332
rect 8386 19320 8392 19332
rect 8444 19320 8450 19372
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19329 8631 19363
rect 8573 19323 8631 19329
rect 5184 19264 7604 19292
rect 2424 19196 3280 19224
rect 3320 19227 3378 19233
rect 3320 19193 3332 19227
rect 3366 19224 3378 19227
rect 5344 19227 5402 19233
rect 3366 19196 5028 19224
rect 3366 19193 3378 19196
rect 3320 19187 3378 19193
rect 5000 19168 5028 19196
rect 5344 19193 5356 19227
rect 5390 19224 5402 19227
rect 6730 19224 6736 19236
rect 5390 19196 6736 19224
rect 5390 19193 5402 19196
rect 5344 19187 5402 19193
rect 6730 19184 6736 19196
rect 6788 19224 6794 19236
rect 7377 19227 7435 19233
rect 7377 19224 7389 19227
rect 6788 19196 7389 19224
rect 6788 19184 6794 19196
rect 7377 19193 7389 19196
rect 7423 19193 7435 19227
rect 7576 19224 7604 19264
rect 7650 19252 7656 19304
rect 7708 19292 7714 19304
rect 7837 19295 7895 19301
rect 7837 19292 7849 19295
rect 7708 19264 7849 19292
rect 7708 19252 7714 19264
rect 7837 19261 7849 19264
rect 7883 19292 7895 19295
rect 8588 19292 8616 19323
rect 9306 19320 9312 19372
rect 9364 19360 9370 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 9364 19332 9413 19360
rect 9364 19320 9370 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 9585 19363 9643 19369
rect 9585 19329 9597 19363
rect 9631 19360 9643 19363
rect 9858 19360 9864 19372
rect 9631 19332 9864 19360
rect 9631 19329 9643 19332
rect 9585 19323 9643 19329
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 9968 19369 9996 19400
rect 16960 19400 17172 19428
rect 17236 19400 18696 19428
rect 9953 19363 10011 19369
rect 9953 19329 9965 19363
rect 9999 19329 10011 19363
rect 9953 19323 10011 19329
rect 12805 19363 12863 19369
rect 12805 19329 12817 19363
rect 12851 19360 12863 19363
rect 12851 19332 13768 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 7883 19264 9444 19292
rect 7883 19261 7895 19264
rect 7837 19255 7895 19261
rect 9306 19224 9312 19236
rect 7576 19196 9312 19224
rect 7377 19187 7435 19193
rect 9306 19184 9312 19196
rect 9364 19184 9370 19236
rect 1578 19116 1584 19168
rect 1636 19156 1642 19168
rect 1673 19159 1731 19165
rect 1673 19156 1685 19159
rect 1636 19128 1685 19156
rect 1636 19116 1642 19128
rect 1673 19125 1685 19128
rect 1719 19125 1731 19159
rect 1673 19119 1731 19125
rect 2130 19116 2136 19168
rect 2188 19156 2194 19168
rect 2777 19159 2835 19165
rect 2777 19156 2789 19159
rect 2188 19128 2789 19156
rect 2188 19116 2194 19128
rect 2777 19125 2789 19128
rect 2823 19125 2835 19159
rect 2777 19119 2835 19125
rect 4433 19159 4491 19165
rect 4433 19125 4445 19159
rect 4479 19156 4491 19159
rect 4522 19156 4528 19168
rect 4479 19128 4528 19156
rect 4479 19125 4491 19128
rect 4433 19119 4491 19125
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 4890 19156 4896 19168
rect 4851 19128 4896 19156
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 4982 19116 4988 19168
rect 5040 19156 5046 19168
rect 6457 19159 6515 19165
rect 6457 19156 6469 19159
rect 5040 19128 6469 19156
rect 5040 19116 5046 19128
rect 6457 19125 6469 19128
rect 6503 19125 6515 19159
rect 6457 19119 6515 19125
rect 6638 19116 6644 19168
rect 6696 19156 6702 19168
rect 7009 19159 7067 19165
rect 7009 19156 7021 19159
rect 6696 19128 7021 19156
rect 6696 19116 6702 19128
rect 7009 19125 7021 19128
rect 7055 19125 7067 19159
rect 7009 19119 7067 19125
rect 7929 19159 7987 19165
rect 7929 19125 7941 19159
rect 7975 19156 7987 19159
rect 8202 19156 8208 19168
rect 7975 19128 8208 19156
rect 7975 19125 7987 19128
rect 7929 19119 7987 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 8297 19159 8355 19165
rect 8297 19125 8309 19159
rect 8343 19156 8355 19159
rect 8754 19156 8760 19168
rect 8343 19128 8760 19156
rect 8343 19125 8355 19128
rect 8297 19119 8355 19125
rect 8754 19116 8760 19128
rect 8812 19116 8818 19168
rect 8938 19156 8944 19168
rect 8899 19128 8944 19156
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 9416 19156 9444 19264
rect 9490 19252 9496 19304
rect 9548 19292 9554 19304
rect 11146 19292 11152 19304
rect 9548 19264 11152 19292
rect 9548 19252 9554 19264
rect 11146 19252 11152 19264
rect 11204 19252 11210 19304
rect 11609 19295 11667 19301
rect 11609 19261 11621 19295
rect 11655 19292 11667 19295
rect 12066 19292 12072 19304
rect 11655 19264 12072 19292
rect 11655 19261 11667 19264
rect 11609 19255 11667 19261
rect 12066 19252 12072 19264
rect 12124 19252 12130 19304
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19292 12955 19295
rect 12986 19292 12992 19304
rect 12943 19264 12992 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 13630 19292 13636 19304
rect 13591 19264 13636 19292
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 13740 19292 13768 19332
rect 13998 19292 14004 19304
rect 13740 19264 14004 19292
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 14185 19295 14243 19301
rect 14185 19292 14197 19295
rect 14148 19264 14197 19292
rect 14148 19252 14154 19264
rect 14185 19261 14197 19264
rect 14231 19261 14243 19295
rect 14185 19255 14243 19261
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14737 19295 14795 19301
rect 14737 19292 14749 19295
rect 14332 19264 14749 19292
rect 14332 19252 14338 19264
rect 14737 19261 14749 19264
rect 14783 19261 14795 19295
rect 14737 19255 14795 19261
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19261 15347 19295
rect 15838 19292 15844 19304
rect 15799 19264 15844 19292
rect 15289 19255 15347 19261
rect 9674 19184 9680 19236
rect 9732 19224 9738 19236
rect 10134 19224 10140 19236
rect 9732 19196 10140 19224
rect 9732 19184 9738 19196
rect 10134 19184 10140 19196
rect 10192 19233 10198 19236
rect 10192 19227 10256 19233
rect 10192 19193 10210 19227
rect 10244 19193 10256 19227
rect 11882 19224 11888 19236
rect 11843 19196 11888 19224
rect 10192 19187 10256 19193
rect 10192 19184 10198 19187
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 13173 19227 13231 19233
rect 13173 19193 13185 19227
rect 13219 19224 13231 19227
rect 15304 19224 15332 19255
rect 15838 19252 15844 19264
rect 15896 19252 15902 19304
rect 16390 19292 16396 19304
rect 16351 19264 16396 19292
rect 16390 19252 16396 19264
rect 16448 19252 16454 19304
rect 16960 19301 16988 19400
rect 17236 19369 17264 19400
rect 18690 19388 18696 19400
rect 18748 19388 18754 19440
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 16945 19295 17003 19301
rect 16945 19261 16957 19295
rect 16991 19261 17003 19295
rect 17586 19292 17592 19304
rect 16945 19255 17003 19261
rect 17052 19264 17592 19292
rect 17052 19224 17080 19264
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 17770 19252 17776 19304
rect 17828 19292 17834 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17828 19264 18061 19292
rect 17828 19252 17834 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 18785 19295 18843 19301
rect 18785 19292 18797 19295
rect 18196 19264 18797 19292
rect 18196 19252 18202 19264
rect 18785 19261 18797 19264
rect 18831 19292 18843 19295
rect 19794 19292 19800 19304
rect 18831 19264 19104 19292
rect 19707 19264 19800 19292
rect 18831 19261 18843 19264
rect 18785 19255 18843 19261
rect 13219 19196 17080 19224
rect 13219 19193 13231 19196
rect 13173 19187 13231 19193
rect 17494 19184 17500 19236
rect 17552 19224 17558 19236
rect 17552 19196 18276 19224
rect 17552 19184 17558 19196
rect 11333 19159 11391 19165
rect 11333 19156 11345 19159
rect 9416 19128 11345 19156
rect 11333 19125 11345 19128
rect 11379 19125 11391 19159
rect 11333 19119 11391 19125
rect 12894 19116 12900 19168
rect 12952 19156 12958 19168
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 12952 19128 13829 19156
rect 12952 19116 12958 19128
rect 13817 19125 13829 19128
rect 13863 19125 13875 19159
rect 13817 19119 13875 19125
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 14369 19159 14427 19165
rect 14369 19156 14381 19159
rect 13964 19128 14381 19156
rect 13964 19116 13970 19128
rect 14369 19125 14381 19128
rect 14415 19125 14427 19159
rect 14369 19119 14427 19125
rect 14921 19159 14979 19165
rect 14921 19125 14933 19159
rect 14967 19156 14979 19159
rect 15010 19156 15016 19168
rect 14967 19128 15016 19156
rect 14967 19125 14979 19128
rect 14921 19119 14979 19125
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 15473 19159 15531 19165
rect 15473 19156 15485 19159
rect 15252 19128 15485 19156
rect 15252 19116 15258 19128
rect 15473 19125 15485 19128
rect 15519 19125 15531 19159
rect 15473 19119 15531 19125
rect 15654 19116 15660 19168
rect 15712 19156 15718 19168
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15712 19128 16037 19156
rect 15712 19116 15718 19128
rect 16025 19125 16037 19128
rect 16071 19125 16083 19159
rect 16025 19119 16083 19125
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 16577 19159 16635 19165
rect 16577 19156 16589 19159
rect 16172 19128 16589 19156
rect 16172 19116 16178 19128
rect 16577 19125 16589 19128
rect 16623 19125 16635 19159
rect 17678 19156 17684 19168
rect 17639 19128 17684 19156
rect 16577 19119 16635 19125
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 18248 19156 18276 19196
rect 18322 19184 18328 19236
rect 18380 19224 18386 19236
rect 18380 19196 18425 19224
rect 18380 19184 18386 19196
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 18248 19128 18981 19156
rect 18969 19125 18981 19128
rect 19015 19125 19027 19159
rect 19076 19156 19104 19264
rect 19794 19252 19800 19264
rect 19852 19292 19858 19304
rect 22094 19292 22100 19304
rect 19852 19264 22100 19292
rect 19852 19252 19858 19264
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 19334 19224 19340 19236
rect 19295 19196 19340 19224
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 19610 19184 19616 19236
rect 19668 19224 19674 19236
rect 20441 19227 20499 19233
rect 20441 19224 20453 19227
rect 19668 19196 20453 19224
rect 19668 19184 19674 19196
rect 20441 19193 20453 19196
rect 20487 19193 20499 19227
rect 20441 19187 20499 19193
rect 20806 19156 20812 19168
rect 19076 19128 20812 19156
rect 18969 19119 19027 19125
rect 20806 19116 20812 19128
rect 20864 19116 20870 19168
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 20956 19128 21001 19156
rect 20956 19116 20962 19128
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 2774 18952 2780 18964
rect 1627 18924 2780 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 2774 18912 2780 18924
rect 2832 18912 2838 18964
rect 2866 18912 2872 18964
rect 2924 18952 2930 18964
rect 4525 18955 4583 18961
rect 2924 18924 2969 18952
rect 2924 18912 2930 18924
rect 4525 18921 4537 18955
rect 4571 18952 4583 18955
rect 5166 18952 5172 18964
rect 4571 18924 5172 18952
rect 4571 18921 4583 18924
rect 4525 18915 4583 18921
rect 5166 18912 5172 18924
rect 5224 18912 5230 18964
rect 6730 18952 6736 18964
rect 6691 18924 6736 18952
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 10318 18952 10324 18964
rect 6840 18924 10324 18952
rect 2222 18884 2228 18896
rect 2183 18856 2228 18884
rect 2222 18844 2228 18856
rect 2280 18844 2286 18896
rect 2792 18856 5764 18884
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 1949 18819 2007 18825
rect 1949 18785 1961 18819
rect 1995 18816 2007 18819
rect 2682 18816 2688 18828
rect 1995 18788 2688 18816
rect 1995 18785 2007 18788
rect 1949 18779 2007 18785
rect 2682 18776 2688 18788
rect 2740 18776 2746 18828
rect 198 18708 204 18760
rect 256 18748 262 18760
rect 2792 18748 2820 18856
rect 3237 18819 3295 18825
rect 3237 18785 3249 18819
rect 3283 18785 3295 18819
rect 3237 18779 3295 18785
rect 3329 18819 3387 18825
rect 3329 18785 3341 18819
rect 3375 18816 3387 18819
rect 4433 18819 4491 18825
rect 3375 18788 4108 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 256 18720 2820 18748
rect 256 18708 262 18720
rect 3050 18708 3056 18760
rect 3108 18748 3114 18760
rect 3252 18748 3280 18779
rect 3108 18720 3280 18748
rect 3513 18751 3571 18757
rect 3108 18708 3114 18720
rect 3513 18717 3525 18751
rect 3559 18717 3571 18751
rect 3513 18711 3571 18717
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 2682 18612 2688 18624
rect 1544 18584 2688 18612
rect 1544 18572 1550 18584
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 2777 18615 2835 18621
rect 2777 18581 2789 18615
rect 2823 18612 2835 18615
rect 3234 18612 3240 18624
rect 2823 18584 3240 18612
rect 2823 18581 2835 18584
rect 2777 18575 2835 18581
rect 3234 18572 3240 18584
rect 3292 18612 3298 18624
rect 3528 18612 3556 18711
rect 4080 18692 4108 18788
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 5074 18816 5080 18828
rect 4479 18788 5080 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 5626 18825 5632 18828
rect 5620 18816 5632 18825
rect 5587 18788 5632 18816
rect 5620 18779 5632 18788
rect 5626 18776 5632 18779
rect 5684 18776 5690 18828
rect 5736 18816 5764 18856
rect 5810 18844 5816 18896
rect 5868 18884 5874 18896
rect 6840 18884 6868 18924
rect 10318 18912 10324 18924
rect 10376 18952 10382 18964
rect 13630 18952 13636 18964
rect 10376 18924 12020 18952
rect 13543 18924 13636 18952
rect 10376 18912 10382 18924
rect 5868 18856 6868 18884
rect 6912 18856 7972 18884
rect 5868 18844 5874 18856
rect 6912 18816 6940 18856
rect 5736 18788 6940 18816
rect 7650 18776 7656 18828
rect 7708 18816 7714 18828
rect 7817 18819 7875 18825
rect 7817 18816 7829 18819
rect 7708 18788 7829 18816
rect 7708 18776 7714 18788
rect 7817 18785 7829 18788
rect 7863 18785 7875 18819
rect 7944 18816 7972 18856
rect 8018 18844 8024 18896
rect 8076 18884 8082 18896
rect 8754 18884 8760 18896
rect 8076 18856 8760 18884
rect 8076 18844 8082 18856
rect 8754 18844 8760 18856
rect 8812 18844 8818 18896
rect 9306 18884 9312 18896
rect 9267 18856 9312 18884
rect 9306 18844 9312 18856
rect 9364 18844 9370 18896
rect 9858 18844 9864 18896
rect 9916 18884 9922 18896
rect 10106 18887 10164 18893
rect 10106 18884 10118 18887
rect 9916 18856 10118 18884
rect 9916 18844 9922 18856
rect 10106 18853 10118 18856
rect 10152 18884 10164 18887
rect 10962 18884 10968 18896
rect 10152 18856 10968 18884
rect 10152 18853 10164 18856
rect 10106 18847 10164 18853
rect 10962 18844 10968 18856
rect 11020 18884 11026 18896
rect 11517 18887 11575 18893
rect 11517 18884 11529 18887
rect 11020 18856 11529 18884
rect 11020 18844 11026 18856
rect 11517 18853 11529 18856
rect 11563 18853 11575 18887
rect 11517 18847 11575 18853
rect 10502 18816 10508 18828
rect 7944 18788 10508 18816
rect 7817 18779 7875 18785
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 11606 18776 11612 18828
rect 11664 18816 11670 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11664 18788 11805 18816
rect 11664 18776 11670 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 11992 18816 12020 18924
rect 13556 18893 13584 18924
rect 13630 18912 13636 18924
rect 13688 18952 13694 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 13688 18924 19533 18952
rect 13688 18912 13694 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 19521 18915 19579 18921
rect 12069 18887 12127 18893
rect 12069 18853 12081 18887
rect 12115 18884 12127 18887
rect 13541 18887 13599 18893
rect 12115 18856 13492 18884
rect 12115 18853 12127 18856
rect 12069 18847 12127 18853
rect 12158 18816 12164 18828
rect 11992 18788 12164 18816
rect 11793 18779 11851 18785
rect 12158 18776 12164 18788
rect 12216 18776 12222 18828
rect 12529 18819 12587 18825
rect 12529 18785 12541 18819
rect 12575 18816 12587 18819
rect 12894 18816 12900 18828
rect 12575 18788 12900 18816
rect 12575 18785 12587 18788
rect 12529 18779 12587 18785
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 13262 18816 13268 18828
rect 13223 18788 13268 18816
rect 13262 18776 13268 18788
rect 13320 18776 13326 18828
rect 13464 18816 13492 18856
rect 13541 18853 13553 18887
rect 13587 18853 13599 18887
rect 13541 18847 13599 18853
rect 13998 18844 14004 18896
rect 14056 18884 14062 18896
rect 14274 18884 14280 18896
rect 14056 18856 14280 18884
rect 14056 18844 14062 18856
rect 14274 18844 14280 18856
rect 14332 18844 14338 18896
rect 15565 18887 15623 18893
rect 15565 18853 15577 18887
rect 15611 18884 15623 18887
rect 15838 18884 15844 18896
rect 15611 18856 15844 18884
rect 15611 18853 15623 18856
rect 15565 18847 15623 18853
rect 15838 18844 15844 18856
rect 15896 18884 15902 18896
rect 20257 18887 20315 18893
rect 20257 18884 20269 18887
rect 15896 18856 20269 18884
rect 15896 18844 15902 18856
rect 20257 18853 20269 18856
rect 20303 18853 20315 18887
rect 20257 18847 20315 18853
rect 14090 18816 14096 18828
rect 13464 18788 14096 18816
rect 14090 18776 14096 18788
rect 14148 18776 14154 18828
rect 15289 18819 15347 18825
rect 15289 18785 15301 18819
rect 15335 18816 15347 18819
rect 15470 18816 15476 18828
rect 15335 18788 15476 18816
rect 15335 18785 15347 18788
rect 15289 18779 15347 18785
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 16025 18819 16083 18825
rect 16025 18785 16037 18819
rect 16071 18816 16083 18819
rect 16482 18816 16488 18828
rect 16071 18788 16488 18816
rect 16071 18785 16083 18788
rect 16025 18779 16083 18785
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 16758 18816 16764 18828
rect 16719 18788 16764 18816
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18816 17739 18819
rect 17862 18816 17868 18828
rect 17727 18788 17868 18816
rect 17727 18785 17739 18788
rect 17681 18779 17739 18785
rect 17862 18776 17868 18788
rect 17920 18776 17926 18828
rect 17957 18819 18015 18825
rect 17957 18785 17969 18819
rect 18003 18816 18015 18819
rect 18138 18816 18144 18828
rect 18003 18788 18144 18816
rect 18003 18785 18015 18788
rect 17957 18779 18015 18785
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 18414 18816 18420 18828
rect 18375 18788 18420 18816
rect 18414 18776 18420 18788
rect 18472 18776 18478 18828
rect 20625 18819 20683 18825
rect 20625 18816 20637 18819
rect 18524 18788 20637 18816
rect 4522 18708 4528 18760
rect 4580 18748 4586 18760
rect 4709 18751 4767 18757
rect 4709 18748 4721 18751
rect 4580 18720 4721 18748
rect 4580 18708 4586 18720
rect 4709 18717 4721 18720
rect 4755 18748 4767 18751
rect 4798 18748 4804 18760
rect 4755 18720 4804 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 5350 18748 5356 18760
rect 5311 18720 5356 18748
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 7374 18748 7380 18760
rect 7147 18720 7380 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 7558 18708 7564 18760
rect 7616 18748 7622 18760
rect 7616 18720 7661 18748
rect 7616 18708 7622 18720
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9640 18720 9873 18748
rect 9640 18708 9646 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 12805 18751 12863 18757
rect 12805 18717 12817 18751
rect 12851 18748 12863 18751
rect 13354 18748 13360 18760
rect 12851 18720 13360 18748
rect 12851 18717 12863 18720
rect 12805 18711 12863 18717
rect 13354 18708 13360 18720
rect 13412 18748 13418 18760
rect 16114 18748 16120 18760
rect 13412 18720 16120 18748
rect 13412 18708 13418 18720
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 16301 18751 16359 18757
rect 16301 18717 16313 18751
rect 16347 18748 16359 18751
rect 16390 18748 16396 18760
rect 16347 18720 16396 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 4062 18680 4068 18692
rect 4023 18652 4068 18680
rect 4062 18640 4068 18652
rect 4120 18640 4126 18692
rect 10870 18640 10876 18692
rect 10928 18680 10934 18692
rect 16316 18680 16344 18711
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 16574 18708 16580 18760
rect 16632 18748 16638 18760
rect 17037 18751 17095 18757
rect 17037 18748 17049 18751
rect 16632 18720 17049 18748
rect 16632 18708 16638 18720
rect 17037 18717 17049 18720
rect 17083 18748 17095 18751
rect 18524 18748 18552 18788
rect 20625 18785 20637 18788
rect 20671 18785 20683 18819
rect 20625 18779 20683 18785
rect 17083 18720 18552 18748
rect 18693 18751 18751 18757
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 18693 18717 18705 18751
rect 18739 18748 18751 18751
rect 18966 18748 18972 18760
rect 18739 18720 18972 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 18966 18708 18972 18720
rect 19024 18708 19030 18760
rect 19150 18748 19156 18760
rect 19111 18720 19156 18748
rect 19150 18708 19156 18720
rect 19208 18708 19214 18760
rect 20438 18680 20444 18692
rect 10928 18652 15700 18680
rect 16316 18652 20444 18680
rect 10928 18640 10934 18652
rect 3970 18612 3976 18624
rect 3292 18584 3976 18612
rect 3292 18572 3298 18584
rect 3970 18572 3976 18584
rect 4028 18572 4034 18624
rect 5261 18615 5319 18621
rect 5261 18581 5273 18615
rect 5307 18612 5319 18615
rect 5718 18612 5724 18624
rect 5307 18584 5724 18612
rect 5307 18581 5319 18584
rect 5261 18575 5319 18581
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 8202 18572 8208 18624
rect 8260 18612 8266 18624
rect 8941 18615 8999 18621
rect 8941 18612 8953 18615
rect 8260 18584 8953 18612
rect 8260 18572 8266 18584
rect 8941 18581 8953 18584
rect 8987 18581 8999 18615
rect 8941 18575 8999 18581
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 11241 18615 11299 18621
rect 11241 18612 11253 18615
rect 9732 18584 11253 18612
rect 9732 18572 9738 18584
rect 11241 18581 11253 18584
rect 11287 18581 11299 18615
rect 13998 18612 14004 18624
rect 13959 18584 14004 18612
rect 11241 18575 11299 18581
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 14461 18615 14519 18621
rect 14461 18581 14473 18615
rect 14507 18612 14519 18615
rect 15010 18612 15016 18624
rect 14507 18584 15016 18612
rect 14507 18581 14519 18584
rect 14461 18575 14519 18581
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15105 18615 15163 18621
rect 15105 18581 15117 18615
rect 15151 18612 15163 18615
rect 15562 18612 15568 18624
rect 15151 18584 15568 18612
rect 15151 18581 15163 18584
rect 15105 18575 15163 18581
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15672 18612 15700 18652
rect 20438 18640 20444 18652
rect 20496 18640 20502 18692
rect 16666 18612 16672 18624
rect 15672 18584 16672 18612
rect 16666 18572 16672 18584
rect 16724 18572 16730 18624
rect 16850 18572 16856 18624
rect 16908 18612 16914 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 16908 18584 17509 18612
rect 16908 18572 16914 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 17586 18572 17592 18624
rect 17644 18612 17650 18624
rect 19889 18615 19947 18621
rect 19889 18612 19901 18615
rect 17644 18584 19901 18612
rect 17644 18572 17650 18584
rect 19889 18581 19901 18584
rect 19935 18581 19947 18615
rect 19889 18575 19947 18581
rect 19978 18572 19984 18624
rect 20036 18612 20042 18624
rect 21085 18615 21143 18621
rect 21085 18612 21097 18615
rect 20036 18584 21097 18612
rect 20036 18572 20042 18584
rect 21085 18581 21097 18584
rect 21131 18581 21143 18615
rect 21085 18575 21143 18581
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 2593 18411 2651 18417
rect 2593 18377 2605 18411
rect 2639 18408 2651 18411
rect 3050 18408 3056 18420
rect 2639 18380 3056 18408
rect 2639 18377 2651 18380
rect 2593 18371 2651 18377
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 4065 18411 4123 18417
rect 4065 18408 4077 18411
rect 4028 18380 4077 18408
rect 4028 18368 4034 18380
rect 4065 18377 4077 18380
rect 4111 18377 4123 18411
rect 4065 18371 4123 18377
rect 4985 18411 5043 18417
rect 4985 18377 4997 18411
rect 5031 18408 5043 18411
rect 5166 18408 5172 18420
rect 5031 18380 5172 18408
rect 5031 18377 5043 18380
rect 4985 18371 5043 18377
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 5537 18411 5595 18417
rect 5537 18377 5549 18411
rect 5583 18408 5595 18411
rect 6270 18408 6276 18420
rect 5583 18380 6276 18408
rect 5583 18377 5595 18380
rect 5537 18371 5595 18377
rect 6270 18368 6276 18380
rect 6328 18368 6334 18420
rect 7377 18411 7435 18417
rect 7377 18377 7389 18411
rect 7423 18408 7435 18411
rect 7561 18411 7619 18417
rect 7561 18408 7573 18411
rect 7423 18380 7573 18408
rect 7423 18377 7435 18380
rect 7377 18371 7435 18377
rect 7561 18377 7573 18380
rect 7607 18408 7619 18411
rect 10870 18408 10876 18420
rect 7607 18380 10876 18408
rect 7607 18377 7619 18380
rect 7561 18371 7619 18377
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 11149 18411 11207 18417
rect 11149 18408 11161 18411
rect 11020 18380 11161 18408
rect 11020 18368 11026 18380
rect 11149 18377 11161 18380
rect 11195 18377 11207 18411
rect 11149 18371 11207 18377
rect 12437 18411 12495 18417
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 13265 18411 13323 18417
rect 13265 18408 13277 18411
rect 12483 18380 13277 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 13265 18377 13277 18380
rect 13311 18377 13323 18411
rect 13265 18371 13323 18377
rect 13722 18368 13728 18420
rect 13780 18408 13786 18420
rect 14829 18411 14887 18417
rect 14829 18408 14841 18411
rect 13780 18380 14841 18408
rect 13780 18368 13786 18380
rect 14829 18377 14841 18380
rect 14875 18408 14887 18411
rect 15378 18408 15384 18420
rect 14875 18380 15384 18408
rect 14875 18377 14887 18380
rect 14829 18371 14887 18377
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 15488 18380 18061 18408
rect 2682 18300 2688 18352
rect 2740 18300 2746 18352
rect 3694 18300 3700 18352
rect 3752 18340 3758 18352
rect 3752 18312 5028 18340
rect 3752 18300 3758 18312
rect 1946 18232 1952 18284
rect 2004 18272 2010 18284
rect 2222 18272 2228 18284
rect 2004 18244 2228 18272
rect 2004 18232 2010 18244
rect 2222 18232 2228 18244
rect 2280 18232 2286 18284
rect 2700 18272 2728 18300
rect 2700 18244 2820 18272
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2682 18204 2688 18216
rect 2643 18176 2688 18204
rect 2682 18164 2688 18176
rect 2740 18164 2746 18216
rect 2792 18204 2820 18244
rect 4246 18232 4252 18284
rect 4304 18272 4310 18284
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 4304 18244 4445 18272
rect 4304 18232 4310 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 5000 18272 5028 18312
rect 5074 18300 5080 18352
rect 5132 18340 5138 18352
rect 5353 18343 5411 18349
rect 5353 18340 5365 18343
rect 5132 18312 5365 18340
rect 5132 18300 5138 18312
rect 5353 18309 5365 18312
rect 5399 18340 5411 18343
rect 5399 18312 7788 18340
rect 5399 18309 5411 18312
rect 5353 18303 5411 18309
rect 5442 18272 5448 18284
rect 5000 18244 5448 18272
rect 4433 18235 4491 18241
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 5902 18232 5908 18284
rect 5960 18272 5966 18284
rect 6181 18275 6239 18281
rect 6181 18272 6193 18275
rect 5960 18244 6193 18272
rect 5960 18232 5966 18244
rect 6181 18241 6193 18244
rect 6227 18272 6239 18275
rect 6638 18272 6644 18284
rect 6227 18244 6644 18272
rect 6227 18241 6239 18244
rect 6181 18235 6239 18241
rect 6638 18232 6644 18244
rect 6696 18232 6702 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 6840 18244 7389 18272
rect 5534 18204 5540 18216
rect 2792 18176 5540 18204
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 6840 18213 6868 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 7760 18272 7788 18312
rect 8478 18300 8484 18352
rect 8536 18340 8542 18352
rect 8757 18343 8815 18349
rect 8757 18340 8769 18343
rect 8536 18312 8769 18340
rect 8536 18300 8542 18312
rect 8757 18309 8769 18312
rect 8803 18340 8815 18343
rect 9398 18340 9404 18352
rect 8803 18312 9404 18340
rect 8803 18309 8815 18312
rect 8757 18303 8815 18309
rect 9398 18300 9404 18312
rect 9456 18300 9462 18352
rect 10778 18300 10784 18352
rect 10836 18340 10842 18352
rect 12342 18340 12348 18352
rect 10836 18312 12348 18340
rect 10836 18300 10842 18312
rect 12342 18300 12348 18312
rect 12400 18300 12406 18352
rect 13814 18340 13820 18352
rect 13096 18312 13820 18340
rect 8018 18272 8024 18284
rect 7760 18244 8024 18272
rect 7377 18235 7435 18241
rect 8018 18232 8024 18244
rect 8076 18232 8082 18284
rect 8202 18272 8208 18284
rect 8163 18244 8208 18272
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 9309 18275 9367 18281
rect 9309 18272 9321 18275
rect 8444 18244 9321 18272
rect 8444 18232 8450 18244
rect 9309 18241 9321 18244
rect 9355 18272 9367 18275
rect 9674 18272 9680 18284
rect 9355 18244 9680 18272
rect 9355 18241 9367 18244
rect 9309 18235 9367 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 10870 18232 10876 18284
rect 10928 18272 10934 18284
rect 13096 18281 13124 18312
rect 13814 18300 13820 18312
rect 13872 18340 13878 18352
rect 15010 18340 15016 18352
rect 13872 18312 15016 18340
rect 13872 18300 13878 18312
rect 15010 18300 15016 18312
rect 15068 18300 15074 18352
rect 15488 18340 15516 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 18049 18371 18107 18377
rect 18325 18411 18383 18417
rect 18325 18377 18337 18411
rect 18371 18408 18383 18411
rect 18874 18408 18880 18420
rect 18371 18380 18880 18408
rect 18371 18377 18383 18380
rect 18325 18371 18383 18377
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 18969 18411 19027 18417
rect 18969 18377 18981 18411
rect 19015 18408 19027 18411
rect 19245 18411 19303 18417
rect 19245 18408 19257 18411
rect 19015 18380 19257 18408
rect 19015 18377 19027 18380
rect 18969 18371 19027 18377
rect 19245 18377 19257 18380
rect 19291 18377 19303 18411
rect 19426 18408 19432 18420
rect 19387 18380 19432 18408
rect 19245 18371 19303 18377
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 18693 18343 18751 18349
rect 18693 18340 18705 18343
rect 15120 18312 15516 18340
rect 16684 18312 18705 18340
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 10928 18244 12173 18272
rect 10928 18232 10934 18244
rect 12161 18241 12173 18244
rect 12207 18272 12219 18275
rect 12897 18275 12955 18281
rect 12897 18272 12909 18275
rect 12207 18244 12909 18272
rect 12207 18241 12219 18244
rect 12161 18235 12219 18241
rect 12897 18241 12909 18244
rect 12943 18241 12955 18275
rect 12897 18235 12955 18241
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18241 13139 18275
rect 13998 18272 14004 18284
rect 13959 18244 14004 18272
rect 13081 18235 13139 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 15120 18272 15148 18312
rect 14476 18244 15148 18272
rect 5997 18207 6055 18213
rect 5997 18173 6009 18207
rect 6043 18204 6055 18207
rect 6825 18207 6883 18213
rect 6043 18176 6132 18204
rect 6043 18173 6055 18176
rect 5997 18167 6055 18173
rect 6104 18148 6132 18176
rect 6825 18173 6837 18207
rect 6871 18173 6883 18207
rect 8573 18207 8631 18213
rect 8573 18204 8585 18207
rect 6825 18167 6883 18173
rect 7944 18176 8248 18204
rect 1673 18139 1731 18145
rect 1673 18105 1685 18139
rect 1719 18136 1731 18139
rect 2952 18139 3010 18145
rect 1719 18108 2176 18136
rect 1719 18105 1731 18108
rect 1673 18099 1731 18105
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2148 18068 2176 18108
rect 2952 18105 2964 18139
rect 2998 18105 3010 18139
rect 2952 18099 3010 18105
rect 2967 18068 2995 18099
rect 4062 18096 4068 18148
rect 4120 18136 4126 18148
rect 4120 18108 6040 18136
rect 4120 18096 4126 18108
rect 4246 18068 4252 18080
rect 2148 18040 4252 18068
rect 4246 18028 4252 18040
rect 4304 18068 4310 18080
rect 4798 18068 4804 18080
rect 4304 18040 4804 18068
rect 4304 18028 4310 18040
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 5166 18028 5172 18080
rect 5224 18068 5230 18080
rect 5350 18068 5356 18080
rect 5224 18040 5356 18068
rect 5224 18028 5230 18040
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 5810 18028 5816 18080
rect 5868 18068 5874 18080
rect 5905 18071 5963 18077
rect 5905 18068 5917 18071
rect 5868 18040 5917 18068
rect 5868 18028 5874 18040
rect 5905 18037 5917 18040
rect 5951 18037 5963 18071
rect 6012 18068 6040 18108
rect 6086 18096 6092 18148
rect 6144 18136 6150 18148
rect 6549 18139 6607 18145
rect 6549 18136 6561 18139
rect 6144 18108 6561 18136
rect 6144 18096 6150 18108
rect 6549 18105 6561 18108
rect 6595 18105 6607 18139
rect 6549 18099 6607 18105
rect 7101 18139 7159 18145
rect 7101 18105 7113 18139
rect 7147 18136 7159 18139
rect 7190 18136 7196 18148
rect 7147 18108 7196 18136
rect 7147 18105 7159 18108
rect 7101 18099 7159 18105
rect 7116 18068 7144 18099
rect 7190 18096 7196 18108
rect 7248 18096 7254 18148
rect 7374 18096 7380 18148
rect 7432 18136 7438 18148
rect 7944 18145 7972 18176
rect 7929 18139 7987 18145
rect 7929 18136 7941 18139
rect 7432 18108 7941 18136
rect 7432 18096 7438 18108
rect 7929 18105 7941 18108
rect 7975 18105 7987 18139
rect 7929 18099 7987 18105
rect 8021 18139 8079 18145
rect 8021 18105 8033 18139
rect 8067 18136 8079 18139
rect 8110 18136 8116 18148
rect 8067 18108 8116 18136
rect 8067 18105 8079 18108
rect 8021 18099 8079 18105
rect 8110 18096 8116 18108
rect 8168 18096 8174 18148
rect 8220 18136 8248 18176
rect 8404 18176 8585 18204
rect 8404 18136 8432 18176
rect 8573 18173 8585 18176
rect 8619 18173 8631 18207
rect 9122 18204 9128 18216
rect 9083 18176 9128 18204
rect 8573 18167 8631 18173
rect 9122 18164 9128 18176
rect 9180 18164 9186 18216
rect 9582 18164 9588 18216
rect 9640 18204 9646 18216
rect 9769 18207 9827 18213
rect 9769 18204 9781 18207
rect 9640 18176 9781 18204
rect 9640 18164 9646 18176
rect 9769 18173 9781 18176
rect 9815 18173 9827 18207
rect 14366 18204 14372 18216
rect 9769 18167 9827 18173
rect 9968 18176 14372 18204
rect 8220 18108 8432 18136
rect 8938 18096 8944 18148
rect 8996 18136 9002 18148
rect 9217 18139 9275 18145
rect 9217 18136 9229 18139
rect 8996 18108 9229 18136
rect 8996 18096 9002 18108
rect 9217 18105 9229 18108
rect 9263 18136 9275 18139
rect 9968 18136 9996 18176
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 9263 18108 9996 18136
rect 10036 18139 10094 18145
rect 9263 18105 9275 18108
rect 9217 18099 9275 18105
rect 10036 18105 10048 18139
rect 10082 18136 10094 18139
rect 11885 18139 11943 18145
rect 10082 18108 11008 18136
rect 10082 18105 10094 18108
rect 10036 18099 10094 18105
rect 10980 18080 11008 18108
rect 11885 18105 11897 18139
rect 11931 18136 11943 18139
rect 13265 18139 13323 18145
rect 11931 18108 12848 18136
rect 11931 18105 11943 18108
rect 11885 18099 11943 18105
rect 12820 18080 12848 18108
rect 13265 18105 13277 18139
rect 13311 18136 13323 18139
rect 13817 18139 13875 18145
rect 13817 18136 13829 18139
rect 13311 18108 13829 18136
rect 13311 18105 13323 18108
rect 13265 18099 13323 18105
rect 13817 18105 13829 18108
rect 13863 18136 13875 18139
rect 14476 18136 14504 18244
rect 15378 18232 15384 18284
rect 15436 18272 15442 18284
rect 15473 18275 15531 18281
rect 15473 18272 15485 18275
rect 15436 18244 15485 18272
rect 15436 18232 15442 18244
rect 15473 18241 15485 18244
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 15562 18232 15568 18284
rect 15620 18272 15626 18284
rect 16684 18281 16712 18312
rect 18693 18309 18705 18312
rect 18739 18309 18751 18343
rect 18693 18303 18751 18309
rect 18782 18300 18788 18352
rect 18840 18340 18846 18352
rect 20533 18343 20591 18349
rect 20533 18340 20545 18343
rect 18840 18312 20545 18340
rect 18840 18300 18846 18312
rect 20533 18309 20545 18312
rect 20579 18309 20591 18343
rect 20533 18303 20591 18309
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 15620 18244 15669 18272
rect 15620 18232 15626 18244
rect 15657 18241 15669 18244
rect 15703 18272 15715 18275
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 15703 18244 16681 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 17402 18272 17408 18284
rect 16669 18235 16727 18241
rect 17144 18244 17408 18272
rect 14550 18164 14556 18216
rect 14608 18204 14614 18216
rect 16022 18204 16028 18216
rect 14608 18176 16028 18204
rect 14608 18164 14614 18176
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 16114 18164 16120 18216
rect 16172 18204 16178 18216
rect 17144 18213 17172 18244
rect 17402 18232 17408 18244
rect 17460 18272 17466 18284
rect 20993 18275 21051 18281
rect 20993 18272 21005 18275
rect 17460 18244 21005 18272
rect 17460 18232 17466 18244
rect 20993 18241 21005 18244
rect 21039 18241 21051 18275
rect 20993 18235 21051 18241
rect 17129 18207 17187 18213
rect 16172 18176 16611 18204
rect 16172 18164 16178 18176
rect 13863 18108 14504 18136
rect 14568 18108 15231 18136
rect 13863 18105 13875 18108
rect 13817 18099 13875 18105
rect 6012 18040 7144 18068
rect 5905 18031 5963 18037
rect 7558 18028 7564 18080
rect 7616 18068 7622 18080
rect 9582 18068 9588 18080
rect 7616 18040 9588 18068
rect 7616 18028 7622 18040
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 10870 18068 10876 18080
rect 9732 18040 10876 18068
rect 9732 18028 9738 18040
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 10962 18028 10968 18080
rect 11020 18068 11026 18080
rect 11425 18071 11483 18077
rect 11425 18068 11437 18071
rect 11020 18040 11437 18068
rect 11020 18028 11026 18040
rect 11425 18037 11437 18040
rect 11471 18037 11483 18071
rect 12802 18068 12808 18080
rect 12763 18040 12808 18068
rect 11425 18031 11483 18037
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 12894 18028 12900 18080
rect 12952 18068 12958 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 12952 18040 13461 18068
rect 12952 18028 12958 18040
rect 13449 18037 13461 18040
rect 13495 18068 13507 18071
rect 13722 18068 13728 18080
rect 13495 18040 13728 18068
rect 13495 18037 13507 18040
rect 13449 18031 13507 18037
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 14458 18068 14464 18080
rect 13964 18040 14009 18068
rect 14419 18040 14464 18068
rect 13964 18028 13970 18040
rect 14458 18028 14464 18040
rect 14516 18068 14522 18080
rect 14568 18068 14596 18108
rect 14516 18040 14596 18068
rect 15013 18071 15071 18077
rect 14516 18028 14522 18040
rect 15013 18037 15025 18071
rect 15059 18068 15071 18071
rect 15102 18068 15108 18080
rect 15059 18040 15108 18068
rect 15059 18037 15071 18040
rect 15013 18031 15071 18037
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15203 18068 15231 18108
rect 15286 18096 15292 18148
rect 15344 18136 15350 18148
rect 16482 18136 16488 18148
rect 15344 18108 16488 18136
rect 15344 18096 15350 18108
rect 16482 18096 16488 18108
rect 16540 18096 16546 18148
rect 15378 18068 15384 18080
rect 15203 18040 15384 18068
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 16022 18068 16028 18080
rect 15983 18040 16028 18068
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 16393 18071 16451 18077
rect 16393 18068 16405 18071
rect 16172 18040 16405 18068
rect 16172 18028 16178 18040
rect 16393 18037 16405 18040
rect 16439 18037 16451 18071
rect 16583 18068 16611 18176
rect 17129 18173 17141 18207
rect 17175 18173 17187 18207
rect 17129 18167 17187 18173
rect 18141 18207 18199 18213
rect 18141 18173 18153 18207
rect 18187 18204 18199 18207
rect 18506 18204 18512 18216
rect 18187 18176 18512 18204
rect 18187 18173 18199 18176
rect 18141 18167 18199 18173
rect 18506 18164 18512 18176
rect 18564 18204 18570 18216
rect 18782 18204 18788 18216
rect 18564 18176 18788 18204
rect 18564 18164 18570 18176
rect 18782 18164 18788 18176
rect 18840 18164 18846 18216
rect 19058 18204 19064 18216
rect 19019 18176 19064 18204
rect 19058 18164 19064 18176
rect 19116 18164 19122 18216
rect 19245 18207 19303 18213
rect 19245 18173 19257 18207
rect 19291 18204 19303 18207
rect 19978 18204 19984 18216
rect 19291 18176 19984 18204
rect 19291 18173 19303 18176
rect 19245 18167 19303 18173
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 20898 18164 20904 18216
rect 20956 18204 20962 18216
rect 21634 18204 21640 18216
rect 20956 18176 21640 18204
rect 20956 18164 20962 18176
rect 21634 18164 21640 18176
rect 21692 18164 21698 18216
rect 17310 18096 17316 18148
rect 17368 18136 17374 18148
rect 17405 18139 17463 18145
rect 17405 18136 17417 18139
rect 17368 18108 17417 18136
rect 17368 18096 17374 18108
rect 17405 18105 17417 18108
rect 17451 18105 17463 18139
rect 17405 18099 17463 18105
rect 18049 18139 18107 18145
rect 18049 18105 18061 18139
rect 18095 18136 18107 18139
rect 19702 18136 19708 18148
rect 18095 18108 19708 18136
rect 18095 18105 18107 18108
rect 18049 18099 18107 18105
rect 19702 18096 19708 18108
rect 19760 18096 19766 18148
rect 19886 18096 19892 18148
rect 19944 18136 19950 18148
rect 20254 18136 20260 18148
rect 19944 18108 20260 18136
rect 19944 18096 19950 18108
rect 20254 18096 20260 18108
rect 20312 18096 20318 18148
rect 18969 18071 19027 18077
rect 18969 18068 18981 18071
rect 16583 18040 18981 18068
rect 16393 18031 16451 18037
rect 18969 18037 18981 18040
rect 19015 18037 19027 18071
rect 18969 18031 19027 18037
rect 19242 18028 19248 18080
rect 19300 18068 19306 18080
rect 19797 18071 19855 18077
rect 19797 18068 19809 18071
rect 19300 18040 19809 18068
rect 19300 18028 19306 18040
rect 19797 18037 19809 18040
rect 19843 18037 19855 18071
rect 19797 18031 19855 18037
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 20165 18071 20223 18077
rect 20165 18068 20177 18071
rect 20036 18040 20177 18068
rect 20036 18028 20042 18040
rect 20165 18037 20177 18040
rect 20211 18037 20223 18071
rect 20165 18031 20223 18037
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 2501 17867 2559 17873
rect 2501 17833 2513 17867
rect 2547 17864 2559 17867
rect 2774 17864 2780 17876
rect 2547 17836 2780 17864
rect 2547 17833 2559 17836
rect 2501 17827 2559 17833
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 3108 17836 3433 17864
rect 3108 17824 3114 17836
rect 3421 17833 3433 17836
rect 3467 17833 3479 17867
rect 4246 17864 4252 17876
rect 4207 17836 4252 17864
rect 3421 17827 3479 17833
rect 4246 17824 4252 17836
rect 4304 17824 4310 17876
rect 5626 17824 5632 17876
rect 5684 17824 5690 17876
rect 7558 17824 7564 17876
rect 7616 17864 7622 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7616 17836 7665 17864
rect 7616 17824 7622 17836
rect 7653 17833 7665 17836
rect 7699 17864 7711 17867
rect 8021 17867 8079 17873
rect 8021 17864 8033 17867
rect 7699 17836 8033 17864
rect 7699 17833 7711 17836
rect 7653 17827 7711 17833
rect 8021 17833 8033 17836
rect 8067 17864 8079 17867
rect 8202 17864 8208 17876
rect 8067 17836 8208 17864
rect 8067 17833 8079 17836
rect 8021 17827 8079 17833
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 8386 17864 8392 17876
rect 8347 17836 8392 17864
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 9122 17824 9128 17876
rect 9180 17864 9186 17876
rect 9217 17867 9275 17873
rect 9217 17864 9229 17867
rect 9180 17836 9229 17864
rect 9180 17824 9186 17836
rect 9217 17833 9229 17836
rect 9263 17833 9275 17867
rect 9217 17827 9275 17833
rect 9306 17824 9312 17876
rect 9364 17864 9370 17876
rect 9674 17864 9680 17876
rect 9364 17836 9680 17864
rect 9364 17824 9370 17836
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 10137 17867 10195 17873
rect 10137 17864 10149 17867
rect 9824 17836 10149 17864
rect 9824 17824 9830 17836
rect 10137 17833 10149 17836
rect 10183 17864 10195 17867
rect 10689 17867 10747 17873
rect 10689 17864 10701 17867
rect 10183 17836 10701 17864
rect 10183 17833 10195 17836
rect 10137 17827 10195 17833
rect 10689 17833 10701 17836
rect 10735 17833 10747 17867
rect 10689 17827 10747 17833
rect 11146 17824 11152 17876
rect 11204 17864 11210 17876
rect 12710 17864 12716 17876
rect 11204 17836 12716 17864
rect 11204 17824 11210 17836
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 12802 17824 12808 17876
rect 12860 17864 12866 17876
rect 13633 17867 13691 17873
rect 13633 17864 13645 17867
rect 12860 17836 13645 17864
rect 12860 17824 12866 17836
rect 13633 17833 13645 17836
rect 13679 17833 13691 17867
rect 13633 17827 13691 17833
rect 13906 17824 13912 17876
rect 13964 17864 13970 17876
rect 14185 17867 14243 17873
rect 14185 17864 14197 17867
rect 13964 17836 14197 17864
rect 13964 17824 13970 17836
rect 14185 17833 14197 17836
rect 14231 17864 14243 17867
rect 21085 17867 21143 17873
rect 21085 17864 21097 17867
rect 14231 17836 21097 17864
rect 14231 17833 14243 17836
rect 14185 17827 14243 17833
rect 21085 17833 21097 17836
rect 21131 17833 21143 17867
rect 21085 17827 21143 17833
rect 5528 17799 5586 17805
rect 1780 17768 5488 17796
rect 1780 17737 1808 17768
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17697 2375 17731
rect 2866 17728 2872 17740
rect 2827 17700 2872 17728
rect 2317 17691 2375 17697
rect 1026 17620 1032 17672
rect 1084 17660 1090 17672
rect 2332 17660 2360 17691
rect 2866 17688 2872 17700
rect 2924 17688 2930 17740
rect 5460 17728 5488 17768
rect 5528 17765 5540 17799
rect 5574 17796 5586 17799
rect 5644 17796 5672 17824
rect 5574 17768 5672 17796
rect 5574 17765 5586 17768
rect 5528 17759 5586 17765
rect 6086 17756 6092 17808
rect 6144 17796 6150 17808
rect 14458 17796 14464 17808
rect 6144 17768 14464 17796
rect 6144 17756 6150 17768
rect 14458 17756 14464 17768
rect 14516 17756 14522 17808
rect 16942 17756 16948 17808
rect 17000 17796 17006 17808
rect 17865 17799 17923 17805
rect 17865 17796 17877 17799
rect 17000 17768 17877 17796
rect 17000 17756 17006 17768
rect 17865 17765 17877 17768
rect 17911 17796 17923 17799
rect 20438 17796 20444 17808
rect 17911 17768 20444 17796
rect 17911 17765 17923 17768
rect 17865 17759 17923 17765
rect 20438 17756 20444 17768
rect 20496 17756 20502 17808
rect 7285 17731 7343 17737
rect 5460 17700 6316 17728
rect 2774 17660 2780 17672
rect 1084 17632 2176 17660
rect 2332 17632 2780 17660
rect 1084 17620 1090 17632
rect 1486 17552 1492 17604
rect 1544 17592 1550 17604
rect 2148 17592 2176 17632
rect 2774 17620 2780 17632
rect 2832 17620 2838 17672
rect 4246 17660 4252 17672
rect 2884 17632 4252 17660
rect 2884 17592 2912 17632
rect 4246 17620 4252 17632
rect 4304 17620 4310 17672
rect 4798 17660 4804 17672
rect 4759 17632 4804 17660
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 5166 17620 5172 17672
rect 5224 17660 5230 17672
rect 5261 17663 5319 17669
rect 5261 17660 5273 17663
rect 5224 17632 5273 17660
rect 5224 17620 5230 17632
rect 5261 17629 5273 17632
rect 5307 17629 5319 17663
rect 6288 17660 6316 17700
rect 7285 17697 7297 17731
rect 7331 17728 7343 17731
rect 7650 17728 7656 17740
rect 7331 17700 7656 17728
rect 7331 17697 7343 17700
rect 7285 17691 7343 17697
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 8478 17728 8484 17740
rect 8439 17700 8484 17728
rect 8478 17688 8484 17700
rect 8536 17688 8542 17740
rect 8662 17688 8668 17740
rect 8720 17728 8726 17740
rect 10042 17728 10048 17740
rect 8720 17700 10048 17728
rect 8720 17688 8726 17700
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 11698 17728 11704 17740
rect 10152 17700 11704 17728
rect 8757 17663 8815 17669
rect 8757 17660 8769 17663
rect 6288 17632 8769 17660
rect 5261 17623 5319 17629
rect 8757 17629 8769 17632
rect 8803 17660 8815 17663
rect 10152 17660 10180 17700
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 11882 17688 11888 17740
rect 11940 17728 11946 17740
rect 12233 17731 12291 17737
rect 12233 17728 12245 17731
rect 11940 17700 12245 17728
rect 11940 17688 11946 17700
rect 12233 17697 12245 17700
rect 12279 17728 12291 17731
rect 13814 17728 13820 17740
rect 12279 17700 13820 17728
rect 12279 17697 12291 17700
rect 12233 17691 12291 17697
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 14550 17728 14556 17740
rect 14511 17700 14556 17728
rect 14550 17688 14556 17700
rect 14608 17688 14614 17740
rect 14645 17731 14703 17737
rect 14645 17697 14657 17731
rect 14691 17728 14703 17731
rect 15102 17728 15108 17740
rect 14691 17700 15108 17728
rect 14691 17697 14703 17700
rect 14645 17691 14703 17697
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 15562 17737 15568 17740
rect 15556 17728 15568 17737
rect 15523 17700 15568 17728
rect 15556 17691 15568 17700
rect 15562 17688 15568 17691
rect 15620 17688 15626 17740
rect 16758 17688 16764 17740
rect 16816 17728 16822 17740
rect 17678 17728 17684 17740
rect 16816 17700 17684 17728
rect 16816 17688 16822 17700
rect 17678 17688 17684 17700
rect 17736 17688 17742 17740
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 18417 17731 18475 17737
rect 18417 17728 18429 17731
rect 17819 17700 18429 17728
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 18417 17697 18429 17700
rect 18463 17728 18475 17731
rect 18463 17700 18644 17728
rect 18463 17697 18475 17700
rect 18417 17691 18475 17697
rect 8803 17632 10180 17660
rect 10321 17663 10379 17669
rect 8803 17629 8815 17632
rect 8757 17623 8815 17629
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 10594 17660 10600 17672
rect 10367 17632 10600 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 11790 17620 11796 17672
rect 11848 17660 11854 17672
rect 11977 17663 12035 17669
rect 11977 17660 11989 17663
rect 11848 17632 11989 17660
rect 11848 17620 11854 17632
rect 11977 17629 11989 17632
rect 12023 17629 12035 17663
rect 11977 17623 12035 17629
rect 12986 17620 12992 17672
rect 13044 17660 13050 17672
rect 14829 17663 14887 17669
rect 13044 17632 14780 17660
rect 13044 17620 13050 17632
rect 1544 17564 2084 17592
rect 2148 17564 2912 17592
rect 3053 17595 3111 17601
rect 1544 17552 1550 17564
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 2056 17524 2084 17564
rect 3053 17561 3065 17595
rect 3099 17592 3111 17595
rect 3326 17592 3332 17604
rect 3099 17564 3332 17592
rect 3099 17561 3111 17564
rect 3053 17555 3111 17561
rect 3326 17552 3332 17564
rect 3384 17552 3390 17604
rect 6270 17552 6276 17604
rect 6328 17592 6334 17604
rect 6328 17564 6776 17592
rect 6328 17552 6334 17564
rect 4062 17524 4068 17536
rect 2056 17496 4068 17524
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 4709 17527 4767 17533
rect 4709 17493 4721 17527
rect 4755 17524 4767 17527
rect 5994 17524 6000 17536
rect 4755 17496 6000 17524
rect 4755 17493 4767 17496
rect 4709 17487 4767 17493
rect 5994 17484 6000 17496
rect 6052 17524 6058 17536
rect 6638 17524 6644 17536
rect 6052 17496 6644 17524
rect 6052 17484 6058 17496
rect 6638 17484 6644 17496
rect 6696 17484 6702 17536
rect 6748 17524 6776 17564
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 9306 17592 9312 17604
rect 7340 17564 9312 17592
rect 7340 17552 7346 17564
rect 9306 17552 9312 17564
rect 9364 17552 9370 17604
rect 9677 17595 9735 17601
rect 9677 17561 9689 17595
rect 9723 17592 9735 17595
rect 10410 17592 10416 17604
rect 9723 17564 10416 17592
rect 9723 17561 9735 17564
rect 9677 17555 9735 17561
rect 10410 17552 10416 17564
rect 10468 17552 10474 17604
rect 13354 17592 13360 17604
rect 10520 17564 12020 17592
rect 13267 17564 13360 17592
rect 10520 17524 10548 17564
rect 6748 17496 10548 17524
rect 11149 17527 11207 17533
rect 11149 17493 11161 17527
rect 11195 17524 11207 17527
rect 11425 17527 11483 17533
rect 11425 17524 11437 17527
rect 11195 17496 11437 17524
rect 11195 17493 11207 17496
rect 11149 17487 11207 17493
rect 11425 17493 11437 17496
rect 11471 17524 11483 17527
rect 11698 17524 11704 17536
rect 11471 17496 11704 17524
rect 11471 17493 11483 17496
rect 11425 17487 11483 17493
rect 11698 17484 11704 17496
rect 11756 17484 11762 17536
rect 11882 17524 11888 17536
rect 11843 17496 11888 17524
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 11992 17524 12020 17564
rect 13354 17552 13360 17564
rect 13412 17592 13418 17604
rect 13998 17592 14004 17604
rect 13412 17564 14004 17592
rect 13412 17552 13418 17564
rect 13998 17552 14004 17564
rect 14056 17552 14062 17604
rect 14752 17592 14780 17632
rect 14829 17629 14841 17663
rect 14875 17660 14887 17663
rect 15010 17660 15016 17672
rect 14875 17632 15016 17660
rect 14875 17629 14887 17632
rect 14829 17623 14887 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15286 17660 15292 17672
rect 15247 17632 15292 17660
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 16945 17663 17003 17669
rect 16945 17660 16957 17663
rect 16540 17632 16957 17660
rect 16540 17620 16546 17632
rect 16945 17629 16957 17632
rect 16991 17660 17003 17663
rect 17310 17660 17316 17672
rect 16991 17632 17316 17660
rect 16991 17629 17003 17632
rect 16945 17623 17003 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 17957 17663 18015 17669
rect 17957 17660 17969 17663
rect 17920 17632 17969 17660
rect 17920 17620 17926 17632
rect 17957 17629 17969 17632
rect 18003 17629 18015 17663
rect 18616 17660 18644 17700
rect 19058 17688 19064 17740
rect 19116 17728 19122 17740
rect 20349 17731 20407 17737
rect 20349 17728 20361 17731
rect 19116 17700 20361 17728
rect 19116 17688 19122 17700
rect 20349 17697 20361 17700
rect 20395 17697 20407 17731
rect 20349 17691 20407 17697
rect 18877 17663 18935 17669
rect 18877 17660 18889 17663
rect 18616 17632 18889 17660
rect 17957 17623 18015 17629
rect 18877 17629 18889 17632
rect 18923 17629 18935 17663
rect 18877 17623 18935 17629
rect 15194 17592 15200 17604
rect 14752 17564 15200 17592
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 17402 17592 17408 17604
rect 17363 17564 17408 17592
rect 17402 17552 17408 17564
rect 17460 17552 17466 17604
rect 17586 17552 17592 17604
rect 17644 17592 17650 17604
rect 19981 17595 20039 17601
rect 19981 17592 19993 17595
rect 17644 17564 19993 17592
rect 17644 17552 17650 17564
rect 19981 17561 19993 17564
rect 20027 17561 20039 17595
rect 19981 17555 20039 17561
rect 16206 17524 16212 17536
rect 11992 17496 16212 17524
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16298 17484 16304 17536
rect 16356 17524 16362 17536
rect 16669 17527 16727 17533
rect 16669 17524 16681 17527
rect 16356 17496 16681 17524
rect 16356 17484 16362 17496
rect 16669 17493 16681 17496
rect 16715 17493 16727 17527
rect 16669 17487 16727 17493
rect 17494 17484 17500 17536
rect 17552 17524 17558 17536
rect 19245 17527 19303 17533
rect 19245 17524 19257 17527
rect 17552 17496 19257 17524
rect 17552 17484 17558 17496
rect 19245 17493 19257 17496
rect 19291 17493 19303 17527
rect 19245 17487 19303 17493
rect 19334 17484 19340 17536
rect 19392 17524 19398 17536
rect 19613 17527 19671 17533
rect 19613 17524 19625 17527
rect 19392 17496 19625 17524
rect 19392 17484 19398 17496
rect 19613 17493 19625 17496
rect 19659 17493 19671 17527
rect 19613 17487 19671 17493
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 2774 17320 2780 17332
rect 2056 17292 2780 17320
rect 1486 17116 1492 17128
rect 1447 17088 1492 17116
rect 1486 17076 1492 17088
rect 1544 17076 1550 17128
rect 2056 17125 2084 17292
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 2869 17323 2927 17329
rect 2869 17289 2881 17323
rect 2915 17320 2927 17323
rect 3234 17320 3240 17332
rect 2915 17292 3240 17320
rect 2915 17289 2927 17292
rect 2869 17283 2927 17289
rect 3234 17280 3240 17292
rect 3292 17280 3298 17332
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 10962 17320 10968 17332
rect 4120 17292 10824 17320
rect 10923 17292 10968 17320
rect 4120 17280 4126 17292
rect 4709 17255 4767 17261
rect 4709 17221 4721 17255
rect 4755 17252 4767 17255
rect 5902 17252 5908 17264
rect 4755 17224 5908 17252
rect 4755 17221 4767 17224
rect 4709 17215 4767 17221
rect 5902 17212 5908 17224
rect 5960 17212 5966 17264
rect 10796 17252 10824 17292
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 11882 17320 11888 17332
rect 11843 17292 11888 17320
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 19242 17320 19248 17332
rect 11992 17292 19248 17320
rect 11992 17252 12020 17292
rect 19242 17280 19248 17292
rect 19300 17280 19306 17332
rect 20438 17320 20444 17332
rect 20399 17292 20444 17320
rect 20438 17280 20444 17292
rect 20496 17280 20502 17332
rect 10796 17224 12020 17252
rect 14093 17255 14151 17261
rect 14093 17221 14105 17255
rect 14139 17252 14151 17255
rect 14274 17252 14280 17264
rect 14139 17224 14280 17252
rect 14139 17221 14151 17224
rect 14093 17215 14151 17221
rect 14274 17212 14280 17224
rect 14332 17212 14338 17264
rect 15654 17212 15660 17264
rect 15712 17252 15718 17264
rect 16025 17255 16083 17261
rect 16025 17252 16037 17255
rect 15712 17224 16037 17252
rect 15712 17212 15718 17224
rect 16025 17221 16037 17224
rect 16071 17221 16083 17255
rect 16482 17252 16488 17264
rect 16443 17224 16488 17252
rect 16025 17215 16083 17221
rect 16482 17212 16488 17224
rect 16540 17212 16546 17264
rect 16942 17252 16948 17264
rect 16903 17224 16948 17252
rect 16942 17212 16948 17224
rect 17000 17212 17006 17264
rect 17052 17224 17724 17252
rect 2314 17184 2320 17196
rect 2275 17156 2320 17184
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 2682 17144 2688 17196
rect 2740 17184 2746 17196
rect 2961 17187 3019 17193
rect 2961 17184 2973 17187
rect 2740 17156 2973 17184
rect 2740 17144 2746 17156
rect 2961 17153 2973 17156
rect 3007 17153 3019 17187
rect 2961 17147 3019 17153
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17184 5135 17187
rect 5813 17187 5871 17193
rect 5813 17184 5825 17187
rect 5123 17156 5825 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 5813 17153 5825 17156
rect 5859 17184 5871 17187
rect 6638 17184 6644 17196
rect 5859 17156 6644 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 8478 17144 8484 17196
rect 8536 17184 8542 17196
rect 9582 17184 9588 17196
rect 8536 17156 9588 17184
rect 8536 17144 8542 17156
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 11241 17187 11299 17193
rect 11241 17184 11253 17187
rect 10652 17156 11253 17184
rect 10652 17144 10658 17156
rect 11241 17153 11253 17156
rect 11287 17153 11299 17187
rect 11241 17147 11299 17153
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 12299 17156 12848 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 3234 17125 3240 17128
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17085 2099 17119
rect 3228 17116 3240 17125
rect 3195 17088 3240 17116
rect 2041 17079 2099 17085
rect 3228 17079 3240 17088
rect 3234 17076 3240 17079
rect 3292 17076 3298 17128
rect 4798 17076 4804 17128
rect 4856 17116 4862 17128
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 4856 17088 5549 17116
rect 4856 17076 4862 17088
rect 5537 17085 5549 17088
rect 5583 17116 5595 17119
rect 6181 17119 6239 17125
rect 6181 17116 6193 17119
rect 5583 17088 6193 17116
rect 5583 17085 5595 17088
rect 5537 17079 5595 17085
rect 6181 17085 6193 17088
rect 6227 17085 6239 17119
rect 6181 17079 6239 17085
rect 7098 17076 7104 17128
rect 7156 17116 7162 17128
rect 7558 17125 7564 17128
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 7156 17088 7297 17116
rect 7156 17076 7162 17088
rect 7285 17085 7297 17088
rect 7331 17085 7343 17119
rect 7552 17116 7564 17125
rect 7519 17088 7564 17116
rect 7285 17079 7343 17085
rect 7552 17079 7564 17088
rect 7558 17076 7564 17079
rect 7616 17076 7622 17128
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 7668 17088 9505 17116
rect 4246 17008 4252 17060
rect 4304 17048 4310 17060
rect 7668 17048 7696 17088
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 9852 17119 9910 17125
rect 9852 17116 9864 17119
rect 9493 17079 9551 17085
rect 9784 17088 9864 17116
rect 4304 17020 7696 17048
rect 9033 17051 9091 17057
rect 4304 17008 4310 17020
rect 9033 17017 9045 17051
rect 9079 17048 9091 17051
rect 9784 17048 9812 17088
rect 9852 17085 9864 17088
rect 9898 17116 9910 17119
rect 10612 17116 10640 17144
rect 9898 17088 10640 17116
rect 9898 17085 9910 17088
rect 9852 17079 9910 17085
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 11940 17088 12725 17116
rect 11940 17076 11946 17088
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 12820 17116 12848 17156
rect 16206 17144 16212 17196
rect 16264 17184 16270 17196
rect 17052 17184 17080 17224
rect 16264 17156 17080 17184
rect 16264 17144 16270 17156
rect 17310 17144 17316 17196
rect 17368 17184 17374 17196
rect 17405 17187 17463 17193
rect 17405 17184 17417 17187
rect 17368 17156 17417 17184
rect 17368 17144 17374 17156
rect 17405 17153 17417 17156
rect 17451 17153 17463 17187
rect 17586 17184 17592 17196
rect 17547 17156 17592 17184
rect 17405 17147 17463 17153
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 17696 17184 17724 17224
rect 17770 17212 17776 17264
rect 17828 17252 17834 17264
rect 17828 17224 18092 17252
rect 17828 17212 17834 17224
rect 18064 17193 18092 17224
rect 18049 17187 18107 17193
rect 17696 17156 18000 17184
rect 12980 17119 13038 17125
rect 12980 17116 12992 17119
rect 12820 17088 12992 17116
rect 12713 17079 12771 17085
rect 12980 17085 12992 17088
rect 13026 17116 13038 17119
rect 13354 17116 13360 17128
rect 13026 17088 13360 17116
rect 13026 17085 13038 17088
rect 12980 17079 13038 17085
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 14458 17076 14464 17128
rect 14516 17116 14522 17128
rect 14645 17119 14703 17125
rect 14645 17116 14657 17119
rect 14516 17088 14657 17116
rect 14516 17076 14522 17088
rect 14645 17085 14657 17088
rect 14691 17085 14703 17119
rect 17972 17116 18000 17156
rect 18049 17153 18061 17187
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 19058 17144 19064 17196
rect 19116 17184 19122 17196
rect 21177 17187 21235 17193
rect 21177 17184 21189 17187
rect 19116 17156 21189 17184
rect 19116 17144 19122 17156
rect 21177 17153 21189 17156
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 20073 17119 20131 17125
rect 20073 17116 20085 17119
rect 17972 17088 20085 17116
rect 14645 17079 14703 17085
rect 20073 17085 20085 17088
rect 20119 17085 20131 17119
rect 20073 17079 20131 17085
rect 13814 17048 13820 17060
rect 9079 17020 9812 17048
rect 9876 17020 13820 17048
rect 9079 17017 9091 17020
rect 9033 17011 9091 17017
rect 1673 16983 1731 16989
rect 1673 16949 1685 16983
rect 1719 16980 1731 16983
rect 2958 16980 2964 16992
rect 1719 16952 2964 16980
rect 1719 16949 1731 16952
rect 1673 16943 1731 16949
rect 2958 16940 2964 16952
rect 3016 16940 3022 16992
rect 4338 16980 4344 16992
rect 4299 16952 4344 16980
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 5169 16983 5227 16989
rect 5169 16949 5181 16983
rect 5215 16980 5227 16983
rect 5258 16980 5264 16992
rect 5215 16952 5264 16980
rect 5215 16949 5227 16952
rect 5169 16943 5227 16949
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 5629 16983 5687 16989
rect 5629 16949 5641 16983
rect 5675 16980 5687 16983
rect 6270 16980 6276 16992
rect 5675 16952 6276 16980
rect 5675 16949 5687 16952
rect 5629 16943 5687 16949
rect 6270 16940 6276 16952
rect 6328 16940 6334 16992
rect 6362 16940 6368 16992
rect 6420 16980 6426 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6420 16952 6561 16980
rect 6420 16940 6426 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 6549 16943 6607 16949
rect 7193 16983 7251 16989
rect 7193 16949 7205 16983
rect 7239 16980 7251 16983
rect 7374 16980 7380 16992
rect 7239 16952 7380 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7374 16940 7380 16952
rect 7432 16980 7438 16992
rect 8202 16980 8208 16992
rect 7432 16952 8208 16980
rect 7432 16940 7438 16952
rect 8202 16940 8208 16952
rect 8260 16980 8266 16992
rect 8665 16983 8723 16989
rect 8665 16980 8677 16983
rect 8260 16952 8677 16980
rect 8260 16940 8266 16952
rect 8665 16949 8677 16952
rect 8711 16949 8723 16983
rect 8665 16943 8723 16949
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16980 9183 16983
rect 9398 16980 9404 16992
rect 9171 16952 9404 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 9493 16983 9551 16989
rect 9493 16949 9505 16983
rect 9539 16980 9551 16983
rect 9876 16980 9904 17020
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 14890 17051 14948 17057
rect 14890 17048 14902 17051
rect 14568 17020 14902 17048
rect 14568 16992 14596 17020
rect 14890 17017 14902 17020
rect 14936 17017 14948 17051
rect 14890 17011 14948 17017
rect 15010 17008 15016 17060
rect 15068 17048 15074 17060
rect 16206 17048 16212 17060
rect 15068 17020 16212 17048
rect 15068 17008 15074 17020
rect 16206 17008 16212 17020
rect 16264 17008 16270 17060
rect 16316 17020 17540 17048
rect 9539 16952 9904 16980
rect 9539 16949 9551 16952
rect 9493 16943 9551 16949
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 13906 16980 13912 16992
rect 10560 16952 13912 16980
rect 10560 16940 10566 16952
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 14550 16980 14556 16992
rect 14511 16952 14556 16980
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 16316 16980 16344 17020
rect 15160 16952 16344 16980
rect 15160 16940 15166 16952
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 16761 16983 16819 16989
rect 16761 16980 16773 16983
rect 16724 16952 16773 16980
rect 16724 16940 16730 16952
rect 16761 16949 16773 16952
rect 16807 16980 16819 16983
rect 17313 16983 17371 16989
rect 17313 16980 17325 16983
rect 16807 16952 17325 16980
rect 16807 16949 16819 16952
rect 16761 16943 16819 16949
rect 17313 16949 17325 16952
rect 17359 16949 17371 16983
rect 17512 16980 17540 17020
rect 17862 17008 17868 17060
rect 17920 17048 17926 17060
rect 18294 17051 18352 17057
rect 18294 17048 18306 17051
rect 17920 17020 18306 17048
rect 17920 17008 17926 17020
rect 18294 17017 18306 17020
rect 18340 17048 18352 17051
rect 19610 17048 19616 17060
rect 18340 17020 19616 17048
rect 18340 17017 18352 17020
rect 18294 17011 18352 17017
rect 19610 17008 19616 17020
rect 19668 17048 19674 17060
rect 19705 17051 19763 17057
rect 19705 17048 19717 17051
rect 19668 17020 19717 17048
rect 19668 17008 19674 17020
rect 19705 17017 19717 17020
rect 19751 17017 19763 17051
rect 19705 17011 19763 17017
rect 19334 16980 19340 16992
rect 17512 16952 19340 16980
rect 17313 16943 17371 16949
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 19484 16952 19529 16980
rect 19484 16940 19490 16952
rect 19978 16940 19984 16992
rect 20036 16980 20042 16992
rect 20809 16983 20867 16989
rect 20809 16980 20821 16983
rect 20036 16952 20821 16980
rect 20036 16940 20042 16952
rect 20809 16949 20821 16952
rect 20855 16949 20867 16983
rect 20809 16943 20867 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1762 16776 1768 16788
rect 1723 16748 1768 16776
rect 1762 16736 1768 16748
rect 1820 16736 1826 16788
rect 2314 16736 2320 16788
rect 2372 16736 2378 16788
rect 4525 16779 4583 16785
rect 4525 16745 4537 16779
rect 4571 16776 4583 16779
rect 4706 16776 4712 16788
rect 4571 16748 4712 16776
rect 4571 16745 4583 16748
rect 4525 16739 4583 16745
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 6638 16776 6644 16788
rect 4816 16748 6644 16776
rect 2332 16708 2360 16736
rect 1596 16680 2360 16708
rect 1596 16649 1624 16680
rect 3050 16668 3056 16720
rect 3108 16708 3114 16720
rect 4816 16708 4844 16748
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 7558 16736 7564 16788
rect 7616 16776 7622 16788
rect 7837 16779 7895 16785
rect 7837 16776 7849 16779
rect 7616 16748 7849 16776
rect 7616 16736 7622 16748
rect 7837 16745 7849 16748
rect 7883 16745 7895 16779
rect 7837 16739 7895 16745
rect 7929 16779 7987 16785
rect 7929 16745 7941 16779
rect 7975 16776 7987 16779
rect 8294 16776 8300 16788
rect 7975 16748 8300 16776
rect 7975 16745 7987 16748
rect 7929 16739 7987 16745
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 9398 16776 9404 16788
rect 9359 16748 9404 16776
rect 9398 16736 9404 16748
rect 9456 16776 9462 16788
rect 10045 16779 10103 16785
rect 10045 16776 10057 16779
rect 9456 16748 10057 16776
rect 9456 16736 9462 16748
rect 10045 16745 10057 16748
rect 10091 16745 10103 16779
rect 10045 16739 10103 16745
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 10410 16776 10416 16788
rect 10183 16748 10416 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 10962 16736 10968 16788
rect 11020 16776 11026 16788
rect 11057 16779 11115 16785
rect 11057 16776 11069 16779
rect 11020 16748 11069 16776
rect 11020 16736 11026 16748
rect 11057 16745 11069 16748
rect 11103 16745 11115 16779
rect 11057 16739 11115 16745
rect 11425 16779 11483 16785
rect 11425 16745 11437 16779
rect 11471 16776 11483 16779
rect 11606 16776 11612 16788
rect 11471 16748 11612 16776
rect 11471 16745 11483 16748
rect 11425 16739 11483 16745
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 11885 16779 11943 16785
rect 11885 16745 11897 16779
rect 11931 16776 11943 16779
rect 12342 16776 12348 16788
rect 11931 16748 12348 16776
rect 11931 16745 11943 16748
rect 11885 16739 11943 16745
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 12897 16779 12955 16785
rect 12897 16745 12909 16779
rect 12943 16776 12955 16779
rect 13354 16776 13360 16788
rect 12943 16748 13360 16776
rect 12943 16745 12955 16748
rect 12897 16739 12955 16745
rect 13354 16736 13360 16748
rect 13412 16776 13418 16788
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 13412 16748 13461 16776
rect 13412 16736 13418 16748
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 13814 16776 13820 16788
rect 13775 16748 13820 16776
rect 13449 16739 13507 16745
rect 13814 16736 13820 16748
rect 13872 16736 13878 16788
rect 13906 16736 13912 16788
rect 13964 16776 13970 16788
rect 13964 16748 14009 16776
rect 13964 16736 13970 16748
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 15286 16776 15292 16788
rect 14516 16748 15292 16776
rect 14516 16736 14522 16748
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15654 16776 15660 16788
rect 15615 16748 15660 16776
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 16301 16779 16359 16785
rect 16301 16745 16313 16779
rect 16347 16776 16359 16779
rect 17586 16776 17592 16788
rect 16347 16748 17592 16776
rect 16347 16745 16359 16748
rect 16301 16739 16359 16745
rect 17586 16736 17592 16748
rect 17644 16776 17650 16788
rect 17773 16779 17831 16785
rect 17773 16776 17785 16779
rect 17644 16748 17785 16776
rect 17644 16736 17650 16748
rect 17773 16745 17785 16748
rect 17819 16745 17831 16779
rect 17773 16739 17831 16745
rect 19429 16779 19487 16785
rect 19429 16745 19441 16779
rect 19475 16776 19487 16779
rect 19610 16776 19616 16788
rect 19475 16748 19616 16776
rect 19475 16745 19487 16748
rect 19429 16739 19487 16745
rect 6914 16708 6920 16720
rect 3108 16680 4844 16708
rect 6380 16680 6920 16708
rect 3108 16668 3114 16680
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16609 1639 16643
rect 1581 16603 1639 16609
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16640 2191 16643
rect 2314 16640 2320 16652
rect 2179 16612 2320 16640
rect 2179 16609 2191 16612
rect 2133 16603 2191 16609
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 3234 16640 3240 16652
rect 3195 16612 3240 16640
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 3329 16643 3387 16649
rect 3329 16609 3341 16643
rect 3375 16609 3387 16643
rect 3329 16603 3387 16609
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 5169 16643 5227 16649
rect 5169 16640 5181 16643
rect 4479 16612 5181 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 5169 16609 5181 16612
rect 5215 16640 5227 16643
rect 5718 16640 5724 16652
rect 5215 16612 5724 16640
rect 5215 16609 5227 16612
rect 5169 16603 5227 16609
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16572 2467 16575
rect 2866 16572 2872 16584
rect 2455 16544 2872 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 3344 16504 3372 16603
rect 5718 16600 5724 16612
rect 5776 16600 5782 16652
rect 6380 16649 6408 16680
rect 6914 16668 6920 16680
rect 6972 16708 6978 16720
rect 9950 16708 9956 16720
rect 6972 16680 9956 16708
rect 6972 16668 6978 16680
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 17494 16708 17500 16720
rect 10060 16680 17500 16708
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 6365 16643 6423 16649
rect 5951 16612 6316 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 3513 16575 3571 16581
rect 3513 16541 3525 16575
rect 3559 16572 3571 16575
rect 4062 16572 4068 16584
rect 3559 16544 4068 16572
rect 3559 16541 3571 16544
rect 3513 16535 3571 16541
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4396 16544 4629 16572
rect 4396 16532 4402 16544
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 5258 16572 5264 16584
rect 5219 16544 5264 16572
rect 4617 16535 4675 16541
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 6288 16572 6316 16612
rect 6365 16609 6377 16643
rect 6411 16609 6423 16643
rect 6638 16640 6644 16652
rect 6599 16612 6644 16640
rect 6365 16603 6423 16609
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 7650 16640 7656 16652
rect 6748 16612 7656 16640
rect 6748 16572 6776 16612
rect 7650 16600 7656 16612
rect 7708 16640 7714 16652
rect 8665 16643 8723 16649
rect 8665 16640 8677 16643
rect 7708 16612 7788 16640
rect 7708 16600 7714 16612
rect 6288 16544 6776 16572
rect 7377 16575 7435 16581
rect 7377 16541 7389 16575
rect 7423 16572 7435 16575
rect 7466 16572 7472 16584
rect 7423 16544 7472 16572
rect 7423 16541 7435 16544
rect 7377 16535 7435 16541
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 7760 16572 7788 16612
rect 8036 16612 8677 16640
rect 8036 16572 8064 16612
rect 8665 16609 8677 16612
rect 8711 16609 8723 16643
rect 8665 16603 8723 16609
rect 8754 16600 8760 16652
rect 8812 16640 8818 16652
rect 10060 16640 10088 16680
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 17788 16708 17816 16739
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 19794 16736 19800 16788
rect 19852 16776 19858 16788
rect 20441 16779 20499 16785
rect 20441 16776 20453 16779
rect 19852 16748 20453 16776
rect 19852 16736 19858 16748
rect 20441 16745 20453 16748
rect 20487 16745 20499 16779
rect 20441 16739 20499 16745
rect 20806 16736 20812 16788
rect 20864 16776 20870 16788
rect 21085 16779 21143 16785
rect 21085 16776 21097 16779
rect 20864 16748 21097 16776
rect 20864 16736 20870 16748
rect 21085 16745 21097 16748
rect 21131 16745 21143 16779
rect 21085 16739 21143 16745
rect 17788 16680 17908 16708
rect 8812 16612 10088 16640
rect 11793 16643 11851 16649
rect 8812 16600 8818 16612
rect 11793 16609 11805 16643
rect 11839 16640 11851 16643
rect 11839 16612 12296 16640
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 7760 16544 8064 16572
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16572 8171 16575
rect 8202 16572 8208 16584
rect 8159 16544 8208 16572
rect 8159 16541 8171 16544
rect 8113 16535 8171 16541
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 10962 16572 10968 16584
rect 10367 16544 10968 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11977 16575 12035 16581
rect 11977 16541 11989 16575
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 3344 16476 11652 16504
rect 2406 16396 2412 16448
rect 2464 16436 2470 16448
rect 4080 16445 4108 16476
rect 2869 16439 2927 16445
rect 2869 16436 2881 16439
rect 2464 16408 2881 16436
rect 2464 16396 2470 16408
rect 2869 16405 2881 16408
rect 2915 16405 2927 16439
rect 2869 16399 2927 16405
rect 4065 16439 4123 16445
rect 4065 16405 4077 16439
rect 4111 16405 4123 16439
rect 4065 16399 4123 16405
rect 4798 16396 4804 16448
rect 4856 16436 4862 16448
rect 5166 16436 5172 16448
rect 4856 16408 5172 16436
rect 4856 16396 4862 16408
rect 5166 16396 5172 16408
rect 5224 16436 5230 16448
rect 5721 16439 5779 16445
rect 5721 16436 5733 16439
rect 5224 16408 5733 16436
rect 5224 16396 5230 16408
rect 5721 16405 5733 16408
rect 5767 16405 5779 16439
rect 6178 16436 6184 16448
rect 6139 16408 6184 16436
rect 5721 16399 5779 16405
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 7469 16439 7527 16445
rect 7469 16436 7481 16439
rect 7340 16408 7481 16436
rect 7340 16396 7346 16408
rect 7469 16405 7481 16408
rect 7515 16405 7527 16439
rect 8478 16436 8484 16448
rect 8439 16408 8484 16436
rect 7469 16399 7527 16405
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 9122 16436 9128 16448
rect 9083 16408 9128 16436
rect 9122 16396 9128 16408
rect 9180 16396 9186 16448
rect 9306 16396 9312 16448
rect 9364 16436 9370 16448
rect 9677 16439 9735 16445
rect 9677 16436 9689 16439
rect 9364 16408 9689 16436
rect 9364 16396 9370 16408
rect 9677 16405 9689 16408
rect 9723 16405 9735 16439
rect 9677 16399 9735 16405
rect 9950 16396 9956 16448
rect 10008 16436 10014 16448
rect 10689 16439 10747 16445
rect 10689 16436 10701 16439
rect 10008 16408 10701 16436
rect 10008 16396 10014 16408
rect 10689 16405 10701 16408
rect 10735 16405 10747 16439
rect 11624 16436 11652 16476
rect 11698 16464 11704 16516
rect 11756 16504 11762 16516
rect 11992 16504 12020 16535
rect 11756 16476 12020 16504
rect 11756 16464 11762 16476
rect 12158 16436 12164 16448
rect 11624 16408 12164 16436
rect 10689 16399 10747 16405
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 12268 16436 12296 16612
rect 12342 16600 12348 16652
rect 12400 16640 12406 16652
rect 12805 16643 12863 16649
rect 12400 16612 12480 16640
rect 12400 16600 12406 16612
rect 12452 16513 12480 16612
rect 12805 16609 12817 16643
rect 12851 16640 12863 16643
rect 13538 16640 13544 16652
rect 12851 16612 13544 16640
rect 12851 16609 12863 16612
rect 12805 16603 12863 16609
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 13630 16600 13636 16652
rect 13688 16640 13694 16652
rect 13906 16640 13912 16652
rect 13688 16612 13912 16640
rect 13688 16600 13694 16612
rect 13906 16600 13912 16612
rect 13964 16640 13970 16652
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 13964 16612 14473 16640
rect 13964 16600 13970 16612
rect 14461 16609 14473 16612
rect 14507 16609 14519 16643
rect 14461 16603 14519 16609
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 16660 16643 16718 16649
rect 16080 16612 16252 16640
rect 16080 16600 16086 16612
rect 12710 16532 12716 16584
rect 12768 16572 12774 16584
rect 13081 16575 13139 16581
rect 13081 16572 13093 16575
rect 12768 16544 13093 16572
rect 12768 16532 12774 16544
rect 13081 16541 13093 16544
rect 13127 16572 13139 16575
rect 13998 16572 14004 16584
rect 13127 16544 14004 16572
rect 13127 16541 13139 16544
rect 13081 16535 13139 16541
rect 13998 16532 14004 16544
rect 14056 16532 14062 16584
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 14274 16572 14280 16584
rect 14139 16544 14280 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 12437 16507 12495 16513
rect 12437 16473 12449 16507
rect 12483 16473 12495 16507
rect 16224 16504 16252 16612
rect 16660 16609 16672 16643
rect 16706 16640 16718 16643
rect 17126 16640 17132 16652
rect 16706 16612 17132 16640
rect 16706 16609 16718 16612
rect 16660 16603 16718 16609
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 17678 16600 17684 16652
rect 17736 16640 17742 16652
rect 17880 16640 17908 16680
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 19705 16711 19763 16717
rect 19705 16708 19717 16711
rect 18104 16680 19717 16708
rect 18104 16668 18110 16680
rect 19705 16677 19717 16680
rect 19751 16677 19763 16711
rect 19705 16671 19763 16677
rect 18316 16643 18374 16649
rect 18316 16640 18328 16643
rect 17736 16612 17816 16640
rect 17880 16612 18328 16640
rect 17736 16600 17742 16612
rect 16298 16532 16304 16584
rect 16356 16572 16362 16584
rect 16400 16575 16458 16581
rect 16400 16572 16412 16575
rect 16356 16544 16412 16572
rect 16356 16532 16362 16544
rect 16400 16541 16412 16544
rect 16446 16541 16458 16575
rect 17788 16572 17816 16612
rect 18316 16609 18328 16612
rect 18362 16640 18374 16643
rect 19334 16640 19340 16652
rect 18362 16612 19340 16640
rect 18362 16609 18374 16612
rect 18316 16603 18374 16609
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 20073 16643 20131 16649
rect 20073 16640 20085 16643
rect 19435 16612 20085 16640
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17788 16544 18061 16572
rect 16400 16535 16458 16541
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 16224 16476 16436 16504
rect 12437 16467 12495 16473
rect 12618 16436 12624 16448
rect 12268 16408 12624 16436
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 14921 16439 14979 16445
rect 14921 16405 14933 16439
rect 14967 16436 14979 16439
rect 15194 16436 15200 16448
rect 14967 16408 15200 16436
rect 14967 16405 14979 16408
rect 14921 16399 14979 16405
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 16408 16436 16436 16476
rect 19435 16436 19463 16612
rect 20073 16609 20085 16612
rect 20119 16609 20131 16643
rect 20073 16603 20131 16609
rect 16408 16408 19463 16436
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2130 16192 2136 16244
rect 2188 16192 2194 16244
rect 4062 16232 4068 16244
rect 4023 16204 4068 16232
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 4525 16235 4583 16241
rect 4525 16201 4537 16235
rect 4571 16232 4583 16235
rect 4706 16232 4712 16244
rect 4571 16204 4712 16232
rect 4571 16201 4583 16204
rect 4525 16195 4583 16201
rect 4706 16192 4712 16204
rect 4764 16192 4770 16244
rect 5902 16192 5908 16244
rect 5960 16232 5966 16244
rect 6273 16235 6331 16241
rect 6273 16232 6285 16235
rect 5960 16204 6285 16232
rect 5960 16192 5966 16204
rect 6273 16201 6285 16204
rect 6319 16201 6331 16235
rect 6273 16195 6331 16201
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 8352 16204 8769 16232
rect 8352 16192 8358 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 8757 16195 8815 16201
rect 10321 16235 10379 16241
rect 10321 16201 10333 16235
rect 10367 16232 10379 16235
rect 10594 16232 10600 16244
rect 10367 16204 10600 16232
rect 10367 16201 10379 16204
rect 10321 16195 10379 16201
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 10704 16204 11652 16232
rect 2148 16164 2176 16192
rect 2314 16164 2320 16176
rect 1412 16136 2320 16164
rect 1412 16037 1440 16136
rect 2314 16124 2320 16136
rect 2372 16124 2378 16176
rect 1486 16056 1492 16108
rect 1544 16096 1550 16108
rect 2133 16099 2191 16105
rect 2133 16096 2145 16099
rect 1544 16068 2145 16096
rect 1544 16056 1550 16068
rect 2133 16065 2145 16068
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 6641 16099 6699 16105
rect 6641 16065 6653 16099
rect 6687 16096 6699 16099
rect 6687 16068 7236 16096
rect 6687 16065 6699 16068
rect 6641 16059 6699 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 15997 2007 16031
rect 2682 16028 2688 16040
rect 2643 16000 2688 16028
rect 1949 15991 2007 15997
rect 1964 15960 1992 15991
rect 2682 15988 2688 16000
rect 2740 15988 2746 16040
rect 2958 16037 2964 16040
rect 2952 16028 2964 16037
rect 2871 16000 2964 16028
rect 2952 15991 2964 16000
rect 3016 16028 3022 16040
rect 4246 16028 4252 16040
rect 3016 16000 4252 16028
rect 2958 15988 2964 15991
rect 3016 15988 3022 16000
rect 4246 15988 4252 16000
rect 4304 15988 4310 16040
rect 4798 15988 4804 16040
rect 4856 16028 4862 16040
rect 4893 16031 4951 16037
rect 4893 16028 4905 16031
rect 4856 16000 4905 16028
rect 4856 15988 4862 16000
rect 4893 15997 4905 16000
rect 4939 15997 4951 16031
rect 7098 16028 7104 16040
rect 7011 16000 7104 16028
rect 4893 15991 4951 15997
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 7208 16028 7236 16068
rect 7374 16037 7380 16040
rect 7368 16028 7380 16037
rect 7208 16000 7380 16028
rect 7368 15991 7380 16000
rect 7374 15988 7380 15991
rect 7432 15988 7438 16040
rect 8478 15988 8484 16040
rect 8536 16028 8542 16040
rect 8941 16031 8999 16037
rect 8941 16028 8953 16031
rect 8536 16000 8953 16028
rect 8536 15988 8542 16000
rect 8941 15997 8953 16000
rect 8987 15997 8999 16031
rect 8941 15991 8999 15997
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 10704 16037 10732 16204
rect 11624 16164 11652 16204
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 12069 16235 12127 16241
rect 12069 16232 12081 16235
rect 11756 16204 12081 16232
rect 11756 16192 11762 16204
rect 12069 16201 12081 16204
rect 12115 16201 12127 16235
rect 12069 16195 12127 16201
rect 12158 16192 12164 16244
rect 12216 16232 12222 16244
rect 17862 16232 17868 16244
rect 12216 16204 16528 16232
rect 17823 16204 17868 16232
rect 12216 16192 12222 16204
rect 11882 16164 11888 16176
rect 11624 16136 11888 16164
rect 11882 16124 11888 16136
rect 11940 16164 11946 16176
rect 14921 16167 14979 16173
rect 14921 16164 14933 16167
rect 11940 16136 13308 16164
rect 11940 16124 11946 16136
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 12986 16096 12992 16108
rect 12667 16068 12992 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 10689 16031 10747 16037
rect 10689 16028 10701 16031
rect 10652 16000 10701 16028
rect 10652 15988 10658 16000
rect 10689 15997 10701 16000
rect 10735 15997 10747 16031
rect 10689 15991 10747 15997
rect 10956 16031 11014 16037
rect 10956 15997 10968 16031
rect 11002 16028 11014 16031
rect 12710 16028 12716 16040
rect 11002 16000 12716 16028
rect 11002 15997 11014 16000
rect 10956 15991 11014 15997
rect 12710 15988 12716 16000
rect 12768 15988 12774 16040
rect 13280 16037 13308 16136
rect 14292 16136 14933 16164
rect 13265 16031 13323 16037
rect 13265 15997 13277 16031
rect 13311 16028 13323 16031
rect 14292 16028 14320 16136
rect 14921 16133 14933 16136
rect 14967 16133 14979 16167
rect 14921 16127 14979 16133
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 15933 16167 15991 16173
rect 15933 16164 15945 16167
rect 15344 16136 15945 16164
rect 15344 16124 15350 16136
rect 15933 16133 15945 16136
rect 15979 16164 15991 16167
rect 16390 16164 16396 16176
rect 15979 16136 16396 16164
rect 15979 16133 15991 16136
rect 15933 16127 15991 16133
rect 16390 16124 16396 16136
rect 16448 16124 16454 16176
rect 16500 16164 16528 16204
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 18012 16204 18061 16232
rect 18012 16192 18018 16204
rect 18049 16201 18061 16204
rect 18095 16201 18107 16235
rect 18049 16195 18107 16201
rect 19334 16192 19340 16244
rect 19392 16232 19398 16244
rect 19429 16235 19487 16241
rect 19429 16232 19441 16235
rect 19392 16204 19441 16232
rect 19392 16192 19398 16204
rect 19429 16201 19441 16204
rect 19475 16201 19487 16235
rect 19429 16195 19487 16201
rect 20533 16167 20591 16173
rect 20533 16164 20545 16167
rect 16500 16136 20545 16164
rect 20533 16133 20545 16136
rect 20579 16133 20591 16167
rect 20533 16127 20591 16133
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16096 18751 16099
rect 19242 16096 19248 16108
rect 18739 16068 19248 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 13311 16000 14320 16028
rect 15105 16031 15163 16037
rect 13311 15997 13323 16000
rect 13265 15991 13323 15997
rect 15105 15997 15117 16031
rect 15151 16028 15163 16031
rect 16114 16028 16120 16040
rect 15151 16000 16120 16028
rect 15151 15997 15163 16000
rect 15105 15991 15163 15997
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 17920 16000 18521 16028
rect 17920 15988 17926 16000
rect 18509 15997 18521 16000
rect 18555 16028 18567 16031
rect 20901 16031 20959 16037
rect 20901 16028 20913 16031
rect 18555 16000 20913 16028
rect 18555 15997 18567 16000
rect 18509 15991 18567 15997
rect 20901 15997 20913 16000
rect 20947 15997 20959 16031
rect 20901 15991 20959 15997
rect 2130 15960 2136 15972
rect 1964 15932 2136 15960
rect 2130 15920 2136 15932
rect 2188 15920 2194 15972
rect 5160 15963 5218 15969
rect 5160 15929 5172 15963
rect 5206 15960 5218 15963
rect 6178 15960 6184 15972
rect 5206 15932 6184 15960
rect 5206 15929 5218 15932
rect 5160 15923 5218 15929
rect 6178 15920 6184 15932
rect 6236 15920 6242 15972
rect 7116 15960 7144 15988
rect 8496 15960 8524 15988
rect 7116 15932 8524 15960
rect 9122 15920 9128 15972
rect 9180 15969 9186 15972
rect 9180 15963 9244 15969
rect 9180 15929 9198 15963
rect 9232 15929 9244 15963
rect 9180 15923 9244 15929
rect 9180 15920 9186 15923
rect 9582 15920 9588 15972
rect 9640 15960 9646 15972
rect 13532 15963 13590 15969
rect 9640 15932 13492 15960
rect 9640 15920 9646 15932
rect 2222 15852 2228 15904
rect 2280 15892 2286 15904
rect 3970 15892 3976 15904
rect 2280 15864 3976 15892
rect 2280 15852 2286 15864
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 8481 15895 8539 15901
rect 8481 15892 8493 15895
rect 7524 15864 8493 15892
rect 7524 15852 7530 15864
rect 8481 15861 8493 15864
rect 8527 15861 8539 15895
rect 12802 15892 12808 15904
rect 12763 15864 12808 15892
rect 8481 15855 8539 15861
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 13464 15892 13492 15932
rect 13532 15929 13544 15963
rect 13578 15960 13590 15963
rect 14274 15960 14280 15972
rect 13578 15932 14280 15960
rect 13578 15929 13590 15932
rect 13532 15923 13590 15929
rect 14274 15920 14280 15932
rect 14332 15920 14338 15972
rect 18417 15963 18475 15969
rect 14660 15932 17264 15960
rect 13906 15892 13912 15904
rect 13464 15864 13912 15892
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 13998 15852 14004 15904
rect 14056 15892 14062 15904
rect 14660 15901 14688 15932
rect 14645 15895 14703 15901
rect 14645 15892 14657 15895
rect 14056 15864 14657 15892
rect 14056 15852 14062 15864
rect 14645 15861 14657 15864
rect 14691 15861 14703 15895
rect 14645 15855 14703 15861
rect 15102 15852 15108 15904
rect 15160 15892 15166 15904
rect 15381 15895 15439 15901
rect 15381 15892 15393 15895
rect 15160 15864 15393 15892
rect 15160 15852 15166 15864
rect 15381 15861 15393 15864
rect 15427 15861 15439 15895
rect 15381 15855 15439 15861
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 15749 15895 15807 15901
rect 15749 15892 15761 15895
rect 15620 15864 15761 15892
rect 15620 15852 15626 15864
rect 15749 15861 15761 15864
rect 15795 15861 15807 15895
rect 15749 15855 15807 15861
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 16393 15895 16451 15901
rect 16393 15892 16405 15895
rect 16264 15864 16405 15892
rect 16264 15852 16270 15864
rect 16393 15861 16405 15864
rect 16439 15861 16451 15895
rect 16393 15855 16451 15861
rect 16853 15895 16911 15901
rect 16853 15861 16865 15895
rect 16899 15892 16911 15895
rect 17126 15892 17132 15904
rect 16899 15864 17132 15892
rect 16899 15861 16911 15864
rect 16853 15855 16911 15861
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 17236 15892 17264 15932
rect 18417 15929 18429 15963
rect 18463 15960 18475 15963
rect 18874 15960 18880 15972
rect 18463 15932 18880 15960
rect 18463 15929 18475 15932
rect 18417 15923 18475 15929
rect 18874 15920 18880 15932
rect 18932 15960 18938 15972
rect 19061 15963 19119 15969
rect 19061 15960 19073 15963
rect 18932 15932 19073 15960
rect 18932 15920 18938 15932
rect 19061 15929 19073 15932
rect 19107 15929 19119 15963
rect 19061 15923 19119 15929
rect 19242 15920 19248 15972
rect 19300 15960 19306 15972
rect 19797 15963 19855 15969
rect 19797 15960 19809 15963
rect 19300 15932 19809 15960
rect 19300 15920 19306 15932
rect 19797 15929 19809 15932
rect 19843 15929 19855 15963
rect 19797 15923 19855 15929
rect 19610 15892 19616 15904
rect 17236 15864 19616 15892
rect 19610 15852 19616 15864
rect 19668 15852 19674 15904
rect 20162 15892 20168 15904
rect 20123 15864 20168 15892
rect 20162 15852 20168 15864
rect 20220 15852 20226 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 2041 15691 2099 15697
rect 2041 15657 2053 15691
rect 2087 15688 2099 15691
rect 2409 15691 2467 15697
rect 2409 15688 2421 15691
rect 2087 15660 2421 15688
rect 2087 15657 2099 15660
rect 2041 15651 2099 15657
rect 2409 15657 2421 15660
rect 2455 15688 2467 15691
rect 2958 15688 2964 15700
rect 2455 15660 2964 15688
rect 2455 15657 2467 15660
rect 2409 15651 2467 15657
rect 2958 15648 2964 15660
rect 3016 15648 3022 15700
rect 3234 15688 3240 15700
rect 3195 15660 3240 15688
rect 3234 15648 3240 15660
rect 3292 15688 3298 15700
rect 3697 15691 3755 15697
rect 3697 15688 3709 15691
rect 3292 15660 3709 15688
rect 3292 15648 3298 15660
rect 3697 15657 3709 15660
rect 3743 15657 3755 15691
rect 3697 15651 3755 15657
rect 4706 15648 4712 15700
rect 4764 15688 4770 15700
rect 4985 15691 5043 15697
rect 4985 15688 4997 15691
rect 4764 15660 4997 15688
rect 4764 15648 4770 15660
rect 4985 15657 4997 15660
rect 5031 15688 5043 15691
rect 5258 15688 5264 15700
rect 5031 15660 5264 15688
rect 5031 15657 5043 15660
rect 4985 15651 5043 15657
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 6089 15691 6147 15697
rect 6089 15657 6101 15691
rect 6135 15688 6147 15691
rect 6546 15688 6552 15700
rect 6135 15660 6552 15688
rect 6135 15657 6147 15660
rect 6089 15651 6147 15657
rect 6546 15648 6552 15660
rect 6604 15648 6610 15700
rect 6914 15688 6920 15700
rect 6875 15660 6920 15688
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 8570 15648 8576 15700
rect 8628 15688 8634 15700
rect 9033 15691 9091 15697
rect 9033 15688 9045 15691
rect 8628 15660 9045 15688
rect 8628 15648 8634 15660
rect 9033 15657 9045 15660
rect 9079 15688 9091 15691
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 9079 15660 9689 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 9677 15651 9735 15657
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 10226 15688 10232 15700
rect 10183 15660 10232 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 12342 15688 12348 15700
rect 12124 15660 12348 15688
rect 12124 15648 12130 15660
rect 12342 15648 12348 15660
rect 12400 15648 12406 15700
rect 12897 15691 12955 15697
rect 12897 15657 12909 15691
rect 12943 15688 12955 15691
rect 13170 15688 13176 15700
rect 12943 15660 13176 15688
rect 12943 15657 12955 15660
rect 12897 15651 12955 15657
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 13906 15688 13912 15700
rect 13867 15660 13912 15688
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 15841 15691 15899 15697
rect 15841 15657 15853 15691
rect 15887 15657 15899 15691
rect 16206 15688 16212 15700
rect 16167 15660 16212 15688
rect 15841 15651 15899 15657
rect 3970 15580 3976 15632
rect 4028 15620 4034 15632
rect 14001 15623 14059 15629
rect 14001 15620 14013 15623
rect 4028 15592 14013 15620
rect 4028 15580 4034 15592
rect 14001 15589 14013 15592
rect 14047 15620 14059 15623
rect 14918 15620 14924 15632
rect 14047 15592 14924 15620
rect 14047 15589 14059 15592
rect 14001 15583 14059 15589
rect 14918 15580 14924 15592
rect 14976 15580 14982 15632
rect 15856 15620 15884 15651
rect 16206 15648 16212 15660
rect 16264 15688 16270 15700
rect 16853 15691 16911 15697
rect 16853 15688 16865 15691
rect 16264 15660 16865 15688
rect 16264 15648 16270 15660
rect 16853 15657 16865 15660
rect 16899 15657 16911 15691
rect 17862 15688 17868 15700
rect 17823 15660 17868 15688
rect 16853 15651 16911 15657
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 17954 15648 17960 15700
rect 18012 15648 18018 15700
rect 18874 15688 18880 15700
rect 18835 15660 18880 15688
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 19426 15688 19432 15700
rect 19387 15660 19432 15688
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19610 15648 19616 15700
rect 19668 15688 19674 15700
rect 20073 15691 20131 15697
rect 20073 15688 20085 15691
rect 19668 15660 20085 15688
rect 19668 15648 19674 15660
rect 20073 15657 20085 15660
rect 20119 15657 20131 15691
rect 20073 15651 20131 15657
rect 16758 15620 16764 15632
rect 15856 15592 16764 15620
rect 16758 15580 16764 15592
rect 16816 15580 16822 15632
rect 17972 15620 18000 15648
rect 20441 15623 20499 15629
rect 20441 15620 20453 15623
rect 17972 15592 20453 15620
rect 20441 15589 20453 15592
rect 20487 15589 20499 15623
rect 20441 15583 20499 15589
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 3142 15552 3148 15564
rect 2823 15524 3148 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 3142 15512 3148 15524
rect 3200 15552 3206 15564
rect 4062 15552 4068 15564
rect 3200 15524 4068 15552
rect 3200 15512 3206 15524
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 4571 15524 5304 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 5276 15493 5304 15524
rect 5810 15512 5816 15564
rect 5868 15552 5874 15564
rect 5997 15555 6055 15561
rect 5997 15552 6009 15555
rect 5868 15524 6009 15552
rect 5868 15512 5874 15524
rect 5997 15521 6009 15524
rect 6043 15552 6055 15555
rect 6641 15555 6699 15561
rect 6641 15552 6653 15555
rect 6043 15524 6653 15552
rect 6043 15521 6055 15524
rect 5997 15515 6055 15521
rect 6641 15521 6653 15524
rect 6687 15521 6699 15555
rect 6641 15515 6699 15521
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 7926 15552 7932 15564
rect 7331 15524 7932 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 5077 15487 5135 15493
rect 5077 15453 5089 15487
rect 5123 15453 5135 15487
rect 5077 15447 5135 15453
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15484 5319 15487
rect 6086 15484 6092 15496
rect 5307 15456 6092 15484
rect 5307 15453 5319 15456
rect 5261 15447 5319 15453
rect 5092 15416 5120 15447
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15484 6331 15487
rect 6362 15484 6368 15496
rect 6319 15456 6368 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 6362 15444 6368 15456
rect 6420 15444 6426 15496
rect 6656 15416 6684 15515
rect 7926 15512 7932 15524
rect 7984 15512 7990 15564
rect 8938 15552 8944 15564
rect 8036 15524 8800 15552
rect 8899 15524 8944 15552
rect 7374 15484 7380 15496
rect 7335 15456 7380 15484
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 7524 15456 7569 15484
rect 7524 15444 7530 15456
rect 8036 15416 8064 15524
rect 8772 15484 8800 15524
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9048 15524 10057 15552
rect 9048 15484 9076 15524
rect 10045 15521 10057 15524
rect 10091 15552 10103 15555
rect 10502 15552 10508 15564
rect 10091 15524 10508 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 11048 15555 11106 15561
rect 11048 15521 11060 15555
rect 11094 15552 11106 15555
rect 11606 15552 11612 15564
rect 11094 15524 11612 15552
rect 11094 15521 11106 15524
rect 11048 15515 11106 15521
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 13906 15512 13912 15564
rect 13964 15552 13970 15564
rect 14734 15552 14740 15564
rect 13964 15524 14740 15552
rect 13964 15512 13970 15524
rect 14734 15512 14740 15524
rect 14792 15552 14798 15564
rect 15102 15552 15108 15564
rect 14792 15524 15108 15552
rect 14792 15512 14798 15524
rect 15102 15512 15108 15524
rect 15160 15552 15166 15564
rect 15473 15555 15531 15561
rect 15473 15552 15485 15555
rect 15160 15524 15485 15552
rect 15160 15512 15166 15524
rect 15473 15521 15485 15524
rect 15519 15552 15531 15555
rect 15519 15524 17264 15552
rect 15519 15521 15531 15524
rect 15473 15515 15531 15521
rect 8772 15456 9076 15484
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9180 15456 9225 15484
rect 9180 15444 9186 15456
rect 10134 15444 10140 15496
rect 10192 15484 10198 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 10192 15456 10241 15484
rect 10192 15444 10198 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10594 15444 10600 15496
rect 10652 15484 10658 15496
rect 10781 15487 10839 15493
rect 10781 15484 10793 15487
rect 10652 15456 10793 15484
rect 10652 15444 10658 15456
rect 10781 15453 10793 15456
rect 10827 15453 10839 15487
rect 12986 15484 12992 15496
rect 12947 15456 12992 15484
rect 10781 15447 10839 15453
rect 12986 15444 12992 15456
rect 13044 15444 13050 15496
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15484 13231 15487
rect 14185 15487 14243 15493
rect 14185 15484 14197 15487
rect 13219 15456 14197 15484
rect 13219 15453 13231 15456
rect 13173 15447 13231 15453
rect 14185 15453 14197 15456
rect 14231 15484 14243 15487
rect 14274 15484 14280 15496
rect 14231 15456 14280 15484
rect 14231 15453 14243 15456
rect 14185 15447 14243 15453
rect 14274 15444 14280 15456
rect 14332 15484 14338 15496
rect 16298 15484 16304 15496
rect 14332 15456 15783 15484
rect 16259 15456 16304 15484
rect 14332 15444 14338 15456
rect 8570 15416 8576 15428
rect 5092 15388 5672 15416
rect 6656 15388 8064 15416
rect 8531 15388 8576 15416
rect 5644 15360 5672 15388
rect 8570 15376 8576 15388
rect 8628 15376 8634 15428
rect 13814 15376 13820 15428
rect 13872 15416 13878 15428
rect 14553 15419 14611 15425
rect 14553 15416 14565 15419
rect 13872 15388 14565 15416
rect 13872 15376 13878 15388
rect 14553 15385 14565 15388
rect 14599 15385 14611 15419
rect 15755 15416 15783 15456
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 16485 15487 16543 15493
rect 16485 15453 16497 15487
rect 16531 15484 16543 15487
rect 17126 15484 17132 15496
rect 16531 15456 17132 15484
rect 16531 15453 16543 15456
rect 16485 15447 16543 15453
rect 17126 15444 17132 15456
rect 17184 15444 17190 15496
rect 17236 15484 17264 15524
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18233 15555 18291 15561
rect 18233 15552 18245 15555
rect 18012 15524 18245 15552
rect 18012 15512 18018 15524
rect 18233 15521 18245 15524
rect 18279 15521 18291 15555
rect 18233 15515 18291 15521
rect 18690 15512 18696 15564
rect 18748 15552 18754 15564
rect 21085 15555 21143 15561
rect 21085 15552 21097 15555
rect 18748 15524 21097 15552
rect 18748 15512 18754 15524
rect 21085 15521 21097 15524
rect 21131 15521 21143 15555
rect 21085 15515 21143 15521
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 17236 15456 18337 15484
rect 18325 15453 18337 15456
rect 18371 15484 18383 15487
rect 18414 15484 18420 15496
rect 18371 15456 18420 15484
rect 18371 15453 18383 15456
rect 18325 15447 18383 15453
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15484 18567 15487
rect 19426 15484 19432 15496
rect 18555 15456 19432 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19705 15419 19763 15425
rect 19705 15416 19717 15419
rect 15755 15388 19717 15416
rect 14553 15379 14611 15385
rect 19705 15385 19717 15388
rect 19751 15416 19763 15419
rect 20162 15416 20168 15428
rect 19751 15388 20168 15416
rect 19751 15385 19763 15388
rect 19705 15379 19763 15385
rect 20162 15376 20168 15388
rect 20220 15376 20226 15428
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 2130 15308 2136 15360
rect 2188 15348 2194 15360
rect 4617 15351 4675 15357
rect 4617 15348 4629 15351
rect 2188 15320 4629 15348
rect 2188 15308 2194 15320
rect 4617 15317 4629 15320
rect 4663 15317 4675 15351
rect 5626 15348 5632 15360
rect 5587 15320 5632 15348
rect 4617 15311 4675 15317
rect 5626 15308 5632 15320
rect 5684 15308 5690 15360
rect 5718 15308 5724 15360
rect 5776 15348 5782 15360
rect 6638 15348 6644 15360
rect 5776 15320 6644 15348
rect 5776 15308 5782 15320
rect 6638 15308 6644 15320
rect 6696 15348 6702 15360
rect 7558 15348 7564 15360
rect 6696 15320 7564 15348
rect 6696 15308 6702 15320
rect 7558 15308 7564 15320
rect 7616 15348 7622 15360
rect 8389 15351 8447 15357
rect 8389 15348 8401 15351
rect 7616 15320 8401 15348
rect 7616 15308 7622 15320
rect 8389 15317 8401 15320
rect 8435 15317 8447 15351
rect 8389 15311 8447 15317
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 12161 15351 12219 15357
rect 12161 15348 12173 15351
rect 11112 15320 12173 15348
rect 11112 15308 11118 15320
rect 12161 15317 12173 15320
rect 12207 15348 12219 15351
rect 12342 15348 12348 15360
rect 12207 15320 12348 15348
rect 12207 15317 12219 15320
rect 12161 15311 12219 15317
rect 12342 15308 12348 15320
rect 12400 15308 12406 15360
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 13078 15348 13084 15360
rect 12575 15320 13084 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 13078 15308 13084 15320
rect 13136 15308 13142 15360
rect 13538 15348 13544 15360
rect 13499 15320 13544 15348
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 15746 15308 15752 15360
rect 15804 15348 15810 15360
rect 16390 15348 16396 15360
rect 15804 15320 16396 15348
rect 15804 15308 15810 15320
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 16758 15308 16764 15360
rect 16816 15348 16822 15360
rect 17405 15351 17463 15357
rect 17405 15348 17417 15351
rect 16816 15320 17417 15348
rect 16816 15308 16822 15320
rect 17405 15317 17417 15320
rect 17451 15348 17463 15351
rect 17494 15348 17500 15360
rect 17451 15320 17500 15348
rect 17451 15317 17463 15320
rect 17405 15311 17463 15317
rect 17494 15308 17500 15320
rect 17552 15308 17558 15360
rect 17770 15348 17776 15360
rect 17731 15320 17776 15348
rect 17770 15308 17776 15320
rect 17828 15308 17834 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 4706 15144 4712 15156
rect 4667 15116 4712 15144
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 6178 15144 6184 15156
rect 6139 15116 6184 15144
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 6546 15144 6552 15156
rect 6507 15116 6552 15144
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 7926 15144 7932 15156
rect 7887 15116 7932 15144
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 8573 15147 8631 15153
rect 8573 15113 8585 15147
rect 8619 15144 8631 15147
rect 8938 15144 8944 15156
rect 8619 15116 8944 15144
rect 8619 15113 8631 15116
rect 8573 15107 8631 15113
rect 8938 15104 8944 15116
rect 8996 15104 9002 15156
rect 10226 15104 10232 15156
rect 10284 15144 10290 15156
rect 10321 15147 10379 15153
rect 10321 15144 10333 15147
rect 10284 15116 10333 15144
rect 10284 15104 10290 15116
rect 10321 15113 10333 15116
rect 10367 15113 10379 15147
rect 10321 15107 10379 15113
rect 10502 15104 10508 15156
rect 10560 15144 10566 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 10560 15116 10701 15144
rect 10560 15104 10566 15116
rect 10689 15113 10701 15116
rect 10735 15113 10747 15147
rect 11146 15144 11152 15156
rect 11107 15116 11152 15144
rect 10689 15107 10747 15113
rect 11146 15104 11152 15116
rect 11204 15104 11210 15156
rect 14001 15147 14059 15153
rect 12636 15116 13952 15144
rect 1302 15036 1308 15088
rect 1360 15076 1366 15088
rect 1581 15079 1639 15085
rect 1581 15076 1593 15079
rect 1360 15048 1593 15076
rect 1360 15036 1366 15048
rect 1581 15045 1593 15048
rect 1627 15045 1639 15079
rect 1581 15039 1639 15045
rect 7101 15079 7159 15085
rect 7101 15045 7113 15079
rect 7147 15076 7159 15079
rect 7650 15076 7656 15088
rect 7147 15048 7656 15076
rect 7147 15045 7159 15048
rect 7101 15039 7159 15045
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 15008 2283 15011
rect 2314 15008 2320 15020
rect 2271 14980 2320 15008
rect 2271 14977 2283 14980
rect 2225 14971 2283 14977
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 11164 15008 11192 15104
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11164 14980 11805 15008
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 15008 12035 15011
rect 12342 15008 12348 15020
rect 12023 14980 12348 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1486 14940 1492 14952
rect 1443 14912 1492 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1486 14900 1492 14912
rect 1544 14900 1550 14952
rect 1946 14940 1952 14952
rect 1907 14912 1952 14940
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 3142 14949 3148 14952
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14940 2927 14943
rect 2915 14912 3011 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 2590 14832 2596 14884
rect 2648 14872 2654 14884
rect 2685 14875 2743 14881
rect 2685 14872 2697 14875
rect 2648 14844 2697 14872
rect 2648 14832 2654 14844
rect 2685 14841 2697 14844
rect 2731 14841 2743 14875
rect 2685 14835 2743 14841
rect 2983 14804 3011 14912
rect 3136 14903 3148 14949
rect 3200 14940 3206 14952
rect 4798 14940 4804 14952
rect 3200 14912 3236 14940
rect 4759 14912 4804 14940
rect 3142 14900 3148 14903
rect 3200 14900 3206 14912
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 4890 14900 4896 14952
rect 4948 14940 4954 14952
rect 5068 14943 5126 14949
rect 5068 14940 5080 14943
rect 4948 14912 5080 14940
rect 4948 14900 4954 14912
rect 5068 14909 5080 14912
rect 5114 14940 5126 14943
rect 6362 14940 6368 14952
rect 5114 14912 6368 14940
rect 5114 14909 5126 14912
rect 5068 14903 5126 14909
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 7282 14940 7288 14952
rect 7243 14912 7288 14940
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 8478 14900 8484 14952
rect 8536 14940 8542 14952
rect 8665 14943 8723 14949
rect 8665 14940 8677 14943
rect 8536 14912 8677 14940
rect 8536 14900 8542 14912
rect 8665 14909 8677 14912
rect 8711 14909 8723 14943
rect 12636 14940 12664 15116
rect 12894 15036 12900 15088
rect 12952 15076 12958 15088
rect 13262 15076 13268 15088
rect 12952 15048 13268 15076
rect 12952 15036 12958 15048
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 13924 15076 13952 15116
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 16114 15144 16120 15156
rect 14047 15116 16120 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 16390 15104 16396 15156
rect 16448 15144 16454 15156
rect 17126 15144 17132 15156
rect 16448 15116 16712 15144
rect 17087 15116 17132 15144
rect 16448 15104 16454 15116
rect 15654 15076 15660 15088
rect 13924 15048 15660 15076
rect 15654 15036 15660 15048
rect 15712 15036 15718 15088
rect 16684 15076 16712 15116
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 17221 15147 17279 15153
rect 17221 15113 17233 15147
rect 17267 15144 17279 15147
rect 19334 15144 19340 15156
rect 17267 15116 19340 15144
rect 17267 15113 17279 15116
rect 17221 15107 17279 15113
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 20162 15104 20168 15156
rect 20220 15144 20226 15156
rect 20257 15147 20315 15153
rect 20257 15144 20269 15147
rect 20220 15116 20269 15144
rect 20220 15104 20226 15116
rect 20257 15113 20269 15116
rect 20303 15113 20315 15147
rect 20257 15107 20315 15113
rect 16684 15048 17724 15076
rect 17696 15020 17724 15048
rect 19242 15036 19248 15088
rect 19300 15076 19306 15088
rect 19613 15079 19671 15085
rect 19613 15076 19625 15079
rect 19300 15048 19625 15076
rect 19300 15036 19306 15048
rect 19613 15045 19625 15048
rect 19659 15045 19671 15079
rect 19613 15039 19671 15045
rect 12710 14968 12716 15020
rect 12768 15008 12774 15020
rect 13173 15011 13231 15017
rect 13173 15008 13185 15011
rect 12768 14980 13185 15008
rect 12768 14968 12774 14980
rect 13173 14977 13185 14980
rect 13219 14977 13231 15011
rect 13998 15008 14004 15020
rect 13173 14971 13231 14977
rect 13280 14980 14004 15008
rect 8665 14903 8723 14909
rect 9324 14912 12664 14940
rect 9324 14884 9352 14912
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 12989 14943 13047 14949
rect 12989 14940 13001 14943
rect 12860 14912 13001 14940
rect 12860 14900 12866 14912
rect 12989 14909 13001 14912
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 13280 14940 13308 14980
rect 13998 14968 14004 14980
rect 14056 14968 14062 15020
rect 14826 15008 14832 15020
rect 14787 14980 14832 15008
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 15008 15071 15011
rect 15194 15008 15200 15020
rect 15059 14980 15200 15008
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 15746 15008 15752 15020
rect 15707 14980 15752 15008
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 16850 14968 16856 15020
rect 16908 15008 16914 15020
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 16908 14980 17417 15008
rect 16908 14968 16914 14980
rect 17405 14977 17417 14980
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 17678 14968 17684 15020
rect 17736 15008 17742 15020
rect 19889 15011 19947 15017
rect 19889 15008 19901 15011
rect 17736 14980 18276 15008
rect 17736 14968 17742 14980
rect 13136 14912 13308 14940
rect 13136 14900 13142 14912
rect 13906 14900 13912 14952
rect 13964 14940 13970 14952
rect 14185 14943 14243 14949
rect 14185 14940 14197 14943
rect 13964 14912 14197 14940
rect 13964 14900 13970 14912
rect 14185 14909 14197 14912
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 14734 14940 14740 14952
rect 14332 14912 14596 14940
rect 14695 14912 14740 14940
rect 14332 14900 14338 14912
rect 8846 14832 8852 14884
rect 8904 14881 8910 14884
rect 8904 14875 8968 14881
rect 8904 14841 8922 14875
rect 8956 14841 8968 14875
rect 8904 14835 8968 14841
rect 8904 14832 8910 14835
rect 9306 14832 9312 14884
rect 9364 14832 9370 14884
rect 9398 14832 9404 14884
rect 9456 14872 9462 14884
rect 10134 14872 10140 14884
rect 9456 14844 10140 14872
rect 9456 14832 9462 14844
rect 10134 14832 10140 14844
rect 10192 14832 10198 14884
rect 11348 14844 11919 14872
rect 3050 14804 3056 14816
rect 2983 14776 3056 14804
rect 3050 14764 3056 14776
rect 3108 14764 3114 14816
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 4249 14807 4307 14813
rect 4249 14804 4261 14807
rect 4120 14776 4261 14804
rect 4120 14764 4126 14776
rect 4249 14773 4261 14776
rect 4295 14773 4307 14807
rect 7558 14804 7564 14816
rect 7519 14776 7564 14804
rect 4249 14767 4307 14773
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 9122 14764 9128 14816
rect 9180 14804 9186 14816
rect 11348 14813 11376 14844
rect 10045 14807 10103 14813
rect 10045 14804 10057 14807
rect 9180 14776 10057 14804
rect 9180 14764 9186 14776
rect 10045 14773 10057 14776
rect 10091 14773 10103 14807
rect 10045 14767 10103 14773
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14773 11391 14807
rect 11698 14804 11704 14816
rect 11659 14776 11704 14804
rect 11333 14767 11391 14773
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 11891 14804 11919 14844
rect 12526 14804 12532 14816
rect 11891 14776 12532 14804
rect 12526 14764 12532 14776
rect 12584 14764 12590 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 12986 14804 12992 14816
rect 12676 14776 12992 14804
rect 12676 14764 12682 14776
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 13078 14764 13084 14816
rect 13136 14804 13142 14816
rect 13633 14807 13691 14813
rect 13633 14804 13645 14807
rect 13136 14776 13645 14804
rect 13136 14764 13142 14776
rect 13633 14773 13645 14776
rect 13679 14773 13691 14807
rect 14366 14804 14372 14816
rect 14327 14776 14372 14804
rect 13633 14767 13691 14773
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 14568 14804 14596 14912
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 14844 14940 14872 14968
rect 15378 14940 15384 14952
rect 14844 14912 15384 14940
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 18248 14949 18276 14980
rect 19444 14980 19901 15008
rect 19444 14952 19472 14980
rect 19889 14977 19901 14980
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 18233 14943 18291 14949
rect 16356 14912 18092 14940
rect 16356 14900 16362 14912
rect 16016 14875 16074 14881
rect 16016 14841 16028 14875
rect 16062 14872 16074 14875
rect 16758 14872 16764 14884
rect 16062 14844 16764 14872
rect 16062 14841 16074 14844
rect 16016 14835 16074 14841
rect 16758 14832 16764 14844
rect 16816 14832 16822 14884
rect 17310 14832 17316 14884
rect 17368 14872 17374 14884
rect 17773 14875 17831 14881
rect 17773 14872 17785 14875
rect 17368 14844 17785 14872
rect 17368 14832 17374 14844
rect 17773 14841 17785 14844
rect 17819 14872 17831 14875
rect 17954 14872 17960 14884
rect 17819 14844 17960 14872
rect 17819 14841 17831 14844
rect 17773 14835 17831 14841
rect 17954 14832 17960 14844
rect 18012 14832 18018 14884
rect 18064 14872 18092 14912
rect 18233 14909 18245 14943
rect 18279 14940 18291 14943
rect 18322 14940 18328 14952
rect 18279 14912 18328 14940
rect 18279 14909 18291 14912
rect 18233 14903 18291 14909
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 18500 14943 18558 14949
rect 18500 14909 18512 14943
rect 18546 14940 18558 14943
rect 19426 14940 19432 14952
rect 18546 14912 19432 14940
rect 18546 14909 18558 14912
rect 18500 14903 18558 14909
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 19610 14900 19616 14952
rect 19668 14940 19674 14952
rect 20993 14943 21051 14949
rect 20993 14940 21005 14943
rect 19668 14912 21005 14940
rect 19668 14900 19674 14912
rect 20993 14909 21005 14912
rect 21039 14909 21051 14943
rect 20993 14903 21051 14909
rect 20625 14875 20683 14881
rect 20625 14872 20637 14875
rect 18064 14844 20637 14872
rect 20625 14841 20637 14844
rect 20671 14841 20683 14875
rect 20625 14835 20683 14841
rect 17221 14807 17279 14813
rect 17221 14804 17233 14807
rect 14568 14776 17233 14804
rect 17221 14773 17233 14776
rect 17267 14773 17279 14807
rect 17221 14767 17279 14773
rect 17494 14764 17500 14816
rect 17552 14804 17558 14816
rect 19426 14804 19432 14816
rect 17552 14776 19432 14804
rect 17552 14764 17558 14776
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 2038 14600 2044 14612
rect 1627 14572 2044 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 2038 14560 2044 14572
rect 2096 14560 2102 14612
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4525 14603 4583 14609
rect 4525 14600 4537 14603
rect 4212 14572 4537 14600
rect 4212 14560 4218 14572
rect 4525 14569 4537 14572
rect 4571 14600 4583 14603
rect 5077 14603 5135 14609
rect 5077 14600 5089 14603
rect 4571 14572 5089 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 5077 14569 5089 14572
rect 5123 14569 5135 14603
rect 5077 14563 5135 14569
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 7742 14600 7748 14612
rect 6595 14572 7748 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 8996 14572 9045 14600
rect 8996 14560 9002 14572
rect 9033 14569 9045 14572
rect 9079 14569 9091 14603
rect 10134 14600 10140 14612
rect 10095 14572 10140 14600
rect 9033 14563 9091 14569
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 12802 14600 12808 14612
rect 10643 14572 12808 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 13633 14603 13691 14609
rect 13633 14600 13645 14603
rect 13219 14572 13645 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 13633 14569 13645 14572
rect 13679 14569 13691 14603
rect 13633 14563 13691 14569
rect 14016 14572 14320 14600
rect 5718 14532 5724 14544
rect 2240 14504 5724 14532
rect 2240 14476 2268 14504
rect 5718 14492 5724 14504
rect 5776 14492 5782 14544
rect 7374 14492 7380 14544
rect 7432 14532 7438 14544
rect 8389 14535 8447 14541
rect 7432 14504 7604 14532
rect 7432 14492 7438 14504
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2222 14464 2228 14476
rect 1995 14436 2228 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 2222 14424 2228 14436
rect 2280 14424 2286 14476
rect 3326 14464 3332 14476
rect 3287 14436 3332 14464
rect 3326 14424 3332 14436
rect 3384 14424 3390 14476
rect 3421 14467 3479 14473
rect 3421 14433 3433 14467
rect 3467 14464 3479 14467
rect 3602 14464 3608 14476
rect 3467 14436 3608 14464
rect 3467 14433 3479 14436
rect 3421 14427 3479 14433
rect 3602 14424 3608 14436
rect 3660 14424 3666 14476
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 4706 14464 4712 14476
rect 4479 14436 4712 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 6914 14473 6920 14476
rect 6908 14464 6920 14473
rect 6875 14436 6920 14464
rect 6908 14427 6920 14436
rect 6972 14464 6978 14476
rect 7466 14464 7472 14476
rect 6972 14436 7472 14464
rect 6914 14424 6920 14427
rect 6972 14424 6978 14436
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 7576 14464 7604 14504
rect 8389 14501 8401 14535
rect 8435 14532 8447 14535
rect 9122 14532 9128 14544
rect 8435 14504 9128 14532
rect 8435 14501 8447 14504
rect 8389 14495 8447 14501
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 14016 14532 14044 14572
rect 14185 14535 14243 14541
rect 14185 14532 14197 14535
rect 9232 14504 14044 14532
rect 14108 14504 14197 14532
rect 9232 14464 9260 14504
rect 14108 14476 14136 14504
rect 14185 14501 14197 14504
rect 14231 14501 14243 14535
rect 14292 14532 14320 14572
rect 15654 14560 15660 14612
rect 15712 14600 15718 14612
rect 15933 14603 15991 14609
rect 15933 14600 15945 14603
rect 15712 14572 15945 14600
rect 15712 14560 15718 14572
rect 15933 14569 15945 14572
rect 15979 14569 15991 14603
rect 15933 14563 15991 14569
rect 16577 14603 16635 14609
rect 16577 14569 16589 14603
rect 16623 14600 16635 14603
rect 18506 14600 18512 14612
rect 16623 14572 18512 14600
rect 16623 14569 16635 14572
rect 16577 14563 16635 14569
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 18966 14560 18972 14612
rect 19024 14600 19030 14612
rect 21085 14603 21143 14609
rect 21085 14600 21097 14603
rect 19024 14572 21097 14600
rect 19024 14560 19030 14572
rect 21085 14569 21097 14572
rect 21131 14569 21143 14603
rect 21085 14563 21143 14569
rect 18325 14535 18383 14541
rect 14292 14504 17080 14532
rect 14185 14495 14243 14501
rect 7576 14436 9260 14464
rect 10318 14424 10324 14476
rect 10376 14464 10382 14476
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 10376 14436 11253 14464
rect 10376 14424 10382 14436
rect 11241 14433 11253 14436
rect 11287 14464 11299 14467
rect 11793 14467 11851 14473
rect 11793 14464 11805 14467
rect 11287 14436 11805 14464
rect 11287 14433 11299 14436
rect 11241 14427 11299 14433
rect 11793 14433 11805 14436
rect 11839 14433 11851 14467
rect 12342 14464 12348 14476
rect 11793 14427 11851 14433
rect 12084 14436 12348 14464
rect 1486 14356 1492 14408
rect 1544 14396 1550 14408
rect 2133 14399 2191 14405
rect 2133 14396 2145 14399
rect 1544 14368 2145 14396
rect 1544 14356 1550 14368
rect 2133 14365 2145 14368
rect 2179 14396 2191 14399
rect 2314 14396 2320 14408
rect 2179 14368 2320 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 3513 14399 3571 14405
rect 3513 14365 3525 14399
rect 3559 14396 3571 14399
rect 4154 14396 4160 14408
rect 3559 14368 4160 14396
rect 3559 14365 3571 14368
rect 3513 14359 3571 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 2590 14288 2596 14340
rect 2648 14328 2654 14340
rect 2961 14331 3019 14337
rect 2961 14328 2973 14331
rect 2648 14300 2973 14328
rect 2648 14288 2654 14300
rect 2961 14297 2973 14300
rect 3007 14297 3019 14331
rect 3970 14328 3976 14340
rect 2961 14291 3019 14297
rect 3528 14300 3976 14328
rect 2866 14260 2872 14272
rect 2827 14232 2872 14260
rect 2866 14220 2872 14232
rect 2924 14260 2930 14272
rect 3528 14260 3556 14300
rect 3970 14288 3976 14300
rect 4028 14328 4034 14340
rect 4632 14328 4660 14359
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 6638 14396 6644 14408
rect 4856 14368 6644 14396
rect 4856 14356 4862 14368
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11698 14396 11704 14408
rect 11011 14368 11704 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 11882 14396 11888 14408
rect 11843 14368 11888 14396
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 12084 14405 12112 14436
rect 12342 14424 12348 14436
rect 12400 14464 12406 14476
rect 13722 14464 13728 14476
rect 12400 14436 13728 14464
rect 12400 14424 12406 14436
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 14090 14464 14096 14476
rect 13872 14436 14096 14464
rect 13872 14424 13878 14436
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 14550 14464 14556 14476
rect 14200 14436 14556 14464
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14365 12127 14399
rect 12069 14359 12127 14365
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 13262 14396 13268 14408
rect 12492 14368 12537 14396
rect 13223 14368 13268 14396
rect 12492 14356 12498 14368
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14396 13507 14399
rect 14200 14396 14228 14436
rect 14550 14424 14556 14436
rect 14608 14464 14614 14476
rect 14608 14436 15332 14464
rect 14608 14424 14614 14436
rect 13495 14368 14228 14396
rect 14277 14399 14335 14405
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 14277 14365 14289 14399
rect 14323 14396 14335 14399
rect 14461 14399 14519 14405
rect 14323 14368 14403 14396
rect 14323 14365 14335 14368
rect 14277 14359 14335 14365
rect 4028 14300 4660 14328
rect 5813 14331 5871 14337
rect 4028 14288 4034 14300
rect 5813 14297 5825 14331
rect 5859 14328 5871 14331
rect 6270 14328 6276 14340
rect 5859 14300 6276 14328
rect 5859 14297 5871 14300
rect 5813 14291 5871 14297
rect 6270 14288 6276 14300
rect 6328 14288 6334 14340
rect 11425 14331 11483 14337
rect 11425 14297 11437 14331
rect 11471 14328 11483 14331
rect 12618 14328 12624 14340
rect 11471 14300 12624 14328
rect 11471 14297 11483 14300
rect 11425 14291 11483 14297
rect 12618 14288 12624 14300
rect 12676 14288 12682 14340
rect 12805 14331 12863 14337
rect 12805 14297 12817 14331
rect 12851 14328 12863 14331
rect 12894 14328 12900 14340
rect 12851 14300 12900 14328
rect 12851 14297 12863 14300
rect 12805 14291 12863 14297
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13633 14331 13691 14337
rect 13633 14297 13645 14331
rect 13679 14328 13691 14331
rect 14375 14328 14403 14368
rect 14461 14365 14473 14399
rect 14507 14396 14519 14399
rect 15194 14396 15200 14408
rect 14507 14368 15200 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 15304 14396 15332 14436
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 15930 14464 15936 14476
rect 15436 14436 15936 14464
rect 15436 14424 15442 14436
rect 15930 14424 15936 14436
rect 15988 14464 15994 14476
rect 16025 14467 16083 14473
rect 16025 14464 16037 14467
rect 15988 14436 16037 14464
rect 15988 14424 15994 14436
rect 16025 14433 16037 14436
rect 16071 14433 16083 14467
rect 16942 14464 16948 14476
rect 16903 14436 16948 14464
rect 16025 14427 16083 14433
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17052 14464 17080 14504
rect 18325 14501 18337 14535
rect 18371 14532 18383 14535
rect 18414 14532 18420 14544
rect 18371 14504 18420 14532
rect 18371 14501 18383 14504
rect 18325 14495 18383 14501
rect 18414 14492 18420 14504
rect 18472 14492 18478 14544
rect 18684 14535 18742 14541
rect 18684 14501 18696 14535
rect 18730 14532 18742 14535
rect 18782 14532 18788 14544
rect 18730 14504 18788 14532
rect 18730 14501 18742 14504
rect 18684 14495 18742 14501
rect 18782 14492 18788 14504
rect 18840 14532 18846 14544
rect 19242 14532 19248 14544
rect 18840 14504 19248 14532
rect 18840 14492 18846 14504
rect 19242 14492 19248 14504
rect 19300 14492 19306 14544
rect 19334 14492 19340 14544
rect 19392 14532 19398 14544
rect 20441 14535 20499 14541
rect 20441 14532 20453 14535
rect 19392 14504 20453 14532
rect 19392 14492 19398 14504
rect 20441 14501 20453 14504
rect 20487 14501 20499 14535
rect 20441 14495 20499 14501
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 17052 14436 20085 14464
rect 20073 14433 20085 14436
rect 20119 14433 20131 14467
rect 20073 14427 20131 14433
rect 16209 14399 16267 14405
rect 15304 14368 15424 14396
rect 15396 14340 15424 14368
rect 16209 14365 16221 14399
rect 16255 14396 16267 14399
rect 16758 14396 16764 14408
rect 16255 14368 16764 14396
rect 16255 14365 16267 14368
rect 16209 14359 16267 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 17037 14399 17095 14405
rect 17037 14396 17049 14399
rect 16908 14368 17049 14396
rect 16908 14356 16914 14368
rect 17037 14365 17049 14368
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 17221 14399 17279 14405
rect 17221 14365 17233 14399
rect 17267 14365 17279 14399
rect 17221 14359 17279 14365
rect 17589 14399 17647 14405
rect 17589 14365 17601 14399
rect 17635 14396 17647 14399
rect 17954 14396 17960 14408
rect 17635 14368 17960 14396
rect 17635 14365 17647 14368
rect 17589 14359 17647 14365
rect 13679 14300 14320 14328
rect 14375 14300 14504 14328
rect 13679 14297 13691 14300
rect 13633 14291 13691 14297
rect 14292 14272 14320 14300
rect 14476 14272 14504 14300
rect 15378 14288 15384 14340
rect 15436 14288 15442 14340
rect 15565 14331 15623 14337
rect 15565 14297 15577 14331
rect 15611 14328 15623 14331
rect 16298 14328 16304 14340
rect 15611 14300 16304 14328
rect 15611 14297 15623 14300
rect 15565 14291 15623 14297
rect 16298 14288 16304 14300
rect 16356 14288 16362 14340
rect 16574 14288 16580 14340
rect 16632 14328 16638 14340
rect 17236 14328 17264 14359
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 18414 14396 18420 14408
rect 18375 14368 18420 14396
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 17770 14328 17776 14340
rect 16632 14300 17776 14328
rect 16632 14288 16638 14300
rect 17770 14288 17776 14300
rect 17828 14328 17834 14340
rect 17828 14300 18368 14328
rect 17828 14288 17834 14300
rect 2924 14232 3556 14260
rect 2924 14220 2930 14232
rect 3602 14220 3608 14272
rect 3660 14260 3666 14272
rect 4065 14263 4123 14269
rect 4065 14260 4077 14263
rect 3660 14232 4077 14260
rect 3660 14220 3666 14232
rect 4065 14229 4077 14232
rect 4111 14229 4123 14263
rect 6086 14260 6092 14272
rect 6047 14232 6092 14260
rect 4065 14223 4123 14229
rect 6086 14220 6092 14232
rect 6144 14220 6150 14272
rect 7374 14220 7380 14272
rect 7432 14260 7438 14272
rect 8021 14263 8079 14269
rect 8021 14260 8033 14263
rect 7432 14232 8033 14260
rect 7432 14220 7438 14232
rect 8021 14229 8033 14232
rect 8067 14229 8079 14263
rect 8662 14260 8668 14272
rect 8623 14232 8668 14260
rect 8021 14223 8079 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 13814 14260 13820 14272
rect 13775 14232 13820 14260
rect 13814 14220 13820 14232
rect 13872 14220 13878 14272
rect 14274 14220 14280 14272
rect 14332 14220 14338 14272
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 14829 14263 14887 14269
rect 14829 14260 14841 14263
rect 14516 14232 14841 14260
rect 14516 14220 14522 14232
rect 14829 14229 14841 14232
rect 14875 14229 14887 14263
rect 18340 14260 18368 14300
rect 19794 14260 19800 14272
rect 18340 14232 19800 14260
rect 14829 14223 14887 14229
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1765 14059 1823 14065
rect 1765 14025 1777 14059
rect 1811 14056 1823 14059
rect 2774 14056 2780 14068
rect 1811 14028 2780 14056
rect 1811 14025 1823 14028
rect 1765 14019 1823 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 3145 14059 3203 14065
rect 3145 14025 3157 14059
rect 3191 14056 3203 14059
rect 3326 14056 3332 14068
rect 3191 14028 3332 14056
rect 3191 14025 3203 14028
rect 3145 14019 3203 14025
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 3252 13929 3280 14028
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 3789 14059 3847 14065
rect 3789 14025 3801 14059
rect 3835 14056 3847 14059
rect 4154 14056 4160 14068
rect 3835 14028 4160 14056
rect 3835 14025 3847 14028
rect 3789 14019 3847 14025
rect 4154 14016 4160 14028
rect 4212 14056 4218 14068
rect 5718 14056 5724 14068
rect 4212 14028 5304 14056
rect 5679 14028 5724 14056
rect 4212 14016 4218 14028
rect 5276 14000 5304 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 6914 14056 6920 14068
rect 6104 14028 6920 14056
rect 5258 13988 5264 14000
rect 5219 13960 5264 13988
rect 5258 13948 5264 13960
rect 5316 13948 5322 14000
rect 5629 13991 5687 13997
rect 5629 13957 5641 13991
rect 5675 13988 5687 13991
rect 6104 13988 6132 14028
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 10134 14056 10140 14068
rect 9815 14028 10140 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 10134 14016 10140 14028
rect 10192 14056 10198 14068
rect 10413 14059 10471 14065
rect 10413 14056 10425 14059
rect 10192 14028 10425 14056
rect 10192 14016 10198 14028
rect 10413 14025 10425 14028
rect 10459 14025 10471 14059
rect 13814 14056 13820 14068
rect 10413 14019 10471 14025
rect 13556 14028 13820 14056
rect 6825 13991 6883 13997
rect 6825 13988 6837 13991
rect 5675 13960 6132 13988
rect 6196 13960 6837 13988
rect 5675 13957 5687 13960
rect 5629 13951 5687 13957
rect 2317 13923 2375 13929
rect 2317 13920 2329 13923
rect 1452 13892 2329 13920
rect 1452 13880 1458 13892
rect 2317 13889 2329 13892
rect 2363 13920 2375 13923
rect 3237 13923 3295 13929
rect 2363 13892 2728 13920
rect 2363 13889 2375 13892
rect 2317 13883 2375 13889
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 2590 13852 2596 13864
rect 2179 13824 2596 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 2700 13852 2728 13892
rect 3237 13889 3249 13923
rect 3283 13889 3295 13923
rect 3237 13883 3295 13889
rect 3694 13852 3700 13864
rect 2700 13824 3700 13852
rect 3694 13812 3700 13824
rect 3752 13812 3758 13864
rect 4154 13861 4160 13864
rect 3881 13855 3939 13861
rect 3881 13821 3893 13855
rect 3927 13821 3939 13855
rect 4148 13852 4160 13861
rect 4115 13824 4160 13852
rect 3881 13815 3939 13821
rect 4148 13815 4160 13824
rect 3896 13784 3924 13815
rect 4154 13812 4160 13815
rect 4212 13812 4218 13864
rect 5902 13812 5908 13864
rect 5960 13852 5966 13864
rect 6196 13861 6224 13960
rect 6825 13957 6837 13960
rect 6871 13957 6883 13991
rect 13556 13988 13584 14028
rect 13814 14016 13820 14028
rect 13872 14056 13878 14068
rect 20165 14059 20223 14065
rect 20165 14056 20177 14059
rect 13872 14028 20177 14056
rect 13872 14016 13878 14028
rect 20165 14025 20177 14028
rect 20211 14025 20223 14059
rect 20165 14019 20223 14025
rect 6825 13951 6883 13957
rect 13464 13960 13584 13988
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 7374 13920 7380 13932
rect 6328 13892 6373 13920
rect 7335 13892 7380 13920
rect 6328 13880 6334 13892
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 13464 13929 13492 13960
rect 15654 13948 15660 14000
rect 15712 13988 15718 14000
rect 15933 13991 15991 13997
rect 15933 13988 15945 13991
rect 15712 13960 15945 13988
rect 15712 13948 15718 13960
rect 15933 13957 15945 13960
rect 15979 13957 15991 13991
rect 15933 13951 15991 13957
rect 18598 13948 18604 14000
rect 18656 13988 18662 14000
rect 19426 13988 19432 14000
rect 18656 13960 19196 13988
rect 19387 13960 19432 13988
rect 18656 13948 18662 13960
rect 13449 13923 13507 13929
rect 13449 13889 13461 13923
rect 13495 13889 13507 13923
rect 13449 13883 13507 13889
rect 13633 13923 13691 13929
rect 13633 13889 13645 13923
rect 13679 13920 13691 13923
rect 18693 13923 18751 13929
rect 18693 13920 18705 13923
rect 13679 13892 13768 13920
rect 13679 13889 13691 13892
rect 13633 13883 13691 13889
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 5960 13824 6193 13852
rect 5960 13812 5966 13824
rect 6181 13821 6193 13824
rect 6227 13821 6239 13855
rect 7190 13852 7196 13864
rect 7103 13824 7196 13852
rect 6181 13815 6239 13821
rect 7190 13812 7196 13824
rect 7248 13852 7254 13864
rect 7558 13852 7564 13864
rect 7248 13824 7564 13852
rect 7248 13812 7254 13824
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 8389 13855 8447 13861
rect 8389 13821 8401 13855
rect 8435 13852 8447 13855
rect 8478 13852 8484 13864
rect 8435 13824 8484 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 8662 13861 8668 13864
rect 8656 13852 8668 13861
rect 8623 13824 8668 13852
rect 8656 13815 8668 13824
rect 8720 13852 8726 13864
rect 9582 13852 9588 13864
rect 8720 13824 9588 13852
rect 8662 13812 8668 13815
rect 8720 13812 8726 13824
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 10594 13852 10600 13864
rect 10555 13824 10600 13852
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 10864 13855 10922 13861
rect 10864 13821 10876 13855
rect 10910 13852 10922 13855
rect 11146 13852 11152 13864
rect 10910 13824 11152 13852
rect 10910 13821 10922 13824
rect 10864 13815 10922 13821
rect 11146 13812 11152 13824
rect 11204 13852 11210 13864
rect 12342 13852 12348 13864
rect 11204 13824 12348 13852
rect 11204 13812 11210 13824
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 4798 13784 4804 13796
rect 3896 13756 4804 13784
rect 4798 13744 4804 13756
rect 4856 13744 4862 13796
rect 6086 13784 6092 13796
rect 5999 13756 6092 13784
rect 6086 13744 6092 13756
rect 6144 13784 6150 13796
rect 7837 13787 7895 13793
rect 7837 13784 7849 13787
rect 6144 13756 7849 13784
rect 6144 13744 6150 13756
rect 7837 13753 7849 13756
rect 7883 13753 7895 13787
rect 7837 13747 7895 13753
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 10686 13784 10692 13796
rect 9824 13756 10692 13784
rect 9824 13744 9830 13756
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 13740 13784 13768 13892
rect 17880 13892 18705 13920
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13872 13824 14013 13852
rect 13872 13812 13878 13824
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 16301 13855 16359 13861
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 16390 13852 16396 13864
rect 16347 13824 16396 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 16574 13861 16580 13864
rect 16568 13852 16580 13861
rect 16535 13824 16580 13852
rect 16568 13815 16580 13824
rect 16574 13812 16580 13815
rect 16632 13812 16638 13864
rect 14268 13787 14326 13793
rect 14268 13784 14280 13787
rect 13740 13756 14280 13784
rect 14268 13753 14280 13756
rect 14314 13784 14326 13787
rect 14366 13784 14372 13796
rect 14314 13756 14372 13784
rect 14314 13753 14326 13756
rect 14268 13747 14326 13753
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 7285 13719 7343 13725
rect 7285 13685 7297 13719
rect 7331 13716 7343 13719
rect 7742 13716 7748 13728
rect 7331 13688 7748 13716
rect 7331 13685 7343 13688
rect 7285 13679 7343 13685
rect 7742 13676 7748 13688
rect 7800 13676 7806 13728
rect 9674 13676 9680 13728
rect 9732 13716 9738 13728
rect 10045 13719 10103 13725
rect 10045 13716 10057 13719
rect 9732 13688 10057 13716
rect 9732 13676 9738 13688
rect 10045 13685 10057 13688
rect 10091 13685 10103 13719
rect 11974 13716 11980 13728
rect 11935 13688 11980 13716
rect 10045 13679 10103 13685
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 12894 13716 12900 13728
rect 12855 13688 12900 13716
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 12989 13719 13047 13725
rect 12989 13685 13001 13719
rect 13035 13716 13047 13719
rect 13262 13716 13268 13728
rect 13035 13688 13268 13716
rect 13035 13685 13047 13688
rect 12989 13679 13047 13685
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 13357 13719 13415 13725
rect 13357 13685 13369 13719
rect 13403 13716 13415 13719
rect 13722 13716 13728 13728
rect 13403 13688 13728 13716
rect 13403 13685 13415 13688
rect 13357 13679 13415 13685
rect 13722 13676 13728 13688
rect 13780 13676 13786 13728
rect 15378 13716 15384 13728
rect 15339 13688 15384 13716
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 17678 13716 17684 13728
rect 17591 13688 17684 13716
rect 17678 13676 17684 13688
rect 17736 13716 17742 13728
rect 17880 13716 17908 13892
rect 18693 13889 18705 13892
rect 18739 13920 18751 13923
rect 18966 13920 18972 13932
rect 18739 13892 18972 13920
rect 18739 13889 18751 13892
rect 18693 13883 18751 13889
rect 18966 13880 18972 13892
rect 19024 13880 19030 13932
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18417 13855 18475 13861
rect 18417 13852 18429 13855
rect 18012 13824 18429 13852
rect 18012 13812 18018 13824
rect 18417 13821 18429 13824
rect 18463 13852 18475 13855
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 18463 13824 19073 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19168 13852 19196 13960
rect 19426 13948 19432 13960
rect 19484 13948 19490 14000
rect 19794 13988 19800 14000
rect 19755 13960 19800 13988
rect 19794 13948 19800 13960
rect 19852 13948 19858 14000
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 20533 13923 20591 13929
rect 20533 13920 20545 13923
rect 19300 13892 20545 13920
rect 19300 13880 19306 13892
rect 20533 13889 20545 13892
rect 20579 13889 20591 13923
rect 20533 13883 20591 13889
rect 20901 13855 20959 13861
rect 20901 13852 20913 13855
rect 19168 13824 20913 13852
rect 19061 13815 19119 13821
rect 20901 13821 20913 13824
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 18506 13784 18512 13796
rect 18467 13756 18512 13784
rect 18506 13744 18512 13756
rect 18564 13744 18570 13796
rect 17736 13688 17908 13716
rect 18049 13719 18107 13725
rect 17736 13676 17742 13688
rect 18049 13685 18061 13719
rect 18095 13716 18107 13719
rect 19150 13716 19156 13728
rect 18095 13688 19156 13716
rect 18095 13685 18107 13688
rect 18049 13679 18107 13685
rect 19150 13676 19156 13688
rect 19208 13676 19214 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 2777 13515 2835 13521
rect 2777 13481 2789 13515
rect 2823 13512 2835 13515
rect 2866 13512 2872 13524
rect 2823 13484 2872 13512
rect 2823 13481 2835 13484
rect 2777 13475 2835 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 4433 13515 4491 13521
rect 4433 13481 4445 13515
rect 4479 13512 4491 13515
rect 4706 13512 4712 13524
rect 4479 13484 4712 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 4706 13472 4712 13484
rect 4764 13512 4770 13524
rect 5350 13512 5356 13524
rect 4764 13484 5356 13512
rect 4764 13472 4770 13484
rect 5350 13472 5356 13484
rect 5408 13512 5414 13524
rect 7190 13512 7196 13524
rect 5408 13484 7196 13512
rect 5408 13472 5414 13484
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7282 13472 7288 13524
rect 7340 13512 7346 13524
rect 8202 13512 8208 13524
rect 7340 13484 8208 13512
rect 7340 13472 7346 13484
rect 8202 13472 8208 13484
rect 8260 13512 8266 13524
rect 8297 13515 8355 13521
rect 8297 13512 8309 13515
rect 8260 13484 8309 13512
rect 8260 13472 8266 13484
rect 8297 13481 8309 13484
rect 8343 13481 8355 13515
rect 8297 13475 8355 13481
rect 9033 13515 9091 13521
rect 9033 13481 9045 13515
rect 9079 13512 9091 13515
rect 9766 13512 9772 13524
rect 9079 13484 9772 13512
rect 9079 13481 9091 13484
rect 9033 13475 9091 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 13446 13512 13452 13524
rect 10520 13484 13452 13512
rect 1578 13404 1584 13456
rect 1636 13444 1642 13456
rect 10520 13453 10548 13484
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 13688 13484 13952 13512
rect 13688 13472 13694 13484
rect 2225 13447 2283 13453
rect 2225 13444 2237 13447
rect 1636 13416 2237 13444
rect 1636 13404 1642 13416
rect 2225 13413 2237 13416
rect 2271 13413 2283 13447
rect 2225 13407 2283 13413
rect 9953 13447 10011 13453
rect 9953 13413 9965 13447
rect 9999 13444 10011 13447
rect 10505 13447 10563 13453
rect 10505 13444 10517 13447
rect 9999 13416 10517 13444
rect 9999 13413 10011 13416
rect 9953 13407 10011 13413
rect 10505 13413 10517 13416
rect 10551 13413 10563 13447
rect 13078 13444 13084 13456
rect 10505 13407 10563 13413
rect 12452 13416 13084 13444
rect 1394 13376 1400 13388
rect 1355 13348 1400 13376
rect 1394 13336 1400 13348
rect 1452 13336 1458 13388
rect 1670 13336 1676 13388
rect 1728 13376 1734 13388
rect 1946 13376 1952 13388
rect 1728 13348 1952 13376
rect 1728 13336 1734 13348
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13376 3571 13379
rect 4154 13376 4160 13388
rect 3559 13348 4160 13376
rect 3559 13345 3571 13348
rect 3513 13339 3571 13345
rect 4154 13336 4160 13348
rect 4212 13376 4218 13388
rect 5166 13385 5172 13388
rect 5160 13376 5172 13385
rect 4212 13348 5172 13376
rect 4212 13336 4218 13348
rect 5160 13339 5172 13348
rect 5166 13336 5172 13339
rect 5224 13336 5230 13388
rect 6897 13379 6955 13385
rect 6897 13376 6909 13379
rect 6196 13348 6909 13376
rect 3418 13308 3424 13320
rect 1596 13280 3424 13308
rect 1596 13249 1624 13280
rect 3418 13268 3424 13280
rect 3476 13268 3482 13320
rect 4890 13308 4896 13320
rect 4851 13280 4896 13308
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 1581 13243 1639 13249
rect 1581 13209 1593 13243
rect 1627 13209 1639 13243
rect 1581 13203 1639 13209
rect 3145 13243 3203 13249
rect 3145 13209 3157 13243
rect 3191 13240 3203 13243
rect 4798 13240 4804 13252
rect 3191 13212 4804 13240
rect 3191 13209 3203 13212
rect 3145 13203 3203 13209
rect 4798 13200 4804 13212
rect 4856 13200 4862 13252
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 6086 13172 6092 13184
rect 3927 13144 6092 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 6086 13132 6092 13144
rect 6144 13172 6150 13184
rect 6196 13172 6224 13348
rect 6897 13345 6909 13348
rect 6943 13376 6955 13379
rect 7374 13376 7380 13388
rect 6943 13348 7380 13376
rect 6943 13345 6955 13348
rect 6897 13339 6955 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 8481 13379 8539 13385
rect 8481 13345 8493 13379
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 6362 13308 6368 13320
rect 6288 13280 6368 13308
rect 6288 13249 6316 13280
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 6638 13308 6644 13320
rect 6599 13280 6644 13308
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 6273 13243 6331 13249
rect 6273 13209 6285 13243
rect 6319 13209 6331 13243
rect 8496 13240 8524 13339
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8904 13348 8953 13376
rect 8904 13336 8910 13348
rect 8941 13345 8953 13348
rect 8987 13376 8999 13379
rect 9490 13376 9496 13388
rect 8987 13348 9496 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 12452 13376 12480 13416
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 13532 13447 13590 13453
rect 13532 13413 13544 13447
rect 13578 13444 13590 13447
rect 13722 13444 13728 13456
rect 13578 13416 13728 13444
rect 13578 13413 13590 13416
rect 13532 13407 13590 13413
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 9631 13348 12480 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 12526 13336 12532 13388
rect 12584 13376 12590 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12584 13348 12725 13376
rect 12584 13336 12590 13348
rect 12713 13345 12725 13348
rect 12759 13376 12771 13379
rect 13170 13376 13176 13388
rect 12759 13348 13176 13376
rect 12759 13345 12771 13348
rect 12713 13339 12771 13345
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 13814 13376 13820 13388
rect 13280 13348 13820 13376
rect 13280 13320 13308 13348
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 13924 13376 13952 13484
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 14424 13484 14657 13512
rect 14424 13472 14430 13484
rect 14645 13481 14657 13484
rect 14691 13481 14703 13515
rect 14645 13475 14703 13481
rect 14660 13444 14688 13475
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15436 13484 16313 13512
rect 15436 13472 15442 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16942 13512 16948 13524
rect 16903 13484 16948 13512
rect 16301 13475 16359 13481
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 18782 13512 18788 13524
rect 18743 13484 18788 13512
rect 18782 13472 18788 13484
rect 18840 13472 18846 13524
rect 18874 13472 18880 13524
rect 18932 13512 18938 13524
rect 20533 13515 20591 13521
rect 20533 13512 20545 13515
rect 18932 13484 20545 13512
rect 18932 13472 18938 13484
rect 20533 13481 20545 13484
rect 20579 13481 20591 13515
rect 20533 13475 20591 13481
rect 15562 13444 15568 13456
rect 14660 13416 15568 13444
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 15930 13444 15936 13456
rect 15891 13416 15936 13444
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 17304 13447 17362 13453
rect 17304 13413 17316 13447
rect 17350 13444 17362 13447
rect 17678 13444 17684 13456
rect 17350 13416 17684 13444
rect 17350 13413 17362 13416
rect 17304 13407 17362 13413
rect 17678 13404 17684 13416
rect 17736 13404 17742 13456
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 20165 13447 20223 13453
rect 20165 13444 20177 13447
rect 18564 13416 20177 13444
rect 18564 13404 18570 13416
rect 20165 13413 20177 13416
rect 20211 13413 20223 13447
rect 20165 13407 20223 13413
rect 19429 13379 19487 13385
rect 19429 13376 19441 13379
rect 13924 13348 19441 13376
rect 19429 13345 19441 13348
rect 19475 13345 19487 13379
rect 19429 13339 19487 13345
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9674 13308 9680 13320
rect 9263 13280 9680 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13308 10103 13311
rect 10134 13308 10140 13320
rect 10091 13280 10140 13308
rect 10091 13277 10103 13280
rect 10045 13271 10103 13277
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 12805 13311 12863 13317
rect 12805 13308 12817 13311
rect 12676 13280 12817 13308
rect 12676 13268 12682 13280
rect 12805 13277 12817 13280
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13078 13308 13084 13320
rect 13035 13280 13084 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 11790 13240 11796 13252
rect 8496 13212 11796 13240
rect 6273 13203 6331 13209
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 11974 13200 11980 13252
rect 12032 13240 12038 13252
rect 13004 13240 13032 13271
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 13262 13308 13268 13320
rect 13223 13280 13268 13308
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 14458 13268 14464 13320
rect 14516 13308 14522 13320
rect 14921 13311 14979 13317
rect 14921 13308 14933 13311
rect 14516 13280 14933 13308
rect 14516 13268 14522 13280
rect 14921 13277 14933 13280
rect 14967 13277 14979 13311
rect 14921 13271 14979 13277
rect 15654 13268 15660 13320
rect 15712 13308 15718 13320
rect 17037 13311 17095 13317
rect 17037 13308 17049 13311
rect 15712 13280 17049 13308
rect 15712 13268 15718 13280
rect 17037 13277 17049 13280
rect 17083 13277 17095 13311
rect 17037 13271 17095 13277
rect 18690 13268 18696 13320
rect 18748 13308 18754 13320
rect 19150 13308 19156 13320
rect 18748 13280 19156 13308
rect 18748 13268 18754 13280
rect 19150 13268 19156 13280
rect 19208 13308 19214 13320
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 19208 13280 21097 13308
rect 19208 13268 19214 13280
rect 21085 13277 21097 13280
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 12032 13212 13032 13240
rect 12032 13200 12038 13212
rect 6144 13144 6224 13172
rect 6144 13132 6150 13144
rect 6362 13132 6368 13184
rect 6420 13172 6426 13184
rect 8021 13175 8079 13181
rect 8021 13172 8033 13175
rect 6420 13144 8033 13172
rect 6420 13132 6426 13144
rect 8021 13141 8033 13144
rect 8067 13141 8079 13175
rect 8021 13135 8079 13141
rect 8573 13175 8631 13181
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 8662 13172 8668 13184
rect 8619 13144 8668 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 8812 13144 9505 13172
rect 8812 13132 8818 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9493 13135 9551 13141
rect 12345 13175 12403 13181
rect 12345 13141 12357 13175
rect 12391 13172 12403 13175
rect 12710 13172 12716 13184
rect 12391 13144 12716 13172
rect 12391 13141 12403 13144
rect 12345 13135 12403 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 14476 13172 14504 13268
rect 16574 13200 16580 13252
rect 16632 13240 16638 13252
rect 16942 13240 16948 13252
rect 16632 13212 16948 13240
rect 16632 13200 16638 13212
rect 16942 13200 16948 13212
rect 17000 13200 17006 13252
rect 18046 13200 18052 13252
rect 18104 13240 18110 13252
rect 19797 13243 19855 13249
rect 19797 13240 19809 13243
rect 18104 13212 19809 13240
rect 18104 13200 18110 13212
rect 19797 13209 19809 13212
rect 19843 13209 19855 13243
rect 19797 13203 19855 13209
rect 13688 13144 14504 13172
rect 13688 13132 13694 13144
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 14884 13144 15485 13172
rect 14884 13132 14890 13144
rect 15473 13141 15485 13144
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 18417 13175 18475 13181
rect 18417 13141 18429 13175
rect 18463 13172 18475 13175
rect 18598 13172 18604 13184
rect 18463 13144 18604 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 19058 13172 19064 13184
rect 19019 13144 19064 13172
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 1854 12968 1860 12980
rect 1719 12940 1860 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 4706 12968 4712 12980
rect 4540 12940 4712 12968
rect 1394 12792 1400 12844
rect 1452 12832 1458 12844
rect 1578 12832 1584 12844
rect 1452 12804 1584 12832
rect 1452 12792 1458 12804
rect 1578 12792 1584 12804
rect 1636 12832 1642 12844
rect 2225 12835 2283 12841
rect 2225 12832 2237 12835
rect 1636 12804 2237 12832
rect 1636 12792 1642 12804
rect 2225 12801 2237 12804
rect 2271 12801 2283 12835
rect 2225 12795 2283 12801
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 4154 12832 4160 12844
rect 3099 12804 4160 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4540 12841 4568 12940
rect 4706 12928 4712 12940
rect 4764 12968 4770 12980
rect 4890 12968 4896 12980
rect 4764 12940 4896 12968
rect 4764 12928 4770 12940
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5224 12940 5917 12968
rect 5224 12928 5230 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 9214 12968 9220 12980
rect 5905 12931 5963 12937
rect 8220 12940 9220 12968
rect 5534 12860 5540 12912
rect 5592 12900 5598 12912
rect 8220 12900 8248 12940
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 9582 12968 9588 12980
rect 9543 12940 9588 12968
rect 9582 12928 9588 12940
rect 9640 12928 9646 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 13725 12971 13783 12977
rect 13725 12968 13737 12971
rect 11848 12940 13737 12968
rect 11848 12928 11854 12940
rect 13725 12937 13737 12940
rect 13771 12937 13783 12971
rect 13725 12931 13783 12937
rect 13817 12971 13875 12977
rect 13817 12937 13829 12971
rect 13863 12968 13875 12971
rect 14274 12968 14280 12980
rect 13863 12940 14280 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 16761 12971 16819 12977
rect 16761 12968 16773 12971
rect 15620 12940 16773 12968
rect 15620 12928 15626 12940
rect 16761 12937 16773 12940
rect 16807 12968 16819 12971
rect 17129 12971 17187 12977
rect 17129 12968 17141 12971
rect 16807 12940 17141 12968
rect 16807 12937 16819 12940
rect 16761 12931 16819 12937
rect 17129 12937 17141 12940
rect 17175 12937 17187 12971
rect 17129 12931 17187 12937
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18506 12968 18512 12980
rect 18095 12940 18512 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 19058 12968 19064 12980
rect 19019 12940 19064 12968
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 5592 12872 8248 12900
rect 5592 12860 5598 12872
rect 9490 12860 9496 12912
rect 9548 12900 9554 12912
rect 9861 12903 9919 12909
rect 9861 12900 9873 12903
rect 9548 12872 9873 12900
rect 9548 12860 9554 12872
rect 9861 12869 9873 12872
rect 9907 12869 9919 12903
rect 9861 12863 9919 12869
rect 13449 12903 13507 12909
rect 13449 12869 13461 12903
rect 13495 12900 13507 12903
rect 13906 12900 13912 12912
rect 13495 12872 13912 12900
rect 13495 12869 13507 12872
rect 13449 12863 13507 12869
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 20165 12903 20223 12909
rect 20165 12900 20177 12903
rect 14292 12872 20177 12900
rect 14292 12844 14320 12872
rect 20165 12869 20177 12872
rect 20211 12869 20223 12903
rect 20165 12863 20223 12869
rect 4525 12835 4583 12841
rect 4525 12832 4537 12835
rect 4304 12804 4537 12832
rect 4304 12792 4310 12804
rect 4525 12801 4537 12804
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12832 7711 12835
rect 7699 12804 8340 12832
rect 7699 12801 7711 12804
rect 7653 12795 7711 12801
rect 1486 12764 1492 12776
rect 1447 12736 1492 12764
rect 1486 12724 1492 12736
rect 1544 12724 1550 12776
rect 2038 12764 2044 12776
rect 1999 12736 2044 12764
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12764 3479 12767
rect 6181 12767 6239 12773
rect 6181 12764 6193 12767
rect 3467 12736 3924 12764
rect 3467 12733 3479 12736
rect 3421 12727 3479 12733
rect 1394 12656 1400 12708
rect 1452 12696 1458 12708
rect 2130 12696 2136 12708
rect 1452 12668 2136 12696
rect 1452 12656 1458 12668
rect 2130 12656 2136 12668
rect 2188 12656 2194 12708
rect 3896 12705 3924 12736
rect 4632 12736 6193 12764
rect 3881 12699 3939 12705
rect 3881 12665 3893 12699
rect 3927 12696 3939 12699
rect 4632 12696 4660 12736
rect 6181 12733 6193 12736
rect 6227 12733 6239 12767
rect 6181 12727 6239 12733
rect 7558 12724 7564 12776
rect 7616 12764 7622 12776
rect 8205 12767 8263 12773
rect 8205 12764 8217 12767
rect 7616 12736 8217 12764
rect 7616 12724 7622 12736
rect 8205 12733 8217 12736
rect 8251 12733 8263 12767
rect 8312 12764 8340 12804
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 10192 12804 10609 12832
rect 10192 12792 10198 12804
rect 10597 12801 10609 12804
rect 10643 12832 10655 12835
rect 10643 12804 10824 12832
rect 10643 12801 10655 12804
rect 10597 12795 10655 12801
rect 8461 12767 8519 12773
rect 8461 12764 8473 12767
rect 8312 12736 8473 12764
rect 8205 12727 8263 12733
rect 8461 12733 8473 12736
rect 8507 12764 8519 12767
rect 9674 12764 9680 12776
rect 8507 12736 9680 12764
rect 8507 12733 8519 12736
rect 8461 12727 8519 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12733 10747 12767
rect 10796 12764 10824 12804
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 12434 12832 12440 12844
rect 11848 12804 12440 12832
rect 11848 12792 11854 12804
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 13078 12832 13084 12844
rect 12991 12804 13084 12832
rect 13078 12792 13084 12804
rect 13136 12832 13142 12844
rect 14274 12832 14280 12844
rect 13136 12804 13575 12832
rect 14187 12804 14280 12832
rect 13136 12792 13142 12804
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 10796 12736 12817 12764
rect 10689 12727 10747 12733
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 4798 12705 4804 12708
rect 4792 12696 4804 12705
rect 3927 12668 4660 12696
rect 4759 12668 4804 12696
rect 3927 12665 3939 12668
rect 3881 12659 3939 12665
rect 4792 12659 4804 12668
rect 4856 12696 4862 12708
rect 5534 12696 5540 12708
rect 4856 12668 5540 12696
rect 4798 12656 4804 12659
rect 4856 12656 4862 12668
rect 5534 12656 5540 12668
rect 5592 12656 5598 12708
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 3513 12631 3571 12637
rect 3513 12628 3525 12631
rect 2096 12600 3525 12628
rect 2096 12588 2102 12600
rect 3513 12597 3525 12600
rect 3559 12597 3571 12631
rect 3513 12591 3571 12597
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 5074 12628 5080 12640
rect 4019 12600 5080 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 7190 12628 7196 12640
rect 7151 12600 7196 12628
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 7745 12631 7803 12637
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 8570 12628 8576 12640
rect 7791 12600 8576 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 10704 12628 10732 12727
rect 10956 12699 11014 12705
rect 10956 12665 10968 12699
rect 11002 12696 11014 12699
rect 11974 12696 11980 12708
rect 11002 12668 11980 12696
rect 11002 12665 11014 12668
rect 10956 12659 11014 12665
rect 11974 12656 11980 12668
rect 12032 12656 12038 12708
rect 11698 12628 11704 12640
rect 10704 12600 11704 12628
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 12250 12628 12256 12640
rect 12115 12600 12256 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12894 12628 12900 12640
rect 12492 12600 12537 12628
rect 12855 12600 12900 12628
rect 12492 12588 12498 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 13547 12628 13575 12804
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 14366 12792 14372 12844
rect 14424 12832 14430 12844
rect 14826 12832 14832 12844
rect 14424 12804 14469 12832
rect 14787 12804 14832 12832
rect 14424 12792 14430 12804
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 18693 12835 18751 12841
rect 18693 12801 18705 12835
rect 18739 12832 18751 12835
rect 19426 12832 19432 12844
rect 18739 12804 19432 12832
rect 18739 12801 18751 12804
rect 18693 12795 18751 12801
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 13725 12767 13783 12773
rect 13725 12764 13737 12767
rect 13679 12736 13737 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 13725 12733 13737 12736
rect 13771 12733 13783 12767
rect 13725 12727 13783 12733
rect 14185 12767 14243 12773
rect 14185 12733 14197 12767
rect 14231 12764 14243 12767
rect 14844 12764 14872 12792
rect 14231 12736 14872 12764
rect 14231 12733 14243 12736
rect 14185 12727 14243 12733
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15381 12767 15439 12773
rect 15381 12764 15393 12767
rect 15252 12736 15393 12764
rect 15252 12724 15258 12736
rect 15381 12733 15393 12736
rect 15427 12764 15439 12767
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 15427 12736 15761 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 15749 12733 15761 12736
rect 15795 12764 15807 12767
rect 17586 12764 17592 12776
rect 15795 12736 17592 12764
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 17586 12724 17592 12736
rect 17644 12724 17650 12776
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 18417 12767 18475 12773
rect 18417 12764 18429 12767
rect 18012 12736 18429 12764
rect 18012 12724 18018 12736
rect 18417 12733 18429 12736
rect 18463 12764 18475 12767
rect 20901 12767 20959 12773
rect 20901 12764 20913 12767
rect 18463 12736 20913 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 20901 12733 20913 12736
rect 20947 12733 20959 12767
rect 20901 12727 20959 12733
rect 13906 12656 13912 12708
rect 13964 12696 13970 12708
rect 14550 12696 14556 12708
rect 13964 12668 14556 12696
rect 13964 12656 13970 12668
rect 14550 12656 14556 12668
rect 14608 12656 14614 12708
rect 18506 12696 18512 12708
rect 14660 12668 17724 12696
rect 18419 12668 18512 12696
rect 14660 12628 14688 12668
rect 13547 12600 14688 12628
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15068 12600 16129 12628
rect 15068 12588 15074 12600
rect 16117 12597 16129 12600
rect 16163 12628 16175 12631
rect 16485 12631 16543 12637
rect 16485 12628 16497 12631
rect 16163 12600 16497 12628
rect 16163 12597 16175 12600
rect 16117 12591 16175 12597
rect 16485 12597 16497 12600
rect 16531 12628 16543 12631
rect 17126 12628 17132 12640
rect 16531 12600 17132 12628
rect 16531 12597 16543 12600
rect 16485 12591 16543 12597
rect 17126 12588 17132 12600
rect 17184 12588 17190 12640
rect 17586 12628 17592 12640
rect 17547 12600 17592 12628
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 17696 12628 17724 12668
rect 18506 12656 18512 12668
rect 18564 12696 18570 12708
rect 20533 12699 20591 12705
rect 20533 12696 20545 12699
rect 18564 12668 20545 12696
rect 18564 12656 18570 12668
rect 20533 12665 20545 12668
rect 20579 12665 20591 12699
rect 20533 12659 20591 12665
rect 19797 12631 19855 12637
rect 19797 12628 19809 12631
rect 17696 12600 19809 12628
rect 19797 12597 19809 12600
rect 19843 12597 19855 12631
rect 19797 12591 19855 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1762 12424 1768 12436
rect 1723 12396 1768 12424
rect 1762 12384 1768 12396
rect 1820 12384 1826 12436
rect 2958 12384 2964 12436
rect 3016 12424 3022 12436
rect 3053 12427 3111 12433
rect 3053 12424 3065 12427
rect 3016 12396 3065 12424
rect 3016 12384 3022 12396
rect 3053 12393 3065 12396
rect 3099 12393 3111 12427
rect 5537 12427 5595 12433
rect 5537 12424 5549 12427
rect 3053 12387 3111 12393
rect 3988 12396 5549 12424
rect 1946 12316 1952 12368
rect 2004 12356 2010 12368
rect 3988 12356 4016 12396
rect 5537 12393 5549 12396
rect 5583 12393 5595 12427
rect 5537 12387 5595 12393
rect 5813 12427 5871 12433
rect 5813 12393 5825 12427
rect 5859 12424 5871 12427
rect 6270 12424 6276 12436
rect 5859 12396 6276 12424
rect 5859 12393 5871 12396
rect 5813 12387 5871 12393
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 8846 12424 8852 12436
rect 6420 12396 8852 12424
rect 6420 12384 6426 12396
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 9309 12427 9367 12433
rect 9309 12393 9321 12427
rect 9355 12424 9367 12427
rect 9766 12424 9772 12436
rect 9355 12396 9772 12424
rect 9355 12393 9367 12396
rect 9309 12387 9367 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11882 12424 11888 12436
rect 11112 12396 11888 12424
rect 11112 12384 11118 12396
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12424 13783 12427
rect 14274 12424 14280 12436
rect 13771 12396 14280 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 16758 12384 16764 12436
rect 16816 12424 16822 12436
rect 16853 12427 16911 12433
rect 16853 12424 16865 12427
rect 16816 12396 16865 12424
rect 16816 12384 16822 12396
rect 16853 12393 16865 12396
rect 16899 12393 16911 12427
rect 16853 12387 16911 12393
rect 17126 12384 17132 12436
rect 17184 12424 17190 12436
rect 17497 12427 17555 12433
rect 17184 12396 17448 12424
rect 17184 12384 17190 12396
rect 2004 12328 4016 12356
rect 2004 12316 2010 12328
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 12894 12356 12900 12368
rect 4120 12328 12900 12356
rect 4120 12316 4126 12328
rect 12894 12316 12900 12328
rect 12952 12316 12958 12368
rect 13630 12316 13636 12368
rect 13688 12356 13694 12368
rect 14185 12359 14243 12365
rect 14185 12356 14197 12359
rect 13688 12328 14197 12356
rect 13688 12316 13694 12328
rect 14185 12325 14197 12328
rect 14231 12356 14243 12359
rect 15194 12356 15200 12368
rect 14231 12328 15200 12356
rect 14231 12325 14243 12328
rect 14185 12319 14243 12325
rect 15194 12316 15200 12328
rect 15252 12316 15258 12368
rect 17420 12356 17448 12396
rect 17497 12393 17509 12427
rect 17543 12424 17555 12427
rect 18506 12424 18512 12436
rect 17543 12396 18512 12424
rect 17543 12393 17555 12396
rect 17497 12387 17555 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 20533 12427 20591 12433
rect 20533 12393 20545 12427
rect 20579 12393 20591 12427
rect 20533 12387 20591 12393
rect 21177 12427 21235 12433
rect 21177 12393 21189 12427
rect 21223 12424 21235 12427
rect 21358 12424 21364 12436
rect 21223 12396 21364 12424
rect 21223 12393 21235 12396
rect 21177 12387 21235 12393
rect 20548 12356 20576 12387
rect 21358 12384 21364 12396
rect 21416 12384 21422 12436
rect 17420 12328 20576 12356
rect 1581 12291 1639 12297
rect 1581 12257 1593 12291
rect 1627 12288 1639 12291
rect 1670 12288 1676 12300
rect 1627 12260 1676 12288
rect 1627 12257 1639 12260
rect 1581 12251 1639 12257
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2222 12288 2228 12300
rect 2179 12260 2228 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 3234 12288 3240 12300
rect 2915 12260 3240 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 3234 12248 3240 12260
rect 3292 12248 3298 12300
rect 4321 12291 4379 12297
rect 4321 12288 4333 12291
rect 3804 12260 4333 12288
rect 1486 12180 1492 12232
rect 1544 12220 1550 12232
rect 1762 12220 1768 12232
rect 1544 12192 1768 12220
rect 1544 12180 1550 12192
rect 1762 12180 1768 12192
rect 1820 12220 1826 12232
rect 2317 12223 2375 12229
rect 2317 12220 2329 12223
rect 1820 12192 2329 12220
rect 1820 12180 1826 12192
rect 2317 12189 2329 12192
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 3804 12096 3832 12260
rect 4321 12257 4333 12260
rect 4367 12257 4379 12291
rect 4321 12251 4379 12257
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 5442 12288 5448 12300
rect 4764 12260 5448 12288
rect 4764 12248 4770 12260
rect 5442 12248 5448 12260
rect 5500 12288 5506 12300
rect 6178 12297 6184 12300
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5500 12260 5917 12288
rect 5500 12248 5506 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 6172 12288 6184 12297
rect 6139 12260 6184 12288
rect 5905 12251 5963 12257
rect 6172 12251 6184 12260
rect 6178 12248 6184 12251
rect 6236 12248 6242 12300
rect 7558 12248 7564 12300
rect 7616 12248 7622 12300
rect 7742 12288 7748 12300
rect 7703 12260 7748 12288
rect 7742 12248 7748 12260
rect 7800 12288 7806 12300
rect 8202 12288 8208 12300
rect 7800 12260 8208 12288
rect 7800 12248 7806 12260
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 8570 12288 8576 12300
rect 8483 12260 8576 12288
rect 8570 12248 8576 12260
rect 8628 12288 8634 12300
rect 9490 12288 9496 12300
rect 8628 12260 9496 12288
rect 8628 12248 8634 12260
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 10597 12291 10655 12297
rect 10597 12288 10609 12291
rect 10192 12260 10609 12288
rect 10192 12248 10198 12260
rect 10597 12257 10609 12260
rect 10643 12257 10655 12291
rect 10597 12251 10655 12257
rect 11609 12291 11667 12297
rect 11609 12257 11621 12291
rect 11655 12288 11667 12291
rect 11698 12288 11704 12300
rect 11655 12260 11704 12288
rect 11655 12257 11667 12260
rect 11609 12251 11667 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11876 12291 11934 12297
rect 11876 12257 11888 12291
rect 11922 12288 11934 12291
rect 12250 12288 12256 12300
rect 11922 12260 12256 12288
rect 11922 12257 11934 12260
rect 11876 12251 11934 12257
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 12434 12248 12440 12300
rect 12492 12288 12498 12300
rect 12802 12288 12808 12300
rect 12492 12260 12808 12288
rect 12492 12248 12498 12260
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 14093 12291 14151 12297
rect 14093 12288 14105 12291
rect 13556 12260 14105 12288
rect 4062 12220 4068 12232
rect 4023 12192 4068 12220
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 7576 12220 7604 12248
rect 7834 12220 7840 12232
rect 7576 12192 7840 12220
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 8662 12220 8668 12232
rect 8623 12192 8668 12220
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 8846 12220 8852 12232
rect 8807 12192 8852 12220
rect 8846 12180 8852 12192
rect 8904 12220 8910 12232
rect 9582 12220 9588 12232
rect 8904 12192 9588 12220
rect 8904 12180 8910 12192
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 10689 12223 10747 12229
rect 10689 12220 10701 12223
rect 10100 12192 10701 12220
rect 10100 12180 10106 12192
rect 10689 12189 10701 12192
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 11054 12220 11060 12232
rect 10919 12192 11060 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 5445 12155 5503 12161
rect 5445 12121 5457 12155
rect 5491 12152 5503 12155
rect 5552 12152 5580 12180
rect 5718 12152 5724 12164
rect 5491 12124 5724 12152
rect 5491 12121 5503 12124
rect 5445 12115 5503 12121
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 8205 12155 8263 12161
rect 8205 12152 8217 12155
rect 6840 12124 8217 12152
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 3786 12084 3792 12096
rect 3559 12056 3792 12084
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 5537 12087 5595 12093
rect 5537 12053 5549 12087
rect 5583 12084 5595 12087
rect 6840 12084 6868 12124
rect 8205 12121 8217 12124
rect 8251 12121 8263 12155
rect 10704 12152 10732 12183
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 12894 12220 12900 12232
rect 12768 12192 12900 12220
rect 12768 12180 12774 12192
rect 12894 12180 12900 12192
rect 12952 12180 12958 12232
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 13556 12229 13584 12260
rect 14093 12257 14105 12260
rect 14139 12257 14151 12291
rect 14093 12251 14151 12257
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 14550 12288 14556 12300
rect 14424 12260 14556 12288
rect 14424 12248 14430 12260
rect 14550 12248 14556 12260
rect 14608 12288 14614 12300
rect 14921 12291 14979 12297
rect 14921 12288 14933 12291
rect 14608 12260 14933 12288
rect 14608 12248 14614 12260
rect 14921 12257 14933 12260
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12288 15531 12291
rect 15562 12288 15568 12300
rect 15519 12260 15568 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 15740 12291 15798 12297
rect 15740 12257 15752 12291
rect 15786 12288 15798 12291
rect 16298 12288 16304 12300
rect 15786 12260 16304 12288
rect 15786 12257 15798 12260
rect 15740 12251 15798 12257
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 17678 12248 17684 12300
rect 17736 12288 17742 12300
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 17736 12260 17877 12288
rect 17736 12248 17742 12260
rect 17865 12257 17877 12260
rect 17911 12257 17923 12291
rect 18598 12288 18604 12300
rect 17865 12251 17923 12257
rect 18156 12260 18604 12288
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 13504 12192 13553 12220
rect 13504 12180 13510 12192
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 15010 12220 15016 12232
rect 14323 12192 15016 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 15010 12180 15016 12192
rect 15068 12220 15074 12232
rect 15194 12220 15200 12232
rect 15068 12192 15200 12220
rect 15068 12180 15074 12192
rect 15194 12180 15200 12192
rect 15252 12180 15258 12232
rect 17770 12180 17776 12232
rect 17828 12220 17834 12232
rect 18156 12229 18184 12260
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 19420 12291 19478 12297
rect 19420 12257 19432 12291
rect 19466 12288 19478 12291
rect 19794 12288 19800 12300
rect 19466 12260 19800 12288
rect 19466 12257 19478 12260
rect 19420 12251 19478 12257
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 17957 12223 18015 12229
rect 17957 12220 17969 12223
rect 17828 12192 17969 12220
rect 17828 12180 17834 12192
rect 17957 12189 17969 12192
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12189 18199 12223
rect 18506 12220 18512 12232
rect 18467 12192 18512 12220
rect 18141 12183 18199 12189
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 19153 12223 19211 12229
rect 19153 12189 19165 12223
rect 19199 12189 19211 12223
rect 19153 12183 19211 12189
rect 11241 12155 11299 12161
rect 11241 12152 11253 12155
rect 10704 12124 11253 12152
rect 8205 12115 8263 12121
rect 11241 12121 11253 12124
rect 11287 12121 11299 12155
rect 11241 12115 11299 12121
rect 16666 12112 16672 12164
rect 16724 12152 16730 12164
rect 16942 12152 16948 12164
rect 16724 12124 16948 12152
rect 16724 12112 16730 12124
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 17586 12112 17592 12164
rect 17644 12152 17650 12164
rect 18969 12155 19027 12161
rect 18969 12152 18981 12155
rect 17644 12124 18981 12152
rect 17644 12112 17650 12124
rect 18969 12121 18981 12124
rect 19015 12121 19027 12155
rect 18969 12115 19027 12121
rect 5583 12056 6868 12084
rect 7285 12087 7343 12093
rect 5583 12053 5595 12056
rect 5537 12047 5595 12053
rect 7285 12053 7297 12087
rect 7331 12084 7343 12087
rect 7374 12084 7380 12096
rect 7331 12056 7380 12084
rect 7331 12053 7343 12056
rect 7285 12047 7343 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7561 12087 7619 12093
rect 7561 12084 7573 12087
rect 7524 12056 7573 12084
rect 7524 12044 7530 12056
rect 7561 12053 7573 12056
rect 7607 12053 7619 12087
rect 7561 12047 7619 12053
rect 7650 12044 7656 12096
rect 7708 12084 7714 12096
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7708 12056 8033 12084
rect 7708 12044 7714 12056
rect 8021 12053 8033 12056
rect 8067 12053 8079 12087
rect 8021 12047 8079 12053
rect 8938 12044 8944 12096
rect 8996 12084 9002 12096
rect 9861 12087 9919 12093
rect 9861 12084 9873 12087
rect 8996 12056 9873 12084
rect 8996 12044 9002 12056
rect 9861 12053 9873 12056
rect 9907 12053 9919 12087
rect 9861 12047 9919 12053
rect 10229 12087 10287 12093
rect 10229 12053 10241 12087
rect 10275 12084 10287 12087
rect 11790 12084 11796 12096
rect 10275 12056 11796 12084
rect 10275 12053 10287 12056
rect 10229 12047 10287 12053
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 12989 12087 13047 12093
rect 12989 12084 13001 12087
rect 12768 12056 13001 12084
rect 12768 12044 12774 12056
rect 12989 12053 13001 12056
rect 13035 12053 13047 12087
rect 12989 12047 13047 12053
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 14737 12087 14795 12093
rect 14737 12084 14749 12087
rect 13504 12056 14749 12084
rect 13504 12044 13510 12056
rect 14737 12053 14749 12056
rect 14783 12084 14795 12087
rect 16206 12084 16212 12096
rect 14783 12056 16212 12084
rect 14783 12053 14795 12056
rect 14737 12047 14795 12053
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 17405 12087 17463 12093
rect 17405 12053 17417 12087
rect 17451 12084 17463 12087
rect 17678 12084 17684 12096
rect 17451 12056 17684 12084
rect 17451 12053 17463 12056
rect 17405 12047 17463 12053
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 19168 12084 19196 12183
rect 20438 12084 20444 12096
rect 19168 12056 20444 12084
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 4890 11840 4896 11892
rect 4948 11880 4954 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 4948 11852 6377 11880
rect 4948 11840 4954 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6549 11883 6607 11889
rect 6549 11849 6561 11883
rect 6595 11880 6607 11883
rect 6822 11880 6828 11892
rect 6595 11852 6828 11880
rect 6595 11849 6607 11852
rect 6549 11843 6607 11849
rect 3786 11772 3792 11824
rect 3844 11812 3850 11824
rect 4157 11815 4215 11821
rect 4157 11812 4169 11815
rect 3844 11784 4169 11812
rect 3844 11772 3850 11784
rect 4157 11781 4169 11784
rect 4203 11812 4215 11815
rect 6564 11812 6592 11843
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 9217 11883 9275 11889
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 9674 11880 9680 11892
rect 9263 11852 9680 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 10134 11880 10140 11892
rect 10095 11852 10140 11880
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 11698 11840 11704 11892
rect 11756 11880 11762 11892
rect 12069 11883 12127 11889
rect 12069 11880 12081 11883
rect 11756 11852 12081 11880
rect 11756 11840 11762 11852
rect 12069 11849 12081 11852
rect 12115 11849 12127 11883
rect 12069 11843 12127 11849
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 12437 11883 12495 11889
rect 12437 11880 12449 11883
rect 12216 11852 12449 11880
rect 12216 11840 12222 11852
rect 12437 11849 12449 11852
rect 12483 11849 12495 11883
rect 13446 11880 13452 11892
rect 12437 11843 12495 11849
rect 12544 11852 13452 11880
rect 9490 11812 9496 11824
rect 4203 11784 5028 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 5000 11753 5028 11784
rect 5920 11784 6592 11812
rect 9451 11784 9496 11812
rect 5920 11753 5948 11784
rect 9490 11772 9496 11784
rect 9548 11772 9554 11824
rect 11882 11812 11888 11824
rect 11843 11784 11888 11812
rect 11882 11772 11888 11784
rect 11940 11772 11946 11824
rect 12544 11812 12572 11852
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 19426 11880 19432 11892
rect 14752 11852 19012 11880
rect 19387 11852 19432 11880
rect 12268 11784 12572 11812
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 6089 11747 6147 11753
rect 6089 11713 6101 11747
rect 6135 11744 6147 11747
rect 6362 11744 6368 11756
rect 6135 11716 6368 11744
rect 6135 11713 6147 11716
rect 6089 11707 6147 11713
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11676 2007 11679
rect 2498 11676 2504 11688
rect 1995 11648 2504 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 2866 11676 2872 11688
rect 2823 11648 2872 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 2866 11636 2872 11648
rect 2924 11676 2930 11688
rect 4154 11676 4160 11688
rect 2924 11648 4160 11676
rect 2924 11636 2930 11648
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 5258 11636 5264 11688
rect 5316 11676 5322 11688
rect 5534 11676 5540 11688
rect 5316 11648 5540 11676
rect 5316 11636 5322 11648
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 5718 11636 5724 11688
rect 5776 11676 5782 11688
rect 6104 11676 6132 11707
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 7374 11744 7380 11756
rect 6512 11716 7380 11744
rect 6512 11704 6518 11716
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 7834 11744 7840 11756
rect 7791 11716 7840 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 5776 11648 6132 11676
rect 5776 11636 5782 11648
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 7064 11648 7297 11676
rect 7064 11636 7070 11648
rect 7285 11645 7297 11648
rect 7331 11676 7343 11679
rect 7650 11676 7656 11688
rect 7331 11648 7656 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 10042 11676 10048 11688
rect 8036 11648 10048 11676
rect 3050 11617 3056 11620
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11577 2283 11611
rect 3044 11608 3056 11617
rect 3011 11580 3056 11608
rect 2225 11571 2283 11577
rect 3044 11571 3056 11580
rect 1670 11540 1676 11552
rect 1631 11512 1676 11540
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 2240 11540 2268 11571
rect 3050 11568 3056 11571
rect 3108 11568 3114 11620
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 8036 11608 8064 11648
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 10496 11679 10554 11685
rect 10496 11645 10508 11679
rect 10542 11676 10554 11679
rect 11054 11676 11060 11688
rect 10542 11648 11060 11676
rect 10542 11645 10554 11648
rect 10496 11639 10554 11645
rect 4120 11580 8064 11608
rect 8104 11611 8162 11617
rect 4120 11568 4126 11580
rect 8104 11577 8116 11611
rect 8150 11608 8162 11611
rect 8938 11608 8944 11620
rect 8150 11580 8944 11608
rect 8150 11577 8162 11580
rect 8104 11571 8162 11577
rect 8938 11568 8944 11580
rect 8996 11568 9002 11620
rect 10244 11608 10272 11639
rect 11054 11636 11060 11648
rect 11112 11676 11118 11688
rect 12268 11685 12296 11784
rect 12710 11772 12716 11824
rect 12768 11812 12774 11824
rect 12768 11784 13124 11812
rect 12768 11772 12774 11784
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12544 11716 13001 11744
rect 12253 11679 12311 11685
rect 11112 11648 11928 11676
rect 11112 11636 11118 11648
rect 10060 11580 10272 11608
rect 10060 11552 10088 11580
rect 11900 11552 11928 11648
rect 12253 11645 12265 11679
rect 12299 11645 12311 11679
rect 12544 11676 12572 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 13096 11744 13124 11784
rect 13262 11772 13268 11824
rect 13320 11812 13326 11824
rect 14090 11812 14096 11824
rect 13320 11784 14096 11812
rect 13320 11772 13326 11784
rect 14090 11772 14096 11784
rect 14148 11812 14154 11824
rect 14752 11812 14780 11852
rect 16298 11812 16304 11824
rect 14148 11784 14780 11812
rect 16211 11784 16304 11812
rect 14148 11772 14154 11784
rect 16298 11772 16304 11784
rect 16356 11812 16362 11824
rect 17586 11812 17592 11824
rect 16356 11784 16804 11812
rect 16356 11772 16362 11784
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13096 11716 13829 11744
rect 12989 11707 13047 11713
rect 13817 11713 13829 11716
rect 13863 11713 13875 11747
rect 16776 11744 16804 11784
rect 17144 11784 17592 11812
rect 17144 11753 17172 11784
rect 17586 11772 17592 11784
rect 17644 11772 17650 11824
rect 17770 11812 17776 11824
rect 17731 11784 17776 11812
rect 17770 11772 17776 11784
rect 17828 11772 17834 11824
rect 18984 11812 19012 11852
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 20809 11815 20867 11821
rect 20809 11812 20821 11815
rect 18984 11784 20821 11812
rect 20809 11781 20821 11784
rect 20855 11781 20867 11815
rect 20809 11775 20867 11781
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 13817 11707 13875 11713
rect 14108 11716 15056 11744
rect 16776 11716 17141 11744
rect 12802 11676 12808 11688
rect 12253 11639 12311 11645
rect 12452 11648 12572 11676
rect 12715 11648 12808 11676
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12452 11608 12480 11648
rect 12802 11636 12808 11648
rect 12860 11676 12866 11688
rect 13262 11676 13268 11688
rect 12860 11648 13268 11676
rect 12860 11636 12866 11648
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 14108 11685 14136 11716
rect 14093 11679 14151 11685
rect 14093 11676 14105 11679
rect 13504 11648 14105 11676
rect 13504 11636 13510 11648
rect 14093 11645 14105 11648
rect 14139 11645 14151 11679
rect 14093 11639 14151 11645
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 15028 11676 15056 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17236 11716 18184 11744
rect 17236 11676 17264 11716
rect 18046 11676 18052 11688
rect 15028 11648 17264 11676
rect 18007 11648 18052 11676
rect 14921 11639 14979 11645
rect 12216 11580 12480 11608
rect 12216 11568 12222 11580
rect 12526 11568 12532 11620
rect 12584 11608 12590 11620
rect 13630 11608 13636 11620
rect 12584 11580 13308 11608
rect 13591 11580 13636 11608
rect 12584 11568 12590 11580
rect 3234 11540 3240 11552
rect 2240 11512 3240 11540
rect 3234 11500 3240 11512
rect 3292 11540 3298 11552
rect 3694 11540 3700 11552
rect 3292 11512 3700 11540
rect 3292 11500 3298 11512
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 4430 11540 4436 11552
rect 4391 11512 4436 11540
rect 4430 11500 4436 11512
rect 4488 11500 4494 11552
rect 4798 11540 4804 11552
rect 4759 11512 4804 11540
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 4948 11512 4993 11540
rect 4948 11500 4954 11512
rect 5258 11500 5264 11552
rect 5316 11540 5322 11552
rect 5445 11543 5503 11549
rect 5445 11540 5457 11543
rect 5316 11512 5457 11540
rect 5316 11500 5322 11512
rect 5445 11509 5457 11512
rect 5491 11509 5503 11543
rect 5445 11503 5503 11509
rect 5813 11543 5871 11549
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 6270 11540 6276 11552
rect 5859 11512 6276 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6365 11543 6423 11549
rect 6365 11509 6377 11543
rect 6411 11540 6423 11543
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6411 11512 6837 11540
rect 6411 11509 6423 11512
rect 6365 11503 6423 11509
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 7190 11540 7196 11552
rect 7151 11512 7196 11540
rect 6825 11503 6883 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7708 11512 7757 11540
rect 7708 11500 7714 11512
rect 7745 11509 7757 11512
rect 7791 11540 7803 11543
rect 10042 11540 10048 11552
rect 7791 11512 10048 11540
rect 7791 11509 7803 11512
rect 7745 11503 7803 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 11609 11543 11667 11549
rect 11609 11540 11621 11543
rect 10744 11512 11621 11540
rect 10744 11500 10750 11512
rect 11609 11509 11621 11512
rect 11655 11509 11667 11543
rect 11882 11540 11888 11552
rect 11795 11512 11888 11540
rect 11609 11503 11667 11509
rect 11882 11500 11888 11512
rect 11940 11540 11946 11552
rect 12710 11540 12716 11552
rect 11940 11512 12716 11540
rect 11940 11500 11946 11512
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13280 11549 13308 11580
rect 13630 11568 13636 11580
rect 13688 11568 13694 11620
rect 13722 11568 13728 11620
rect 13780 11608 13786 11620
rect 13780 11580 13825 11608
rect 13780 11568 13786 11580
rect 14182 11568 14188 11620
rect 14240 11608 14246 11620
rect 14366 11608 14372 11620
rect 14240 11580 14372 11608
rect 14240 11568 14246 11580
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 13265 11543 13323 11549
rect 13265 11509 13277 11543
rect 13311 11509 13323 11543
rect 14936 11540 14964 11639
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18156 11676 18184 11716
rect 20441 11679 20499 11685
rect 20441 11676 20453 11679
rect 18156 11648 20453 11676
rect 20441 11645 20453 11648
rect 20487 11645 20499 11679
rect 20441 11639 20499 11645
rect 15188 11611 15246 11617
rect 15188 11577 15200 11611
rect 15234 11608 15246 11611
rect 15470 11608 15476 11620
rect 15234 11580 15476 11608
rect 15234 11577 15246 11580
rect 15188 11571 15246 11577
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 15654 11568 15660 11620
rect 15712 11608 15718 11620
rect 15712 11580 17080 11608
rect 15712 11568 15718 11580
rect 15562 11540 15568 11552
rect 14936 11512 15568 11540
rect 13265 11503 13323 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 16577 11543 16635 11549
rect 16577 11509 16589 11543
rect 16623 11540 16635 11543
rect 16666 11540 16672 11552
rect 16623 11512 16672 11540
rect 16623 11509 16635 11512
rect 16577 11503 16635 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 16942 11540 16948 11552
rect 16903 11512 16948 11540
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17052 11549 17080 11580
rect 18138 11568 18144 11620
rect 18196 11608 18202 11620
rect 18316 11611 18374 11617
rect 18316 11608 18328 11611
rect 18196 11580 18328 11608
rect 18196 11568 18202 11580
rect 18316 11577 18328 11580
rect 18362 11608 18374 11611
rect 18598 11608 18604 11620
rect 18362 11580 18604 11608
rect 18362 11577 18374 11580
rect 18316 11571 18374 11577
rect 18598 11568 18604 11580
rect 18656 11608 18662 11620
rect 19242 11608 19248 11620
rect 18656 11580 19248 11608
rect 18656 11568 18662 11580
rect 19242 11568 19248 11580
rect 19300 11608 19306 11620
rect 20073 11611 20131 11617
rect 20073 11608 20085 11611
rect 19300 11580 20085 11608
rect 19300 11568 19306 11580
rect 20073 11577 20085 11580
rect 20119 11577 20131 11611
rect 20073 11571 20131 11577
rect 17037 11543 17095 11549
rect 17037 11509 17049 11543
rect 17083 11540 17095 11543
rect 19610 11540 19616 11552
rect 17083 11512 19616 11540
rect 17083 11509 17095 11512
rect 17037 11503 17095 11509
rect 19610 11500 19616 11512
rect 19668 11500 19674 11552
rect 19794 11540 19800 11552
rect 19755 11512 19800 11540
rect 19794 11500 19800 11512
rect 19852 11500 19858 11552
rect 20438 11500 20444 11552
rect 20496 11540 20502 11552
rect 21177 11543 21235 11549
rect 21177 11540 21189 11543
rect 20496 11512 21189 11540
rect 20496 11500 20502 11512
rect 21177 11509 21189 11512
rect 21223 11509 21235 11543
rect 21177 11503 21235 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2498 11296 2504 11348
rect 2556 11296 2562 11348
rect 2682 11336 2688 11348
rect 2643 11308 2688 11336
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 4249 11339 4307 11345
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 4522 11336 4528 11348
rect 4295 11308 4528 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 5166 11336 5172 11348
rect 4663 11308 5172 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 5166 11296 5172 11308
rect 5224 11336 5230 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 5224 11308 5273 11336
rect 5224 11296 5230 11308
rect 5261 11305 5273 11308
rect 5307 11305 5319 11339
rect 5261 11299 5319 11305
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 5500 11308 5733 11336
rect 5500 11296 5506 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 5721 11299 5779 11305
rect 6365 11339 6423 11345
rect 6365 11305 6377 11339
rect 6411 11336 6423 11339
rect 7190 11336 7196 11348
rect 6411 11308 7196 11336
rect 6411 11305 6423 11308
rect 6365 11299 6423 11305
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 7377 11339 7435 11345
rect 7377 11305 7389 11339
rect 7423 11336 7435 11339
rect 8938 11336 8944 11348
rect 7423 11308 8944 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9309 11339 9367 11345
rect 9309 11305 9321 11339
rect 9355 11336 9367 11339
rect 9398 11336 9404 11348
rect 9355 11308 9404 11336
rect 9355 11305 9367 11308
rect 9309 11299 9367 11305
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10192 11308 10517 11336
rect 10192 11296 10198 11308
rect 10505 11305 10517 11308
rect 10551 11305 10563 11339
rect 10505 11299 10563 11305
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11517 11339 11575 11345
rect 11517 11336 11529 11339
rect 10928 11308 11529 11336
rect 10928 11296 10934 11308
rect 11517 11305 11529 11308
rect 11563 11305 11575 11339
rect 11517 11299 11575 11305
rect 11977 11339 12035 11345
rect 11977 11305 11989 11339
rect 12023 11336 12035 11339
rect 13446 11336 13452 11348
rect 12023 11308 13452 11336
rect 12023 11305 12035 11308
rect 11977 11299 12035 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13633 11339 13691 11345
rect 13633 11305 13645 11339
rect 13679 11336 13691 11339
rect 13814 11336 13820 11348
rect 13679 11308 13820 11336
rect 13679 11305 13691 11308
rect 13633 11299 13691 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 14185 11339 14243 11345
rect 14185 11305 14197 11339
rect 14231 11305 14243 11339
rect 14185 11299 14243 11305
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15654 11336 15660 11348
rect 15335 11308 15660 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 1670 11228 1676 11280
rect 1728 11268 1734 11280
rect 2041 11271 2099 11277
rect 2041 11268 2053 11271
rect 1728 11240 2053 11268
rect 1728 11228 1734 11240
rect 2041 11237 2053 11240
rect 2087 11237 2099 11271
rect 2516 11268 2544 11296
rect 6457 11271 6515 11277
rect 6457 11268 6469 11271
rect 2516 11240 6469 11268
rect 2041 11231 2099 11237
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11200 1823 11203
rect 1946 11200 1952 11212
rect 1811 11172 1952 11200
rect 1811 11169 1823 11172
rect 1765 11163 1823 11169
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 2498 11200 2504 11212
rect 2459 11172 2504 11200
rect 2498 11160 2504 11172
rect 2556 11160 2562 11212
rect 2038 11092 2044 11144
rect 2096 11132 2102 11144
rect 2222 11132 2228 11144
rect 2096 11104 2228 11132
rect 2096 11092 2102 11104
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2608 11132 2636 11240
rect 6457 11237 6469 11240
rect 6503 11237 6515 11271
rect 6457 11231 6515 11237
rect 6840 11240 8340 11268
rect 4706 11200 4712 11212
rect 4667 11172 4712 11200
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11200 5963 11203
rect 5994 11200 6000 11212
rect 5951 11172 6000 11200
rect 5951 11169 5963 11172
rect 5905 11163 5963 11169
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6270 11200 6276 11212
rect 6231 11172 6276 11200
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 6840 11200 6868 11240
rect 6564 11172 6868 11200
rect 6917 11203 6975 11209
rect 2682 11132 2688 11144
rect 2608 11104 2688 11132
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 3050 11092 3056 11144
rect 3108 11132 3114 11144
rect 3145 11135 3203 11141
rect 3145 11132 3157 11135
rect 3108 11104 3157 11132
rect 3108 11092 3114 11104
rect 3145 11101 3157 11104
rect 3191 11132 3203 11135
rect 3513 11135 3571 11141
rect 3513 11132 3525 11135
rect 3191 11104 3525 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3513 11101 3525 11104
rect 3559 11132 3571 11135
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 3559 11104 4905 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 4893 11101 4905 11104
rect 4939 11132 4951 11135
rect 6454 11132 6460 11144
rect 4939 11104 6460 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 6564 11064 6592 11172
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 7282 11200 7288 11212
rect 6963 11172 7288 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 7650 11200 7656 11212
rect 7607 11172 7656 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 7006 11132 7012 11144
rect 6967 11104 7012 11132
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11132 7251 11135
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7239 11104 7389 11132
rect 7239 11101 7251 11104
rect 7193 11095 7251 11101
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 4120 11036 6592 11064
rect 4120 11024 4126 11036
rect 6638 11024 6644 11076
rect 6696 11064 6702 11076
rect 7208 11064 7236 11095
rect 6696 11036 7236 11064
rect 6696 11024 6702 11036
rect 1673 10999 1731 11005
rect 1673 10965 1685 10999
rect 1719 10996 1731 10999
rect 2222 10996 2228 11008
rect 1719 10968 2228 10996
rect 1719 10965 1731 10968
rect 1673 10959 1731 10965
rect 2222 10956 2228 10968
rect 2280 10956 2286 11008
rect 2498 10956 2504 11008
rect 2556 10996 2562 11008
rect 2866 10996 2872 11008
rect 2556 10968 2872 10996
rect 2556 10956 2562 10968
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 3881 10999 3939 11005
rect 3881 10965 3893 10999
rect 3927 10996 3939 10999
rect 3970 10996 3976 11008
rect 3927 10968 3976 10996
rect 3927 10965 3939 10968
rect 3881 10959 3939 10965
rect 3970 10956 3976 10968
rect 4028 10996 4034 11008
rect 6365 10999 6423 11005
rect 6365 10996 6377 10999
rect 4028 10968 6377 10996
rect 4028 10956 4034 10968
rect 6365 10965 6377 10968
rect 6411 10965 6423 10999
rect 6365 10959 6423 10965
rect 6457 10999 6515 11005
rect 6457 10965 6469 10999
rect 6503 10996 6515 10999
rect 6549 10999 6607 11005
rect 6549 10996 6561 10999
rect 6503 10968 6561 10996
rect 6503 10965 6515 10968
rect 6457 10959 6515 10965
rect 6549 10965 6561 10968
rect 6595 10965 6607 10999
rect 6549 10959 6607 10965
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7576 10996 7604 11163
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 7828 11203 7886 11209
rect 7828 11169 7840 11203
rect 7874 11200 7886 11203
rect 8202 11200 8208 11212
rect 7874 11172 8208 11200
rect 7874 11169 7886 11172
rect 7828 11163 7886 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 8312 11200 8340 11240
rect 8846 11228 8852 11280
rect 8904 11268 8910 11280
rect 10229 11271 10287 11277
rect 10229 11268 10241 11271
rect 8904 11240 10241 11268
rect 8904 11228 8910 11240
rect 10229 11237 10241 11240
rect 10275 11237 10287 11271
rect 10229 11231 10287 11237
rect 11790 11228 11796 11280
rect 11848 11268 11854 11280
rect 12345 11271 12403 11277
rect 12345 11268 12357 11271
rect 11848 11240 12357 11268
rect 11848 11228 11854 11240
rect 12345 11237 12357 11240
rect 12391 11237 12403 11271
rect 12345 11231 12403 11237
rect 12437 11271 12495 11277
rect 12437 11237 12449 11271
rect 12483 11268 12495 11271
rect 12526 11268 12532 11280
rect 12483 11240 12532 11268
rect 12483 11237 12495 11240
rect 12437 11231 12495 11237
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 13906 11268 13912 11280
rect 12952 11240 13912 11268
rect 12952 11228 12958 11240
rect 13906 11228 13912 11240
rect 13964 11228 13970 11280
rect 14200 11268 14228 11299
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16301 11339 16359 11345
rect 16301 11305 16313 11339
rect 16347 11336 16359 11339
rect 16942 11336 16948 11348
rect 16347 11308 16948 11336
rect 16347 11305 16359 11308
rect 16301 11299 16359 11305
rect 16942 11296 16948 11308
rect 17000 11336 17006 11348
rect 17221 11339 17279 11345
rect 17221 11336 17233 11339
rect 17000 11308 17233 11336
rect 17000 11296 17006 11308
rect 17221 11305 17233 11308
rect 17267 11305 17279 11339
rect 17221 11299 17279 11305
rect 17497 11339 17555 11345
rect 17497 11305 17509 11339
rect 17543 11336 17555 11339
rect 17954 11336 17960 11348
rect 17543 11308 17960 11336
rect 17543 11305 17555 11308
rect 17497 11299 17555 11305
rect 17954 11296 17960 11308
rect 18012 11296 18018 11348
rect 18969 11339 19027 11345
rect 18969 11305 18981 11339
rect 19015 11336 19027 11339
rect 19426 11336 19432 11348
rect 19015 11308 19432 11336
rect 19015 11305 19027 11308
rect 18969 11299 19027 11305
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 19610 11336 19616 11348
rect 19571 11308 19616 11336
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 20438 11336 20444 11348
rect 20399 11308 20444 11336
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 15378 11268 15384 11280
rect 14200 11240 15384 11268
rect 15378 11228 15384 11240
rect 15436 11228 15442 11280
rect 17865 11271 17923 11277
rect 17865 11237 17877 11271
rect 17911 11268 17923 11271
rect 18506 11268 18512 11280
rect 17911 11240 18512 11268
rect 17911 11237 17923 11240
rect 17865 11231 17923 11237
rect 18506 11228 18512 11240
rect 18564 11228 18570 11280
rect 19242 11268 19248 11280
rect 19203 11240 19248 11268
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 11054 11200 11060 11212
rect 8312 11172 11060 11200
rect 11054 11160 11060 11172
rect 11112 11200 11118 11212
rect 11149 11203 11207 11209
rect 11149 11200 11161 11203
rect 11112 11172 11161 11200
rect 11112 11160 11118 11172
rect 11149 11169 11161 11172
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 13081 11203 13139 11209
rect 13081 11169 13093 11203
rect 13127 11200 13139 11203
rect 13541 11203 13599 11209
rect 13541 11200 13553 11203
rect 13127 11172 13553 11200
rect 13127 11169 13139 11172
rect 13081 11163 13139 11169
rect 13541 11169 13553 11172
rect 13587 11169 13599 11203
rect 14550 11200 14556 11212
rect 14511 11172 14556 11200
rect 13541 11163 13599 11169
rect 10686 11092 10692 11144
rect 10744 11132 10750 11144
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 10744 11104 12541 11132
rect 10744 11092 10750 11104
rect 12529 11101 12541 11104
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 8570 11024 8576 11076
rect 8628 11064 8634 11076
rect 13096 11064 13124 11163
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 15010 11200 15016 11212
rect 14700 11172 15016 11200
rect 14700 11160 14706 11172
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 15654 11200 15660 11212
rect 15615 11172 15660 11200
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 16206 11160 16212 11212
rect 16264 11200 16270 11212
rect 16945 11203 17003 11209
rect 16945 11200 16957 11203
rect 16264 11172 16957 11200
rect 16264 11160 16270 11172
rect 16945 11169 16957 11172
rect 16991 11200 17003 11203
rect 17770 11200 17776 11212
rect 16991 11172 17776 11200
rect 16991 11169 17003 11172
rect 16945 11163 17003 11169
rect 17770 11160 17776 11172
rect 17828 11160 17834 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 17972 11172 18613 11200
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 14829 11135 14887 11141
rect 13780 11104 13825 11132
rect 13780 11092 13786 11104
rect 14829 11101 14841 11135
rect 14875 11132 14887 11135
rect 15102 11132 15108 11144
rect 14875 11104 15108 11132
rect 14875 11101 14887 11104
rect 14829 11095 14887 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15344 11104 15761 11132
rect 15344 11092 15350 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 8628 11036 13124 11064
rect 13173 11067 13231 11073
rect 8628 11024 8634 11036
rect 13173 11033 13185 11067
rect 13219 11064 13231 11067
rect 14642 11064 14648 11076
rect 13219 11036 14648 11064
rect 13219 11033 13231 11036
rect 13173 11027 13231 11033
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 15470 11024 15476 11076
rect 15528 11064 15534 11076
rect 15856 11064 15884 11095
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 17972 11141 18000 11172
rect 18601 11169 18613 11172
rect 18647 11169 18659 11203
rect 18601 11163 18659 11169
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 16724 11104 17969 11132
rect 16724 11092 16730 11104
rect 17957 11101 17969 11104
rect 18003 11101 18015 11135
rect 18138 11132 18144 11144
rect 18099 11104 18144 11132
rect 17957 11095 18015 11101
rect 18138 11092 18144 11104
rect 18196 11092 18202 11144
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 19392 11104 20576 11132
rect 19392 11092 19398 11104
rect 20548 11076 20576 11104
rect 15528 11036 15884 11064
rect 15528 11024 15534 11036
rect 16114 11024 16120 11076
rect 16172 11064 16178 11076
rect 18782 11064 18788 11076
rect 16172 11036 18788 11064
rect 16172 11024 16178 11036
rect 18782 11024 18788 11036
rect 18840 11064 18846 11076
rect 19981 11067 20039 11073
rect 19981 11064 19993 11067
rect 18840 11036 19993 11064
rect 18840 11024 18846 11036
rect 19981 11033 19993 11036
rect 20027 11033 20039 11067
rect 19981 11027 20039 11033
rect 20530 11024 20536 11076
rect 20588 11064 20594 11076
rect 21085 11067 21143 11073
rect 21085 11064 21097 11067
rect 20588 11036 21097 11064
rect 20588 11024 20594 11036
rect 21085 11033 21097 11036
rect 21131 11033 21143 11067
rect 21085 11027 21143 11033
rect 6972 10968 7604 10996
rect 6972 10956 6978 10968
rect 8202 10956 8208 11008
rect 8260 10996 8266 11008
rect 8938 10996 8944 11008
rect 8260 10968 8944 10996
rect 8260 10956 8266 10968
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 9858 10996 9864 11008
rect 9819 10968 9864 10996
rect 9858 10956 9864 10968
rect 9916 10956 9922 11008
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13078 10996 13084 11008
rect 12952 10968 13084 10996
rect 12952 10956 12958 10968
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 16390 10956 16396 11008
rect 16448 10996 16454 11008
rect 16761 10999 16819 11005
rect 16761 10996 16773 10999
rect 16448 10968 16773 10996
rect 16448 10956 16454 10968
rect 16761 10965 16773 10968
rect 16807 10996 16819 10999
rect 17954 10996 17960 11008
rect 16807 10968 17960 10996
rect 16807 10965 16819 10968
rect 16761 10959 16819 10965
rect 17954 10956 17960 10968
rect 18012 10956 18018 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 5166 10792 5172 10804
rect 4120 10764 4568 10792
rect 5127 10764 5172 10792
rect 4120 10752 4126 10764
rect 4433 10727 4491 10733
rect 4433 10724 4445 10727
rect 3896 10696 4445 10724
rect 3896 10668 3924 10696
rect 4433 10693 4445 10696
rect 4479 10693 4491 10727
rect 4540 10724 4568 10764
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 6086 10752 6092 10804
rect 6144 10792 6150 10804
rect 6181 10795 6239 10801
rect 6181 10792 6193 10795
rect 6144 10764 6193 10792
rect 6144 10752 6150 10764
rect 6181 10761 6193 10764
rect 6227 10761 6239 10795
rect 8570 10792 8576 10804
rect 6181 10755 6239 10761
rect 6288 10764 8576 10792
rect 6288 10724 6316 10764
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 9493 10795 9551 10801
rect 9493 10792 9505 10795
rect 8812 10764 9505 10792
rect 8812 10752 8818 10764
rect 9493 10761 9505 10764
rect 9539 10761 9551 10795
rect 9493 10755 9551 10761
rect 10781 10795 10839 10801
rect 10781 10761 10793 10795
rect 10827 10792 10839 10795
rect 12710 10792 12716 10804
rect 10827 10764 12716 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 15470 10792 15476 10804
rect 15431 10764 15476 10792
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 17954 10752 17960 10804
rect 18012 10792 18018 10804
rect 20530 10792 20536 10804
rect 18012 10764 19656 10792
rect 20491 10764 20536 10792
rect 18012 10752 18018 10764
rect 6638 10724 6644 10736
rect 4540 10696 6316 10724
rect 6599 10696 6644 10724
rect 4433 10687 4491 10693
rect 6638 10684 6644 10696
rect 6696 10684 6702 10736
rect 8202 10724 8208 10736
rect 8163 10696 8208 10724
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 8389 10727 8447 10733
rect 8389 10693 8401 10727
rect 8435 10724 8447 10727
rect 8481 10727 8539 10733
rect 8481 10724 8493 10727
rect 8435 10696 8493 10724
rect 8435 10693 8447 10696
rect 8389 10687 8447 10693
rect 8481 10693 8493 10696
rect 8527 10693 8539 10727
rect 8481 10687 8539 10693
rect 8938 10684 8944 10736
rect 8996 10724 9002 10736
rect 8996 10696 9076 10724
rect 8996 10684 9002 10696
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2498 10656 2504 10668
rect 1719 10628 2504 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 3234 10656 3240 10668
rect 2823 10628 3240 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 3878 10656 3884 10668
rect 3839 10628 3884 10656
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10656 4123 10659
rect 5718 10656 5724 10668
rect 4111 10628 5724 10656
rect 4111 10625 4123 10628
rect 4065 10619 4123 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 9048 10665 9076 10696
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 9079 10628 10057 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 10045 10625 10057 10628
rect 10091 10656 10103 10659
rect 10870 10656 10876 10668
rect 10091 10628 10876 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 11425 10659 11483 10665
rect 11425 10625 11437 10659
rect 11471 10656 11483 10659
rect 11974 10656 11980 10668
rect 11471 10628 11980 10656
rect 11471 10625 11483 10628
rect 11425 10619 11483 10625
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 14090 10656 14096 10668
rect 14051 10628 14096 10656
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 18064 10665 18092 10764
rect 19628 10736 19656 10764
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 19610 10684 19616 10736
rect 19668 10724 19674 10736
rect 19797 10727 19855 10733
rect 19797 10724 19809 10727
rect 19668 10696 19809 10724
rect 19668 10684 19674 10696
rect 19797 10693 19809 10696
rect 19843 10724 19855 10727
rect 20165 10727 20223 10733
rect 20165 10724 20177 10727
rect 19843 10696 20177 10724
rect 19843 10693 19855 10696
rect 19797 10687 19855 10693
rect 20165 10693 20177 10696
rect 20211 10724 20223 10727
rect 20438 10724 20444 10736
rect 20211 10696 20444 10724
rect 20211 10693 20223 10696
rect 20165 10687 20223 10693
rect 20438 10684 20444 10696
rect 20496 10684 20502 10736
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 1397 10591 1455 10597
rect 1397 10588 1409 10591
rect 1360 10560 1409 10588
rect 1360 10548 1366 10560
rect 1397 10557 1409 10560
rect 1443 10557 1455 10591
rect 1397 10551 1455 10557
rect 1486 10548 1492 10600
rect 1544 10588 1550 10600
rect 2314 10588 2320 10600
rect 1544 10560 2320 10588
rect 1544 10548 1550 10560
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 6840 10588 6868 10616
rect 8846 10588 8852 10600
rect 5592 10560 6868 10588
rect 6912 10560 8515 10588
rect 8807 10560 8852 10588
rect 5592 10548 5598 10560
rect 2501 10523 2559 10529
rect 2501 10489 2513 10523
rect 2547 10520 2559 10523
rect 3050 10520 3056 10532
rect 2547 10492 3056 10520
rect 2547 10489 2559 10492
rect 2501 10483 2559 10489
rect 3050 10480 3056 10492
rect 3108 10480 3114 10532
rect 4706 10480 4712 10532
rect 4764 10520 4770 10532
rect 4893 10523 4951 10529
rect 4893 10520 4905 10523
rect 4764 10492 4905 10520
rect 4764 10480 4770 10492
rect 4893 10489 4905 10492
rect 4939 10520 4951 10523
rect 6912 10520 6940 10560
rect 7098 10529 7104 10532
rect 7092 10520 7104 10529
rect 4939 10492 6940 10520
rect 7059 10492 7104 10520
rect 4939 10489 4951 10492
rect 4893 10483 4951 10489
rect 7092 10483 7104 10492
rect 7098 10480 7104 10483
rect 7156 10480 7162 10532
rect 8389 10523 8447 10529
rect 8389 10520 8401 10523
rect 7484 10492 8401 10520
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 2133 10455 2191 10461
rect 2133 10452 2145 10455
rect 2004 10424 2145 10452
rect 2004 10412 2010 10424
rect 2133 10421 2145 10424
rect 2179 10421 2191 10455
rect 2133 10415 2191 10421
rect 2314 10412 2320 10464
rect 2372 10452 2378 10464
rect 2593 10455 2651 10461
rect 2593 10452 2605 10455
rect 2372 10424 2605 10452
rect 2372 10412 2378 10424
rect 2593 10421 2605 10424
rect 2639 10421 2651 10455
rect 3234 10452 3240 10464
rect 3195 10424 3240 10452
rect 2593 10415 2651 10421
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 3326 10412 3332 10464
rect 3384 10452 3390 10464
rect 3421 10455 3479 10461
rect 3421 10452 3433 10455
rect 3384 10424 3433 10452
rect 3384 10412 3390 10424
rect 3421 10421 3433 10424
rect 3467 10421 3479 10455
rect 3421 10415 3479 10421
rect 3789 10455 3847 10461
rect 3789 10421 3801 10455
rect 3835 10452 3847 10455
rect 3970 10452 3976 10464
rect 3835 10424 3976 10452
rect 3835 10421 3847 10424
rect 3789 10415 3847 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10452 5687 10455
rect 5718 10452 5724 10464
rect 5675 10424 5724 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7484 10452 7512 10492
rect 8389 10489 8401 10492
rect 8435 10489 8447 10523
rect 8487 10520 8515 10560
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 8941 10591 8999 10597
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 9398 10588 9404 10600
rect 8987 10560 9404 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 11112 10560 11161 10588
rect 11112 10548 11118 10560
rect 11149 10557 11161 10560
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 11756 10560 12449 10588
rect 11756 10548 11762 10560
rect 12437 10557 12449 10560
rect 12483 10588 12495 10591
rect 13446 10588 13452 10600
rect 12483 10560 13452 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 15562 10548 15568 10600
rect 15620 10588 15626 10600
rect 15749 10591 15807 10597
rect 15749 10588 15761 10591
rect 15620 10560 15761 10588
rect 15620 10548 15626 10560
rect 15749 10557 15761 10560
rect 15795 10588 15807 10591
rect 16390 10588 16396 10600
rect 15795 10560 16396 10588
rect 15795 10557 15807 10560
rect 15749 10551 15807 10557
rect 16390 10548 16396 10560
rect 16448 10548 16454 10600
rect 18316 10591 18374 10597
rect 18316 10557 18328 10591
rect 18362 10588 18374 10591
rect 19426 10588 19432 10600
rect 18362 10560 19432 10588
rect 18362 10557 18374 10560
rect 18316 10551 18374 10557
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 9953 10523 10011 10529
rect 9953 10520 9965 10523
rect 8487 10492 9965 10520
rect 8389 10483 8447 10489
rect 9953 10489 9965 10492
rect 9999 10520 10011 10523
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 9999 10492 10517 10520
rect 9999 10489 10011 10492
rect 9953 10483 10011 10489
rect 10505 10489 10517 10492
rect 10551 10489 10563 10523
rect 10505 10483 10563 10489
rect 10778 10480 10784 10532
rect 10836 10520 10842 10532
rect 11241 10523 11299 10529
rect 11241 10520 11253 10523
rect 10836 10492 11253 10520
rect 10836 10480 10842 10492
rect 11241 10489 11253 10492
rect 11287 10520 11299 10523
rect 11514 10520 11520 10532
rect 11287 10492 11520 10520
rect 11287 10489 11299 10492
rect 11241 10483 11299 10489
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 12704 10523 12762 10529
rect 12704 10489 12716 10523
rect 12750 10520 12762 10523
rect 13078 10520 13084 10532
rect 12750 10492 13084 10520
rect 12750 10489 12762 10492
rect 12704 10483 12762 10489
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 14360 10523 14418 10529
rect 14360 10489 14372 10523
rect 14406 10520 14418 10523
rect 15102 10520 15108 10532
rect 14406 10492 15108 10520
rect 14406 10489 14418 10492
rect 14360 10483 14418 10489
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 16022 10529 16028 10532
rect 16016 10520 16028 10529
rect 15935 10492 16028 10520
rect 16016 10483 16028 10492
rect 16080 10520 16086 10532
rect 16080 10492 19472 10520
rect 16022 10480 16028 10483
rect 16080 10480 16086 10492
rect 9858 10452 9864 10464
rect 7064 10424 7512 10452
rect 9819 10424 9864 10452
rect 7064 10412 7070 10424
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 11885 10455 11943 10461
rect 11885 10421 11897 10455
rect 11931 10452 11943 10455
rect 12802 10452 12808 10464
rect 11931 10424 12808 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13780 10424 13829 10452
rect 13780 10412 13786 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 17126 10452 17132 10464
rect 17087 10424 17132 10452
rect 13817 10415 13875 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17402 10452 17408 10464
rect 17363 10424 17408 10452
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 19444 10461 19472 10492
rect 19429 10455 19487 10461
rect 19429 10421 19441 10455
rect 19475 10421 19487 10455
rect 19429 10415 19487 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2317 10251 2375 10257
rect 2317 10248 2329 10251
rect 2280 10220 2329 10248
rect 2280 10208 2286 10220
rect 2317 10217 2329 10220
rect 2363 10248 2375 10251
rect 2498 10248 2504 10260
rect 2363 10220 2504 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 6178 10208 6184 10260
rect 6236 10248 6242 10260
rect 8021 10251 8079 10257
rect 8021 10248 8033 10251
rect 6236 10220 8033 10248
rect 6236 10208 6242 10220
rect 8021 10217 8033 10220
rect 8067 10217 8079 10251
rect 8021 10211 8079 10217
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 10318 10248 10324 10260
rect 8527 10220 10324 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 13078 10248 13084 10260
rect 10428 10220 12940 10248
rect 13039 10220 13084 10248
rect 1762 10180 1768 10192
rect 1675 10152 1768 10180
rect 1762 10140 1768 10152
rect 1820 10180 1826 10192
rect 1820 10152 2544 10180
rect 1820 10140 1826 10152
rect 2222 10112 2228 10124
rect 2183 10084 2228 10112
rect 2222 10072 2228 10084
rect 2280 10072 2286 10124
rect 2516 10053 2544 10152
rect 2682 10140 2688 10192
rect 2740 10180 2746 10192
rect 2958 10180 2964 10192
rect 2740 10152 2964 10180
rect 2740 10140 2746 10152
rect 2958 10140 2964 10152
rect 3016 10180 3022 10192
rect 4332 10183 4390 10189
rect 3016 10152 4108 10180
rect 3016 10140 3022 10152
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 3510 10112 3516 10124
rect 3283 10084 3516 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 4080 10121 4108 10152
rect 4332 10149 4344 10183
rect 4378 10180 4390 10183
rect 5718 10180 5724 10192
rect 4378 10152 5724 10180
rect 4378 10149 4390 10152
rect 4332 10143 4390 10149
rect 5718 10140 5724 10152
rect 5776 10180 5782 10192
rect 10428 10180 10456 10220
rect 5776 10152 10456 10180
rect 12912 10180 12940 10220
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 13188 10220 17785 10248
rect 13188 10180 13216 10220
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 18141 10251 18199 10257
rect 18141 10217 18153 10251
rect 18187 10248 18199 10251
rect 18506 10248 18512 10260
rect 18187 10220 18512 10248
rect 18187 10217 18199 10220
rect 18141 10211 18199 10217
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 18782 10248 18788 10260
rect 18743 10220 18788 10248
rect 18782 10208 18788 10220
rect 18840 10208 18846 10260
rect 19245 10251 19303 10257
rect 19245 10217 19257 10251
rect 19291 10248 19303 10251
rect 19610 10248 19616 10260
rect 19291 10220 19616 10248
rect 19291 10217 19303 10220
rect 19245 10211 19303 10217
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 19978 10248 19984 10260
rect 19891 10220 19984 10248
rect 19978 10208 19984 10220
rect 20036 10248 20042 10260
rect 20530 10248 20536 10260
rect 20036 10220 20536 10248
rect 20036 10208 20042 10220
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 12912 10152 13216 10180
rect 13624 10183 13682 10189
rect 5776 10140 5782 10152
rect 13624 10149 13636 10183
rect 13670 10180 13682 10183
rect 13722 10180 13728 10192
rect 13670 10152 13728 10180
rect 13670 10149 13682 10152
rect 13624 10143 13682 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 15105 10183 15163 10189
rect 15105 10149 15117 10183
rect 15151 10180 15163 10183
rect 15286 10180 15292 10192
rect 15151 10152 15292 10180
rect 15151 10149 15163 10152
rect 15105 10143 15163 10149
rect 15286 10140 15292 10152
rect 15344 10140 15350 10192
rect 15838 10180 15844 10192
rect 15799 10152 15844 10180
rect 15838 10140 15844 10152
rect 15896 10140 15902 10192
rect 16660 10183 16718 10189
rect 16660 10149 16672 10183
rect 16706 10180 16718 10183
rect 17126 10180 17132 10192
rect 16706 10152 17132 10180
rect 16706 10149 16718 10152
rect 16660 10143 16718 10149
rect 17126 10140 17132 10152
rect 17184 10140 17190 10192
rect 5994 10121 6000 10124
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10081 4123 10115
rect 5988 10112 6000 10121
rect 5955 10084 6000 10112
rect 4065 10075 4123 10081
rect 5988 10075 6000 10084
rect 6052 10112 6058 10124
rect 6822 10112 6828 10124
rect 6052 10084 6828 10112
rect 5994 10072 6000 10075
rect 6052 10072 6058 10084
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7466 10112 7472 10124
rect 6972 10084 7472 10112
rect 6972 10072 6978 10084
rect 7466 10072 7472 10084
rect 7524 10112 7530 10124
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 7524 10084 7941 10112
rect 7524 10072 7530 10084
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 8754 10112 8760 10124
rect 8435 10084 8760 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 8754 10072 8760 10084
rect 8812 10072 8818 10124
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 9033 10115 9091 10121
rect 9033 10112 9045 10115
rect 8904 10084 9045 10112
rect 8904 10072 8910 10084
rect 9033 10081 9045 10084
rect 9079 10081 9091 10115
rect 10042 10112 10048 10124
rect 10003 10084 10048 10112
rect 9033 10075 9091 10081
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10312 10115 10370 10121
rect 10312 10081 10324 10115
rect 10358 10112 10370 10115
rect 10686 10112 10692 10124
rect 10358 10084 10692 10112
rect 10358 10081 10370 10084
rect 10312 10075 10370 10081
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 11698 10112 11704 10124
rect 11659 10084 11704 10112
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11974 10121 11980 10124
rect 11968 10112 11980 10121
rect 11935 10084 11980 10112
rect 11968 10075 11980 10084
rect 11974 10072 11980 10075
rect 12032 10072 12038 10124
rect 13357 10115 13415 10121
rect 13357 10081 13369 10115
rect 13403 10112 13415 10115
rect 13446 10112 13452 10124
rect 13403 10084 13452 10112
rect 13403 10081 13415 10084
rect 13357 10075 13415 10081
rect 13446 10072 13452 10084
rect 13504 10112 13510 10124
rect 14090 10112 14096 10124
rect 13504 10084 14096 10112
rect 13504 10072 13510 10084
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 15749 10115 15807 10121
rect 15749 10081 15761 10115
rect 15795 10112 15807 10115
rect 15930 10112 15936 10124
rect 15795 10084 15936 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 16390 10112 16396 10124
rect 16351 10084 16396 10112
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 18509 10115 18567 10121
rect 18509 10081 18521 10115
rect 18555 10112 18567 10115
rect 18598 10112 18604 10124
rect 18555 10084 18604 10112
rect 18555 10081 18567 10084
rect 18509 10075 18567 10081
rect 18598 10072 18604 10084
rect 18656 10072 18662 10124
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10044 2559 10047
rect 3326 10044 3332 10056
rect 2547 10016 3188 10044
rect 3287 10016 3332 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 1857 9979 1915 9985
rect 1857 9945 1869 9979
rect 1903 9976 1915 9979
rect 3050 9976 3056 9988
rect 1903 9948 3056 9976
rect 1903 9945 1915 9948
rect 1857 9939 1915 9945
rect 3050 9936 3056 9948
rect 3108 9936 3114 9988
rect 3160 9976 3188 10016
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 3436 9976 3464 10007
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5592 10016 5733 10044
rect 5592 10004 5598 10016
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 6840 10044 6868 10072
rect 8570 10044 8576 10056
rect 6840 10016 8576 10044
rect 5721 10007 5779 10013
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 16022 10044 16028 10056
rect 15983 10016 16028 10044
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 7098 9976 7104 9988
rect 3160 9948 3464 9976
rect 7011 9948 7104 9976
rect 2314 9868 2320 9920
rect 2372 9908 2378 9920
rect 2869 9911 2927 9917
rect 2869 9908 2881 9911
rect 2372 9880 2881 9908
rect 2372 9868 2378 9880
rect 2869 9877 2881 9880
rect 2915 9877 2927 9911
rect 3436 9908 3464 9948
rect 7098 9936 7104 9948
rect 7156 9976 7162 9988
rect 9401 9979 9459 9985
rect 9401 9976 9413 9979
rect 7156 9948 9413 9976
rect 7156 9936 7162 9948
rect 9401 9945 9413 9948
rect 9447 9945 9459 9979
rect 9401 9939 9459 9945
rect 14737 9979 14795 9985
rect 14737 9945 14749 9979
rect 14783 9976 14795 9979
rect 15102 9976 15108 9988
rect 14783 9948 15108 9976
rect 14783 9945 14795 9948
rect 14737 9939 14795 9945
rect 15102 9936 15108 9948
rect 15160 9936 15166 9988
rect 3878 9908 3884 9920
rect 3436 9880 3884 9908
rect 2869 9871 2927 9877
rect 3878 9868 3884 9880
rect 3936 9908 3942 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 3936 9880 5457 9908
rect 3936 9868 3942 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 5445 9871 5503 9877
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 6914 9908 6920 9920
rect 6144 9880 6920 9908
rect 6144 9868 6150 9880
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 7377 9911 7435 9917
rect 7377 9908 7389 9911
rect 7248 9880 7389 9908
rect 7248 9868 7254 9880
rect 7377 9877 7389 9880
rect 7423 9877 7435 9911
rect 7377 9871 7435 9877
rect 7650 9868 7656 9920
rect 7708 9908 7714 9920
rect 7745 9911 7803 9917
rect 7745 9908 7757 9911
rect 7708 9880 7757 9908
rect 7708 9868 7714 9880
rect 7745 9877 7757 9880
rect 7791 9877 7803 9911
rect 7745 9871 7803 9877
rect 9953 9911 10011 9917
rect 9953 9877 9965 9911
rect 9999 9908 10011 9911
rect 10962 9908 10968 9920
rect 9999 9880 10968 9908
rect 9999 9877 10011 9880
rect 9953 9871 10011 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11425 9911 11483 9917
rect 11425 9877 11437 9911
rect 11471 9908 11483 9911
rect 11974 9908 11980 9920
rect 11471 9880 11980 9908
rect 11471 9877 11483 9880
rect 11425 9871 11483 9877
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 15381 9911 15439 9917
rect 15381 9877 15393 9911
rect 15427 9908 15439 9911
rect 17034 9908 17040 9920
rect 15427 9880 17040 9908
rect 15427 9877 15439 9880
rect 15381 9871 15439 9877
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 1762 9704 1768 9716
rect 1723 9676 1768 9704
rect 1762 9664 1768 9676
rect 1820 9664 1826 9716
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 2556 9676 2820 9704
rect 2556 9664 2562 9676
rect 1780 9568 1808 9664
rect 2792 9636 2820 9676
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 3418 9704 3424 9716
rect 2924 9676 3424 9704
rect 2924 9664 2930 9676
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 15654 9704 15660 9716
rect 4120 9676 15660 9704
rect 4120 9664 4126 9676
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 15838 9664 15844 9716
rect 15896 9704 15902 9716
rect 16393 9707 16451 9713
rect 16393 9704 16405 9707
rect 15896 9676 16405 9704
rect 15896 9664 15902 9676
rect 16393 9673 16405 9676
rect 16439 9673 16451 9707
rect 16393 9667 16451 9673
rect 17402 9664 17408 9716
rect 17460 9704 17466 9716
rect 17589 9707 17647 9713
rect 17589 9704 17601 9707
rect 17460 9676 17601 9704
rect 17460 9664 17466 9676
rect 17589 9673 17601 9676
rect 17635 9673 17647 9707
rect 17589 9667 17647 9673
rect 18693 9707 18751 9713
rect 18693 9673 18705 9707
rect 18739 9704 18751 9707
rect 19610 9704 19616 9716
rect 18739 9676 19616 9704
rect 18739 9673 18751 9676
rect 18693 9667 18751 9673
rect 19610 9664 19616 9676
rect 19668 9664 19674 9716
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 2792 9608 4537 9636
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 4525 9599 4583 9605
rect 5074 9596 5080 9648
rect 5132 9636 5138 9648
rect 5537 9639 5595 9645
rect 5537 9636 5549 9639
rect 5132 9608 5549 9636
rect 5132 9596 5138 9608
rect 5537 9605 5549 9608
rect 5583 9636 5595 9639
rect 6546 9636 6552 9648
rect 5583 9608 6552 9636
rect 5583 9605 5595 9608
rect 5537 9599 5595 9605
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 6972 9608 7420 9636
rect 6972 9596 6978 9608
rect 4062 9568 4068 9580
rect 1780 9540 1992 9568
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9469 1915 9503
rect 1964 9500 1992 9540
rect 3896 9540 4068 9568
rect 2113 9503 2171 9509
rect 2113 9500 2125 9503
rect 1964 9472 2125 9500
rect 1857 9463 1915 9469
rect 2113 9469 2125 9472
rect 2159 9469 2171 9503
rect 2682 9500 2688 9512
rect 2113 9463 2171 9469
rect 2240 9472 2688 9500
rect 1872 9432 1900 9463
rect 2240 9432 2268 9472
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 3896 9509 3924 9540
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 4203 9540 5181 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 5169 9537 5181 9540
rect 5215 9568 5227 9571
rect 5718 9568 5724 9580
rect 5215 9540 5724 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 7098 9568 7104 9580
rect 6411 9540 7104 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7392 9577 7420 9608
rect 9950 9596 9956 9648
rect 10008 9636 10014 9648
rect 10134 9636 10140 9648
rect 10008 9608 10140 9636
rect 10008 9596 10014 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 11425 9639 11483 9645
rect 11425 9636 11437 9639
rect 10796 9608 11437 9636
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 8202 9568 8208 9580
rect 7708 9540 8208 9568
rect 7708 9528 7714 9540
rect 8202 9528 8208 9540
rect 8260 9568 8266 9580
rect 10796 9577 10824 9608
rect 11425 9605 11437 9608
rect 11471 9636 11483 9639
rect 12434 9636 12440 9648
rect 11471 9608 12440 9636
rect 11471 9605 11483 9608
rect 11425 9599 11483 9605
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 13633 9639 13691 9645
rect 13633 9605 13645 9639
rect 13679 9636 13691 9639
rect 13814 9636 13820 9648
rect 13679 9608 13820 9636
rect 13679 9605 13691 9608
rect 13633 9599 13691 9605
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14550 9636 14556 9648
rect 14384 9608 14556 9636
rect 8665 9571 8723 9577
rect 8665 9568 8677 9571
rect 8260 9540 8677 9568
rect 8260 9528 8266 9540
rect 8665 9537 8677 9540
rect 8711 9537 8723 9571
rect 8665 9531 8723 9537
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10962 9568 10968 9580
rect 10923 9540 10968 9568
rect 10781 9531 10839 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12768 9540 12909 9568
rect 12768 9528 12774 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 12897 9531 12955 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 14384 9577 14412 9608
rect 14550 9596 14556 9608
rect 14608 9636 14614 9648
rect 14829 9639 14887 9645
rect 14829 9636 14841 9639
rect 14608 9608 14841 9636
rect 14608 9596 14614 9608
rect 14829 9605 14841 9608
rect 14875 9605 14887 9639
rect 14829 9599 14887 9605
rect 15672 9577 15700 9664
rect 16577 9639 16635 9645
rect 16577 9605 16589 9639
rect 16623 9636 16635 9639
rect 19150 9636 19156 9648
rect 16623 9608 19156 9636
rect 16623 9605 16635 9608
rect 16577 9599 16635 9605
rect 19150 9596 19156 9608
rect 19208 9596 19214 9648
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 15657 9571 15715 9577
rect 15657 9537 15669 9571
rect 15703 9537 15715 9571
rect 17126 9568 17132 9580
rect 17087 9540 17132 9568
rect 15657 9531 15715 9537
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17770 9528 17776 9580
rect 17828 9568 17834 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 17828 9540 18245 9568
rect 17828 9528 17834 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9568 19119 9571
rect 19334 9568 19340 9580
rect 19107 9540 19340 9568
rect 19107 9537 19119 9540
rect 19061 9531 19119 9537
rect 19334 9528 19340 9540
rect 19392 9568 19398 9580
rect 19978 9568 19984 9580
rect 19392 9540 19984 9568
rect 19392 9528 19398 9540
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9469 3939 9503
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 3881 9463 3939 9469
rect 3988 9472 5457 9500
rect 1872 9404 2268 9432
rect 2498 9392 2504 9444
rect 2556 9432 2562 9444
rect 3988 9432 4016 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 6546 9500 6552 9512
rect 6135 9472 6552 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 6546 9460 6552 9472
rect 6604 9460 6610 9512
rect 7190 9500 7196 9512
rect 7151 9472 7196 9500
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7466 9460 7472 9512
rect 7524 9500 7530 9512
rect 7524 9472 10824 9500
rect 7524 9460 7530 9472
rect 5810 9432 5816 9444
rect 2556 9404 4016 9432
rect 4080 9404 5816 9432
rect 2556 9392 2562 9404
rect 4080 9376 4108 9404
rect 5810 9392 5816 9404
rect 5868 9432 5874 9444
rect 6454 9432 6460 9444
rect 5868 9404 6460 9432
rect 5868 9392 5874 9404
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 8932 9435 8990 9441
rect 8932 9401 8944 9435
rect 8978 9432 8990 9435
rect 9674 9432 9680 9444
rect 8978 9404 9680 9432
rect 8978 9401 8990 9404
rect 8932 9395 8990 9401
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 10796 9432 10824 9472
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 11514 9500 11520 9512
rect 10928 9472 11520 9500
rect 10928 9460 10934 9472
rect 11514 9460 11520 9472
rect 11572 9500 11578 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11572 9472 11713 9500
rect 11572 9460 11578 9472
rect 11701 9469 11713 9472
rect 11747 9500 11759 9503
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 11747 9472 12081 9500
rect 11747 9469 11759 9472
rect 11701 9463 11759 9469
rect 12069 9469 12081 9472
rect 12115 9469 12127 9503
rect 12802 9500 12808 9512
rect 12763 9472 12808 9500
rect 12069 9463 12127 9469
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 14185 9503 14243 9509
rect 14185 9469 14197 9503
rect 14231 9500 14243 9503
rect 15194 9500 15200 9512
rect 14231 9472 15200 9500
rect 14231 9469 14243 9472
rect 14185 9463 14243 9469
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 16945 9503 17003 9509
rect 16945 9469 16957 9503
rect 16991 9500 17003 9503
rect 17402 9500 17408 9512
rect 16991 9472 17408 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 16298 9432 16304 9444
rect 10796 9404 16304 9432
rect 16298 9392 16304 9404
rect 16356 9392 16362 9444
rect 17034 9432 17040 9444
rect 16995 9404 17040 9432
rect 17034 9392 17040 9404
rect 17092 9392 17098 9444
rect 3234 9364 3240 9376
rect 3195 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3510 9364 3516 9376
rect 3471 9336 3516 9364
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 3973 9367 4031 9373
rect 3973 9333 3985 9367
rect 4019 9364 4031 9367
rect 4062 9364 4068 9376
rect 4019 9336 4068 9364
rect 4019 9333 4031 9336
rect 3973 9327 4031 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 4893 9367 4951 9373
rect 4893 9364 4905 9367
rect 4764 9336 4905 9364
rect 4764 9324 4770 9336
rect 4893 9333 4905 9336
rect 4939 9333 4951 9367
rect 4893 9327 4951 9333
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 5074 9364 5080 9376
rect 5031 9336 5080 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5445 9367 5503 9373
rect 5445 9333 5457 9367
rect 5491 9364 5503 9367
rect 5721 9367 5779 9373
rect 5721 9364 5733 9367
rect 5491 9336 5733 9364
rect 5491 9333 5503 9336
rect 5445 9327 5503 9333
rect 5721 9333 5733 9336
rect 5767 9333 5779 9367
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 5721 9327 5779 9333
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 6604 9336 6837 9364
rect 6604 9324 6610 9336
rect 6825 9333 6837 9336
rect 6871 9333 6883 9367
rect 6825 9327 6883 9333
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6972 9336 7297 9364
rect 6972 9324 6978 9336
rect 7285 9333 7297 9336
rect 7331 9364 7343 9367
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7331 9336 7849 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 8113 9367 8171 9373
rect 8113 9333 8125 9367
rect 8159 9364 8171 9367
rect 9490 9364 9496 9376
rect 8159 9336 9496 9364
rect 8159 9333 8171 9336
rect 8113 9327 8171 9333
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 9582 9324 9588 9376
rect 9640 9364 9646 9376
rect 9858 9364 9864 9376
rect 9640 9336 9864 9364
rect 9640 9324 9646 9336
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 10042 9364 10048 9376
rect 10003 9336 10048 9364
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10318 9364 10324 9376
rect 10279 9336 10324 9364
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10689 9367 10747 9373
rect 10689 9333 10701 9367
rect 10735 9364 10747 9367
rect 10778 9364 10784 9376
rect 10735 9336 10784 9364
rect 10735 9333 10747 9336
rect 10689 9327 10747 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12492 9336 12537 9364
rect 12492 9324 12498 9336
rect 15102 9324 15108 9376
rect 15160 9364 15166 9376
rect 15197 9367 15255 9373
rect 15197 9364 15209 9367
rect 15160 9336 15209 9364
rect 15160 9324 15166 9336
rect 15197 9333 15209 9336
rect 15243 9333 15255 9367
rect 15197 9327 15255 9333
rect 15930 9324 15936 9376
rect 15988 9364 15994 9376
rect 16025 9367 16083 9373
rect 16025 9364 16037 9367
rect 15988 9336 16037 9364
rect 15988 9324 15994 9336
rect 16025 9333 16037 9336
rect 16071 9333 16083 9367
rect 16025 9327 16083 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2280 9132 2329 9160
rect 2280 9120 2286 9132
rect 2317 9129 2329 9132
rect 2363 9160 2375 9163
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2363 9132 2789 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 2777 9123 2835 9129
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 5718 9160 5724 9172
rect 3559 9132 5724 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 5718 9120 5724 9132
rect 5776 9160 5782 9172
rect 5997 9163 6055 9169
rect 5997 9160 6009 9163
rect 5776 9132 6009 9160
rect 5776 9120 5782 9132
rect 5997 9129 6009 9132
rect 6043 9129 6055 9163
rect 6362 9160 6368 9172
rect 6323 9132 6368 9160
rect 5997 9123 6055 9129
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9160 6607 9163
rect 7190 9160 7196 9172
rect 6595 9132 7196 9160
rect 6595 9129 6607 9132
rect 6549 9123 6607 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7374 9160 7380 9172
rect 7331 9132 7380 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 8628 9132 9873 9160
rect 8628 9120 8634 9132
rect 9861 9129 9873 9132
rect 9907 9160 9919 9163
rect 10042 9160 10048 9172
rect 9907 9132 10048 9160
rect 9907 9129 9919 9132
rect 9861 9123 9919 9129
rect 10042 9120 10048 9132
rect 10100 9160 10106 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 10100 9132 10241 9160
rect 10100 9120 10106 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11057 9163 11115 9169
rect 11057 9160 11069 9163
rect 11020 9132 11069 9160
rect 11020 9120 11026 9132
rect 11057 9129 11069 9132
rect 11103 9129 11115 9163
rect 11514 9160 11520 9172
rect 11475 9132 11520 9160
rect 11057 9123 11115 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 12802 9160 12808 9172
rect 12763 9132 12808 9160
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 13136 9132 13185 9160
rect 13136 9120 13142 9132
rect 13173 9129 13185 9132
rect 13219 9160 13231 9163
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 13219 9132 13553 9160
rect 13219 9129 13231 9132
rect 13173 9123 13231 9129
rect 13541 9129 13553 9132
rect 13587 9129 13599 9163
rect 13541 9123 13599 9129
rect 14461 9163 14519 9169
rect 14461 9129 14473 9163
rect 14507 9160 14519 9163
rect 15102 9160 15108 9172
rect 14507 9132 15108 9160
rect 14507 9129 14519 9132
rect 14461 9123 14519 9129
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 15470 9120 15476 9172
rect 15528 9160 15534 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 15528 9132 15669 9160
rect 15528 9120 15534 9132
rect 15657 9129 15669 9132
rect 15703 9160 15715 9163
rect 16025 9163 16083 9169
rect 16025 9160 16037 9163
rect 15703 9132 16037 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 16025 9129 16037 9132
rect 16071 9129 16083 9163
rect 16025 9123 16083 9129
rect 17037 9163 17095 9169
rect 17037 9129 17049 9163
rect 17083 9160 17095 9163
rect 17126 9160 17132 9172
rect 17083 9132 17132 9160
rect 17083 9129 17095 9132
rect 17037 9123 17095 9129
rect 17126 9120 17132 9132
rect 17184 9160 17190 9172
rect 17313 9163 17371 9169
rect 17313 9160 17325 9163
rect 17184 9132 17325 9160
rect 17184 9120 17190 9132
rect 17313 9129 17325 9132
rect 17359 9129 17371 9163
rect 17313 9123 17371 9129
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 18141 9163 18199 9169
rect 18141 9160 18153 9163
rect 17552 9132 18153 9160
rect 17552 9120 17558 9132
rect 18141 9129 18153 9132
rect 18187 9160 18199 9163
rect 19334 9160 19340 9172
rect 18187 9132 19340 9160
rect 18187 9129 18199 9132
rect 18141 9123 18199 9129
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 1673 9095 1731 9101
rect 1673 9061 1685 9095
rect 1719 9092 1731 9095
rect 3326 9092 3332 9104
rect 1719 9064 3332 9092
rect 1719 9061 1731 9064
rect 1673 9055 1731 9061
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 14829 9095 14887 9101
rect 4212 9064 13308 9092
rect 4212 9052 4218 9064
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 9024 1823 9027
rect 2130 9024 2136 9036
rect 1811 8996 2136 9024
rect 1811 8993 1823 8996
rect 1765 8987 1823 8993
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 5350 9024 5356 9036
rect 3016 8996 5356 9024
rect 3016 8984 3022 8996
rect 5350 8984 5356 8996
rect 5408 9024 5414 9036
rect 6822 9024 6828 9036
rect 5408 8996 6828 9024
rect 5408 8984 5414 8996
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 8849 9027 8907 9033
rect 8849 8993 8861 9027
rect 8895 9024 8907 9027
rect 9030 9024 9036 9036
rect 8895 8996 9036 9024
rect 8895 8993 8907 8996
rect 8849 8987 8907 8993
rect 9030 8984 9036 8996
rect 9088 9024 9094 9036
rect 9582 9024 9588 9036
rect 9088 8996 9588 9024
rect 9088 8984 9094 8996
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 13280 9024 13308 9064
rect 14829 9061 14841 9095
rect 14875 9092 14887 9095
rect 15010 9092 15016 9104
rect 14875 9064 15016 9092
rect 14875 9061 14887 9064
rect 14829 9055 14887 9061
rect 15010 9052 15016 9064
rect 15068 9052 15074 9104
rect 16850 9092 16856 9104
rect 15120 9064 16856 9092
rect 15120 9024 15148 9064
rect 16850 9052 16856 9064
rect 16908 9052 16914 9104
rect 13280 8996 15148 9024
rect 16022 8984 16028 9036
rect 16080 9024 16086 9036
rect 16393 9027 16451 9033
rect 16393 9024 16405 9027
rect 16080 8996 16405 9024
rect 16080 8984 16086 8996
rect 16393 8993 16405 8996
rect 16439 8993 16451 9027
rect 16393 8987 16451 8993
rect 17034 8984 17040 9036
rect 17092 9024 17098 9036
rect 17681 9027 17739 9033
rect 17681 9024 17693 9027
rect 17092 8996 17693 9024
rect 17092 8984 17098 8996
rect 17681 8993 17693 8996
rect 17727 8993 17739 9027
rect 17681 8987 17739 8993
rect 2498 8916 2504 8968
rect 2556 8956 2562 8968
rect 6914 8956 6920 8968
rect 2556 8928 6920 8956
rect 2556 8916 2562 8928
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 7699 8928 8309 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 8297 8925 8309 8928
rect 8343 8956 8355 8959
rect 8478 8956 8484 8968
rect 8343 8928 8484 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8956 9183 8959
rect 9674 8956 9680 8968
rect 9171 8928 9680 8956
rect 9171 8925 9183 8928
rect 9125 8919 9183 8925
rect 1026 8848 1032 8900
rect 1084 8888 1090 8900
rect 4062 8888 4068 8900
rect 1084 8860 4068 8888
rect 1084 8848 1090 8860
rect 4062 8848 4068 8860
rect 4120 8888 4126 8900
rect 4341 8891 4399 8897
rect 4341 8888 4353 8891
rect 4120 8860 4353 8888
rect 4120 8848 4126 8860
rect 4341 8857 4353 8860
rect 4387 8857 4399 8891
rect 4341 8851 4399 8857
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 8956 8888 8984 8919
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 10744 8928 12449 8956
rect 10744 8916 10750 8928
rect 12437 8925 12449 8928
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 5040 8860 8984 8888
rect 5040 8848 5046 8860
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 3142 8820 3148 8832
rect 1995 8792 3148 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 3881 8823 3939 8829
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 4246 8820 4252 8832
rect 3927 8792 4252 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4764 8792 4905 8820
rect 4764 8780 4770 8792
rect 4893 8789 4905 8792
rect 4939 8820 4951 8823
rect 5074 8820 5080 8832
rect 4939 8792 5080 8820
rect 4939 8789 4951 8792
rect 4893 8783 4951 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5350 8820 5356 8832
rect 5311 8792 5356 8820
rect 5350 8780 5356 8792
rect 5408 8820 5414 8832
rect 6270 8820 6276 8832
rect 5408 8792 6276 8820
rect 5408 8780 5414 8792
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 8481 8823 8539 8829
rect 8481 8789 8493 8823
rect 8527 8820 8539 8823
rect 8754 8820 8760 8832
rect 8527 8792 8760 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 8956 8820 8984 8860
rect 9214 8848 9220 8900
rect 9272 8888 9278 8900
rect 10778 8888 10784 8900
rect 9272 8860 10784 8888
rect 9272 8848 9278 8860
rect 10778 8848 10784 8860
rect 10836 8848 10842 8900
rect 10134 8820 10140 8832
rect 8956 8792 10140 8820
rect 10134 8780 10140 8792
rect 10192 8780 10198 8832
rect 11885 8823 11943 8829
rect 11885 8789 11897 8823
rect 11931 8820 11943 8823
rect 11974 8820 11980 8832
rect 11931 8792 11980 8820
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 13722 8780 13728 8832
rect 13780 8820 13786 8832
rect 13909 8823 13967 8829
rect 13909 8820 13921 8823
rect 13780 8792 13921 8820
rect 13780 8780 13786 8792
rect 13909 8789 13921 8792
rect 13955 8789 13967 8823
rect 13909 8783 13967 8789
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 3510 8616 3516 8628
rect 1811 8588 3516 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 3878 8616 3884 8628
rect 3839 8588 3884 8616
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 5166 8616 5172 8628
rect 4304 8588 5172 8616
rect 4304 8576 4310 8588
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 6914 8616 6920 8628
rect 6875 8588 6920 8616
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9674 8616 9680 8628
rect 9355 8588 9680 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9674 8576 9680 8588
rect 9732 8616 9738 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 9732 8588 10425 8616
rect 9732 8576 9738 8588
rect 10413 8585 10425 8588
rect 10459 8616 10471 8619
rect 10962 8616 10968 8628
rect 10459 8588 10968 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11974 8616 11980 8628
rect 11935 8588 11980 8616
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13173 8619 13231 8625
rect 13173 8616 13185 8619
rect 12952 8588 13185 8616
rect 12952 8576 12958 8588
rect 13173 8585 13185 8588
rect 13219 8585 13231 8619
rect 13722 8616 13728 8628
rect 13683 8588 13728 8616
rect 13173 8579 13231 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 14458 8616 14464 8628
rect 14419 8588 14464 8616
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 16022 8616 16028 8628
rect 15983 8588 16028 8616
rect 16022 8576 16028 8588
rect 16080 8576 16086 8628
rect 16390 8616 16396 8628
rect 16351 8588 16396 8616
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 16850 8616 16856 8628
rect 16763 8588 16856 8616
rect 16850 8576 16856 8588
rect 16908 8616 16914 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 16908 8588 17233 8616
rect 16908 8576 16914 8588
rect 17221 8585 17233 8588
rect 17267 8616 17279 8619
rect 17494 8616 17500 8628
rect 17267 8588 17500 8616
rect 17267 8585 17279 8588
rect 17221 8579 17279 8585
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8517 3663 8551
rect 3605 8511 3663 8517
rect 10045 8551 10103 8557
rect 10045 8517 10057 8551
rect 10091 8548 10103 8551
rect 10134 8548 10140 8560
rect 10091 8520 10140 8548
rect 10091 8517 10103 8520
rect 10045 8511 10103 8517
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3620 8480 3648 8511
rect 10134 8508 10140 8520
rect 10192 8508 10198 8560
rect 10686 8548 10692 8560
rect 10647 8520 10692 8548
rect 10686 8508 10692 8520
rect 10744 8508 10750 8560
rect 11701 8551 11759 8557
rect 11701 8517 11713 8551
rect 11747 8548 11759 8551
rect 12158 8548 12164 8560
rect 11747 8520 12164 8548
rect 11747 8517 11759 8520
rect 11701 8511 11759 8517
rect 12158 8508 12164 8520
rect 12216 8548 12222 8560
rect 12805 8551 12863 8557
rect 12805 8548 12817 8551
rect 12216 8520 12817 8548
rect 12216 8508 12222 8520
rect 12805 8517 12817 8520
rect 12851 8517 12863 8551
rect 12805 8511 12863 8517
rect 13998 8508 14004 8560
rect 14056 8548 14062 8560
rect 14737 8551 14795 8557
rect 14737 8548 14749 8551
rect 14056 8520 14749 8548
rect 14056 8508 14062 8520
rect 14737 8517 14749 8520
rect 14783 8517 14795 8551
rect 14737 8511 14795 8517
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 3384 8452 5365 8480
rect 3384 8440 3390 8452
rect 5353 8449 5365 8452
rect 5399 8480 5411 8483
rect 6089 8483 6147 8489
rect 6089 8480 6101 8483
rect 5399 8452 6101 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 6089 8449 6101 8452
rect 6135 8449 6147 8483
rect 6089 8443 6147 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 7098 8480 7104 8492
rect 6595 8452 7104 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 7607 8452 8064 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 2056 8384 2237 8412
rect 2056 8276 2084 8384
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 3234 8412 3240 8424
rect 2225 8375 2283 8381
rect 2516 8384 3240 8412
rect 2516 8353 2544 8384
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 7282 8412 7288 8424
rect 7243 8384 7288 8412
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 7926 8412 7932 8424
rect 7887 8384 7932 8412
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 2470 8347 2544 8353
rect 2470 8344 2482 8347
rect 2179 8316 2482 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 2470 8313 2482 8316
rect 2516 8316 2544 8347
rect 2682 8344 2688 8356
rect 2608 8316 2688 8344
rect 2516 8313 2528 8316
rect 2470 8307 2528 8313
rect 2608 8276 2636 8316
rect 2682 8304 2688 8316
rect 2740 8344 2746 8356
rect 2866 8344 2872 8356
rect 2740 8316 2872 8344
rect 2740 8304 2746 8316
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 5077 8347 5135 8353
rect 5077 8344 5089 8347
rect 3252 8316 5089 8344
rect 3252 8288 3280 8316
rect 5077 8313 5089 8316
rect 5123 8313 5135 8347
rect 5077 8307 5135 8313
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8344 5227 8347
rect 5810 8344 5816 8356
rect 5215 8316 5816 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 2056 8248 2636 8276
rect 3234 8236 3240 8288
rect 3292 8236 3298 8288
rect 4246 8276 4252 8288
rect 4207 8248 4252 8276
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4706 8276 4712 8288
rect 4667 8248 4712 8276
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 5092 8276 5120 8307
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7377 8347 7435 8353
rect 7377 8344 7389 8347
rect 6972 8316 7389 8344
rect 6972 8304 6978 8316
rect 7377 8313 7389 8316
rect 7423 8313 7435 8347
rect 7377 8307 7435 8313
rect 5350 8276 5356 8288
rect 5092 8248 5356 8276
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 7098 8236 7104 8288
rect 7156 8276 7162 8288
rect 7944 8276 7972 8372
rect 8036 8344 8064 8452
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 8996 8452 14136 8480
rect 8996 8440 9002 8452
rect 8196 8347 8254 8353
rect 8196 8344 8208 8347
rect 8036 8316 8208 8344
rect 8196 8313 8208 8316
rect 8242 8344 8254 8347
rect 8478 8344 8484 8356
rect 8242 8316 8484 8344
rect 8242 8313 8254 8316
rect 8196 8307 8254 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 11882 8304 11888 8356
rect 11940 8344 11946 8356
rect 14001 8347 14059 8353
rect 14001 8344 14013 8347
rect 11940 8316 14013 8344
rect 11940 8304 11946 8316
rect 14001 8313 14013 8316
rect 14047 8313 14059 8347
rect 14108 8344 14136 8452
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14424 8452 15117 8480
rect 14424 8440 14430 8452
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 15473 8415 15531 8421
rect 15473 8412 15485 8415
rect 14332 8384 15485 8412
rect 14332 8372 14338 8384
rect 15473 8381 15485 8384
rect 15519 8381 15531 8415
rect 15473 8375 15531 8381
rect 17310 8344 17316 8356
rect 14108 8316 17316 8344
rect 14001 8307 14059 8313
rect 17310 8304 17316 8316
rect 17368 8304 17374 8356
rect 9582 8276 9588 8288
rect 7156 8248 7972 8276
rect 9543 8248 9588 8276
rect 7156 8236 7162 8248
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 11974 8276 11980 8288
rect 11756 8248 11980 8276
rect 11756 8236 11762 8248
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 1673 8075 1731 8081
rect 1673 8041 1685 8075
rect 1719 8072 1731 8075
rect 2774 8072 2780 8084
rect 1719 8044 2780 8072
rect 1719 8041 1731 8044
rect 1673 8035 1731 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 4246 8072 4252 8084
rect 3375 8044 4252 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 7282 8072 7288 8084
rect 5132 8044 7288 8072
rect 5132 8032 5138 8044
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 8202 8072 8208 8084
rect 7708 8044 8208 8072
rect 7708 8032 7714 8044
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 8478 8072 8484 8084
rect 8439 8044 8484 8072
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 8720 8044 9873 8072
rect 8720 8032 8726 8044
rect 9861 8041 9873 8044
rect 9907 8041 9919 8075
rect 9861 8035 9919 8041
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 11701 8075 11759 8081
rect 11701 8072 11713 8075
rect 10376 8044 11713 8072
rect 10376 8032 10382 8044
rect 11701 8041 11713 8044
rect 11747 8041 11759 8075
rect 12066 8072 12072 8084
rect 12027 8044 12072 8072
rect 11701 8035 11759 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 12986 8072 12992 8084
rect 12575 8044 12992 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 13265 8075 13323 8081
rect 13265 8041 13277 8075
rect 13311 8072 13323 8075
rect 13354 8072 13360 8084
rect 13311 8044 13360 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 13538 8072 13544 8084
rect 13499 8044 13544 8072
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 13906 8072 13912 8084
rect 13867 8044 13912 8072
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14332 8044 14657 8072
rect 14332 8032 14338 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 14645 8035 14703 8041
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 15933 8075 15991 8081
rect 15933 8072 15945 8075
rect 15611 8044 15945 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 15933 8041 15945 8044
rect 15979 8072 15991 8075
rect 16850 8072 16856 8084
rect 15979 8044 16856 8072
rect 15979 8041 15991 8044
rect 15933 8035 15991 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 3142 7964 3148 8016
rect 3200 8004 3206 8016
rect 3786 8004 3792 8016
rect 3200 7976 3792 8004
rect 3200 7964 3206 7976
rect 3786 7964 3792 7976
rect 3844 7964 3850 8016
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 12253 8007 12311 8013
rect 12253 8004 12265 8007
rect 4120 7976 12265 8004
rect 4120 7964 4126 7976
rect 12253 7973 12265 7976
rect 12299 7973 12311 8007
rect 12253 7967 12311 7973
rect 1489 7939 1547 7945
rect 1489 7905 1501 7939
rect 1535 7905 1547 7939
rect 1489 7899 1547 7905
rect 2041 7939 2099 7945
rect 2041 7905 2053 7939
rect 2087 7936 2099 7939
rect 2774 7936 2780 7948
rect 2087 7908 2780 7936
rect 2087 7905 2099 7908
rect 2041 7899 2099 7905
rect 1504 7868 1532 7899
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3421 7939 3479 7945
rect 3421 7936 3433 7939
rect 3016 7908 3433 7936
rect 3016 7896 3022 7908
rect 3421 7905 3433 7908
rect 3467 7905 3479 7939
rect 3421 7899 3479 7905
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4212 7908 4445 7936
rect 4212 7896 4218 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 4433 7899 4491 7905
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7936 4583 7939
rect 4706 7936 4712 7948
rect 4571 7908 4712 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 5350 7945 5356 7948
rect 5344 7936 5356 7945
rect 5311 7908 5356 7936
rect 5344 7899 5356 7908
rect 5350 7896 5356 7899
rect 5408 7896 5414 7948
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 7098 7936 7104 7948
rect 6880 7908 7104 7936
rect 6880 7896 6886 7908
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7368 7939 7426 7945
rect 7368 7905 7380 7939
rect 7414 7936 7426 7939
rect 7742 7936 7748 7948
rect 7414 7908 7748 7936
rect 7414 7905 7426 7908
rect 7368 7899 7426 7905
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 12158 7936 12164 7948
rect 7892 7908 12164 7936
rect 7892 7896 7898 7908
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 12805 7939 12863 7945
rect 12805 7936 12817 7939
rect 12768 7908 12817 7936
rect 12768 7896 12774 7908
rect 12805 7905 12817 7908
rect 12851 7905 12863 7939
rect 12805 7899 12863 7905
rect 2314 7868 2320 7880
rect 1504 7840 2320 7868
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 3513 7871 3571 7877
rect 3513 7868 3525 7871
rect 2915 7840 3525 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3513 7837 3525 7840
rect 3559 7868 3571 7871
rect 3786 7868 3792 7880
rect 3559 7840 3792 7868
rect 3559 7837 3571 7840
rect 3513 7831 3571 7837
rect 3786 7828 3792 7840
rect 3844 7868 3850 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 3844 7840 4629 7868
rect 3844 7828 3850 7840
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 5074 7868 5080 7880
rect 5035 7840 5080 7868
rect 4617 7831 4675 7837
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 10502 7868 10508 7880
rect 8260 7840 10508 7868
rect 8260 7828 8266 7840
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 10735 7840 11345 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 11333 7837 11345 7840
rect 11379 7868 11391 7871
rect 11882 7868 11888 7880
rect 11379 7840 11888 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 12032 7840 14289 7868
rect 12032 7828 12038 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 1118 7760 1124 7812
rect 1176 7800 1182 7812
rect 3234 7800 3240 7812
rect 1176 7772 3240 7800
rect 1176 7760 1182 7772
rect 3234 7760 3240 7772
rect 3292 7760 3298 7812
rect 8938 7800 8944 7812
rect 8851 7772 8944 7800
rect 8938 7760 8944 7772
rect 8996 7800 9002 7812
rect 10962 7800 10968 7812
rect 8996 7772 10968 7800
rect 8996 7760 9002 7772
rect 10962 7760 10968 7772
rect 11020 7760 11026 7812
rect 11057 7803 11115 7809
rect 11057 7769 11069 7803
rect 11103 7800 11115 7803
rect 12253 7803 12311 7809
rect 11103 7772 12204 7800
rect 11103 7769 11115 7772
rect 11057 7763 11115 7769
rect 2958 7732 2964 7744
rect 2919 7704 2964 7732
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 4028 7704 4077 7732
rect 4028 7692 4034 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 6457 7735 6515 7741
rect 6457 7701 6469 7735
rect 6503 7732 6515 7735
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 6503 7704 6929 7732
rect 6503 7701 6515 7704
rect 6457 7695 6515 7701
rect 6917 7701 6929 7704
rect 6963 7732 6975 7735
rect 7006 7732 7012 7744
rect 6963 7704 7012 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 9217 7735 9275 7741
rect 9217 7732 9229 7735
rect 8904 7704 9229 7732
rect 8904 7692 8910 7704
rect 9217 7701 9229 7704
rect 9263 7701 9275 7735
rect 9217 7695 9275 7701
rect 9950 7692 9956 7744
rect 10008 7732 10014 7744
rect 10229 7735 10287 7741
rect 10229 7732 10241 7735
rect 10008 7704 10241 7732
rect 10008 7692 10014 7704
rect 10229 7701 10241 7704
rect 10275 7701 10287 7735
rect 12176 7732 12204 7772
rect 12253 7769 12265 7803
rect 12299 7800 12311 7803
rect 15930 7800 15936 7812
rect 12299 7772 15936 7800
rect 12299 7769 12311 7772
rect 12253 7763 12311 7769
rect 15930 7760 15936 7772
rect 15988 7760 15994 7812
rect 12894 7732 12900 7744
rect 12176 7704 12900 7732
rect 10229 7695 10287 7701
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 15010 7732 15016 7744
rect 14971 7704 15016 7732
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7528 1823 7531
rect 1946 7528 1952 7540
rect 1811 7500 1952 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 3844 7500 4445 7528
rect 3844 7488 3850 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 4433 7491 4491 7497
rect 4617 7531 4675 7537
rect 4617 7497 4629 7531
rect 4663 7528 4675 7531
rect 5074 7528 5080 7540
rect 4663 7500 5080 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 3053 7395 3111 7401
rect 3053 7392 3065 7395
rect 2924 7364 3065 7392
rect 2924 7352 2930 7364
rect 3053 7361 3065 7364
rect 3099 7361 3111 7395
rect 4448 7392 4476 7491
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 9493 7531 9551 7537
rect 9493 7528 9505 7531
rect 7064 7500 9505 7528
rect 7064 7488 7070 7500
rect 9493 7497 9505 7500
rect 9539 7497 9551 7531
rect 9493 7491 9551 7497
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 11241 7531 11299 7537
rect 11241 7528 11253 7531
rect 10560 7500 11253 7528
rect 10560 7488 10566 7500
rect 11241 7497 11253 7500
rect 11287 7497 11299 7531
rect 11241 7491 11299 7497
rect 11606 7488 11612 7540
rect 11664 7528 11670 7540
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11664 7500 11805 7528
rect 11664 7488 11670 7500
rect 11793 7497 11805 7500
rect 11839 7497 11851 7531
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 11793 7491 11851 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 12713 7531 12771 7537
rect 12713 7528 12725 7531
rect 12676 7500 12725 7528
rect 12676 7488 12682 7500
rect 12713 7497 12725 7500
rect 12759 7497 12771 7531
rect 13170 7528 13176 7540
rect 13131 7500 13176 7528
rect 12713 7491 12771 7497
rect 13170 7488 13176 7500
rect 13228 7488 13234 7540
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13320 7500 13461 7528
rect 13320 7488 13326 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 18693 7531 18751 7537
rect 18693 7497 18705 7531
rect 18739 7528 18751 7531
rect 19518 7528 19524 7540
rect 18739 7500 19524 7528
rect 18739 7497 18751 7500
rect 18693 7491 18751 7497
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 8481 7463 8539 7469
rect 8481 7429 8493 7463
rect 8527 7460 8539 7463
rect 8527 7432 9996 7460
rect 8527 7429 8539 7432
rect 8481 7423 8539 7429
rect 9968 7404 9996 7432
rect 12158 7420 12164 7472
rect 12216 7460 12222 7472
rect 19061 7463 19119 7469
rect 19061 7460 19073 7463
rect 12216 7432 19073 7460
rect 12216 7420 12222 7432
rect 4448 7364 4835 7392
rect 3053 7355 3111 7361
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7324 1915 7327
rect 2498 7324 2504 7336
rect 1903 7296 2504 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 2130 7256 2136 7268
rect 2091 7228 2136 7256
rect 2130 7216 2136 7228
rect 2188 7216 2194 7268
rect 3068 7256 3096 7355
rect 3326 7333 3332 7336
rect 3320 7324 3332 7333
rect 3287 7296 3332 7324
rect 3320 7287 3332 7296
rect 3326 7284 3332 7287
rect 3384 7284 3390 7336
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 3804 7296 4629 7324
rect 3234 7256 3240 7268
rect 3068 7228 3240 7256
rect 3234 7216 3240 7228
rect 3292 7256 3298 7268
rect 3804 7256 3832 7296
rect 4617 7293 4629 7296
rect 4663 7324 4675 7327
rect 4709 7327 4767 7333
rect 4709 7324 4721 7327
rect 4663 7296 4721 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 4709 7293 4721 7296
rect 4755 7293 4767 7327
rect 4807 7324 4835 7364
rect 5810 7352 5816 7404
rect 5868 7392 5874 7404
rect 6822 7392 6828 7404
rect 5868 7364 6592 7392
rect 6783 7364 6828 7392
rect 5868 7352 5874 7364
rect 4965 7327 5023 7333
rect 4965 7324 4977 7327
rect 4807 7296 4977 7324
rect 4709 7287 4767 7293
rect 4965 7293 4977 7296
rect 5011 7324 5023 7327
rect 5718 7324 5724 7336
rect 5011 7296 5724 7324
rect 5011 7293 5023 7296
rect 4965 7287 5023 7293
rect 5718 7284 5724 7296
rect 5776 7324 5782 7336
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 5776 7296 6377 7324
rect 5776 7284 5782 7296
rect 6365 7293 6377 7296
rect 6411 7293 6423 7327
rect 6564 7324 6592 7364
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 9030 7392 9036 7404
rect 8991 7364 9036 7392
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 9950 7392 9956 7404
rect 9911 7364 9956 7392
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 10100 7364 10149 7392
rect 10100 7352 10106 7364
rect 10137 7361 10149 7364
rect 10183 7392 10195 7395
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 10183 7364 10517 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13504 7364 13829 7392
rect 13504 7352 13510 7364
rect 13817 7361 13829 7364
rect 13863 7392 13875 7395
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 13863 7364 14197 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 14185 7361 14197 7364
rect 14231 7392 14243 7395
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 14231 7364 14565 7392
rect 14231 7361 14243 7364
rect 14185 7355 14243 7361
rect 14553 7361 14565 7364
rect 14599 7392 14611 7395
rect 15010 7392 15016 7404
rect 14599 7364 15016 7392
rect 14599 7361 14611 7364
rect 14553 7355 14611 7361
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 16666 7324 16672 7336
rect 6564 7296 16672 7324
rect 6365 7287 6423 7293
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 18524 7333 18552 7432
rect 19061 7429 19073 7432
rect 19107 7429 19119 7463
rect 19061 7423 19119 7429
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 7098 7265 7104 7268
rect 7092 7256 7104 7265
rect 3292 7228 3832 7256
rect 7059 7228 7104 7256
rect 3292 7216 3298 7228
rect 7092 7219 7104 7228
rect 7098 7216 7104 7219
rect 7156 7216 7162 7268
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 10873 7259 10931 7265
rect 10873 7256 10885 7259
rect 7432 7228 10885 7256
rect 7432 7216 7438 7228
rect 10873 7225 10885 7228
rect 10919 7225 10931 7259
rect 10873 7219 10931 7225
rect 2866 7188 2872 7200
rect 2827 7160 2872 7188
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 6089 7191 6147 7197
rect 6089 7188 6101 7191
rect 5408 7160 6101 7188
rect 5408 7148 5414 7160
rect 6089 7157 6101 7160
rect 6135 7157 6147 7191
rect 6089 7151 6147 7157
rect 8205 7191 8263 7197
rect 8205 7157 8217 7191
rect 8251 7188 8263 7191
rect 8294 7188 8300 7200
rect 8251 7160 8300 7188
rect 8251 7157 8263 7160
rect 8205 7151 8263 7157
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 8846 7188 8852 7200
rect 8807 7160 8852 7188
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 8938 7148 8944 7200
rect 8996 7188 9002 7200
rect 9858 7188 9864 7200
rect 8996 7160 9041 7188
rect 9819 7160 9864 7188
rect 8996 7148 9002 7160
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 3421 6987 3479 6993
rect 3421 6953 3433 6987
rect 3467 6984 3479 6987
rect 4246 6984 4252 6996
rect 3467 6956 4252 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 5261 6987 5319 6993
rect 5261 6953 5273 6987
rect 5307 6984 5319 6987
rect 5534 6984 5540 6996
rect 5307 6956 5540 6984
rect 5307 6953 5319 6956
rect 5261 6947 5319 6953
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 5718 6984 5724 6996
rect 5679 6956 5724 6984
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 7742 6984 7748 6996
rect 7024 6956 7748 6984
rect 3326 6876 3332 6928
rect 3384 6916 3390 6928
rect 3697 6919 3755 6925
rect 3697 6916 3709 6919
rect 3384 6888 3709 6916
rect 3384 6876 3390 6888
rect 3697 6885 3709 6888
rect 3743 6885 3755 6919
rect 3697 6879 3755 6885
rect 1486 6808 1492 6860
rect 1544 6848 1550 6860
rect 1581 6851 1639 6857
rect 1581 6848 1593 6851
rect 1544 6820 1593 6848
rect 1544 6808 1550 6820
rect 1581 6817 1593 6820
rect 1627 6817 1639 6851
rect 2038 6848 2044 6860
rect 1999 6820 2044 6848
rect 1581 6811 1639 6817
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2222 6808 2228 6860
rect 2280 6848 2286 6860
rect 2501 6851 2559 6857
rect 2501 6848 2513 6851
rect 2280 6820 2513 6848
rect 2280 6808 2286 6820
rect 2501 6817 2513 6820
rect 2547 6817 2559 6851
rect 2501 6811 2559 6817
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 3050 6848 3056 6860
rect 3007 6820 3056 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 3712 6848 3740 6879
rect 4338 6876 4344 6928
rect 4396 6916 4402 6928
rect 4709 6919 4767 6925
rect 4709 6916 4721 6919
rect 4396 6888 4721 6916
rect 4396 6876 4402 6888
rect 4709 6885 4721 6888
rect 4755 6885 4767 6919
rect 4709 6879 4767 6885
rect 4801 6919 4859 6925
rect 4801 6885 4813 6919
rect 4847 6916 4859 6919
rect 5074 6916 5080 6928
rect 4847 6888 5080 6916
rect 4847 6885 4859 6888
rect 4801 6879 4859 6885
rect 5074 6876 5080 6888
rect 5132 6876 5138 6928
rect 6822 6916 6828 6928
rect 6783 6888 6828 6916
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 3712 6820 4936 6848
rect 4908 6789 4936 6820
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 6052 6820 6101 6848
rect 6052 6808 6058 6820
rect 6089 6817 6101 6820
rect 6135 6817 6147 6851
rect 6089 6811 6147 6817
rect 6733 6851 6791 6857
rect 6733 6817 6745 6851
rect 6779 6848 6791 6851
rect 7024 6848 7052 6956
rect 7742 6944 7748 6956
rect 7800 6984 7806 6996
rect 8294 6984 8300 6996
rect 7800 6956 8300 6984
rect 7800 6944 7806 6956
rect 8294 6944 8300 6956
rect 8352 6984 8358 6996
rect 10042 6984 10048 6996
rect 8352 6956 10048 6984
rect 8352 6944 8358 6956
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 7098 6876 7104 6928
rect 7156 6916 7162 6928
rect 8202 6916 8208 6928
rect 7156 6888 8208 6916
rect 7156 6876 7162 6888
rect 6779 6820 7052 6848
rect 7193 6851 7251 6857
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 7282 6848 7288 6860
rect 7239 6820 7288 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 7282 6808 7288 6820
rect 7340 6848 7346 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7340 6820 7665 6848
rect 7340 6808 7346 6820
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7760 6848 7788 6888
rect 8202 6876 8208 6888
rect 8260 6916 8266 6928
rect 8260 6888 8800 6916
rect 8260 6876 8266 6888
rect 8662 6848 8668 6860
rect 7760 6820 7880 6848
rect 8623 6820 8668 6848
rect 7653 6811 7711 6817
rect 4893 6783 4951 6789
rect 4893 6749 4905 6783
rect 4939 6780 4951 6783
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4939 6752 5273 6780
rect 4939 6749 4951 6752
rect 4893 6743 4951 6749
rect 5261 6749 5273 6752
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 7852 6789 7880 6820
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 8772 6848 8800 6888
rect 9030 6848 9036 6860
rect 8772 6820 9036 6848
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 6696 6752 7757 6780
rect 6696 6740 6702 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 4341 6715 4399 6721
rect 4341 6712 4353 6715
rect 4212 6684 4353 6712
rect 4212 6672 4218 6684
rect 4341 6681 4353 6684
rect 4387 6681 4399 6715
rect 7760 6712 7788 6743
rect 8478 6740 8484 6792
rect 8536 6780 8542 6792
rect 8864 6789 8892 6820
rect 9030 6808 9036 6820
rect 9088 6848 9094 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9088 6820 9321 6848
rect 9088 6808 9094 6820
rect 9309 6817 9321 6820
rect 9355 6848 9367 6851
rect 9398 6848 9404 6860
rect 9355 6820 9404 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9398 6808 9404 6820
rect 9456 6808 9462 6860
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 11974 6848 11980 6860
rect 10367 6820 11980 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12437 6851 12495 6857
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 12526 6848 12532 6860
rect 12483 6820 12532 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 13173 6851 13231 6857
rect 13173 6817 13185 6851
rect 13219 6848 13231 6851
rect 14182 6848 14188 6860
rect 13219 6820 14188 6848
rect 13219 6817 13231 6820
rect 13173 6811 13231 6817
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 19058 6848 19064 6860
rect 19019 6820 19064 6848
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 19613 6851 19671 6857
rect 19613 6817 19625 6851
rect 19659 6817 19671 6851
rect 19613 6811 19671 6817
rect 8757 6783 8815 6789
rect 8757 6780 8769 6783
rect 8536 6752 8769 6780
rect 8536 6740 8542 6752
rect 8757 6749 8769 6752
rect 8803 6749 8815 6783
rect 8757 6743 8815 6749
rect 8849 6783 8907 6789
rect 8849 6749 8861 6783
rect 8895 6749 8907 6783
rect 8849 6743 8907 6749
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 11848 6752 12725 6780
rect 11848 6740 11854 6752
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 19628 6724 19656 6811
rect 8110 6712 8116 6724
rect 7760 6684 8116 6712
rect 4341 6675 4399 6681
rect 8110 6672 8116 6684
rect 8168 6672 8174 6724
rect 8297 6715 8355 6721
rect 8297 6681 8309 6715
rect 8343 6712 8355 6715
rect 9858 6712 9864 6724
rect 8343 6684 9864 6712
rect 8343 6681 8355 6684
rect 8297 6675 8355 6681
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 19610 6712 19616 6724
rect 9968 6684 19616 6712
rect 5350 6644 5356 6656
rect 5311 6616 5356 6644
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7282 6644 7288 6656
rect 7243 6616 7288 6644
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7834 6604 7840 6656
rect 7892 6644 7898 6656
rect 9968 6644 9996 6684
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 19797 6715 19855 6721
rect 19797 6681 19809 6715
rect 19843 6712 19855 6715
rect 19886 6712 19892 6724
rect 19843 6684 19892 6712
rect 19843 6681 19855 6684
rect 19797 6675 19855 6681
rect 19886 6672 19892 6684
rect 19944 6672 19950 6724
rect 7892 6616 9996 6644
rect 7892 6604 7898 6616
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10597 6647 10655 6653
rect 10597 6644 10609 6647
rect 10192 6616 10609 6644
rect 10192 6604 10198 6616
rect 10597 6613 10609 6616
rect 10643 6613 10655 6647
rect 10597 6607 10655 6613
rect 10686 6604 10692 6656
rect 10744 6644 10750 6656
rect 11057 6647 11115 6653
rect 11057 6644 11069 6647
rect 10744 6616 11069 6644
rect 10744 6604 10750 6616
rect 11057 6613 11069 6616
rect 11103 6644 11115 6647
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 11103 6616 11345 6644
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 11333 6613 11345 6616
rect 11379 6613 11391 6647
rect 11333 6607 11391 6613
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11664 6616 11713 6644
rect 11664 6604 11670 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 13538 6644 13544 6656
rect 13451 6616 13544 6644
rect 11701 6607 11759 6613
rect 13538 6604 13544 6616
rect 13596 6644 13602 6656
rect 13817 6647 13875 6653
rect 13817 6644 13829 6647
rect 13596 6616 13829 6644
rect 13596 6604 13602 6616
rect 13817 6613 13829 6616
rect 13863 6613 13875 6647
rect 13817 6607 13875 6613
rect 19245 6647 19303 6653
rect 19245 6613 19257 6647
rect 19291 6644 19303 6647
rect 20070 6644 20076 6656
rect 19291 6616 20076 6644
rect 19291 6613 19303 6616
rect 19245 6607 19303 6613
rect 20070 6604 20076 6616
rect 20128 6604 20134 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 1670 6440 1676 6452
rect 1631 6412 1676 6440
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 1854 6400 1860 6452
rect 1912 6440 1918 6452
rect 2501 6443 2559 6449
rect 2501 6440 2513 6443
rect 1912 6412 2513 6440
rect 1912 6400 1918 6412
rect 2501 6409 2513 6412
rect 2547 6409 2559 6443
rect 2501 6403 2559 6409
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3513 6443 3571 6449
rect 3513 6440 3525 6443
rect 2832 6412 3525 6440
rect 2832 6400 2838 6412
rect 3513 6409 3525 6412
rect 3559 6409 3571 6443
rect 5534 6440 5540 6452
rect 5495 6412 5540 6440
rect 3513 6403 3571 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 5960 6412 6101 6440
rect 5960 6400 5966 6412
rect 6089 6409 6101 6412
rect 6135 6409 6147 6443
rect 6089 6403 6147 6409
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 6914 6440 6920 6452
rect 6687 6412 6920 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 7116 6412 7696 6440
rect 1762 6332 1768 6384
rect 1820 6372 1826 6384
rect 2133 6375 2191 6381
rect 2133 6372 2145 6375
rect 1820 6344 2145 6372
rect 1820 6332 1826 6344
rect 2133 6341 2145 6344
rect 2179 6341 2191 6375
rect 2133 6335 2191 6341
rect 3421 6375 3479 6381
rect 3421 6341 3433 6375
rect 3467 6372 3479 6375
rect 5350 6372 5356 6384
rect 3467 6344 5356 6372
rect 3467 6341 3479 6344
rect 3421 6335 3479 6341
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3970 6304 3976 6316
rect 3099 6276 3976 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4080 6313 4108 6344
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 6822 6332 6828 6384
rect 6880 6372 6886 6384
rect 7116 6381 7144 6412
rect 7101 6375 7159 6381
rect 7101 6372 7113 6375
rect 6880 6344 7113 6372
rect 6880 6332 6886 6344
rect 7101 6341 7113 6344
rect 7147 6341 7159 6375
rect 7101 6335 7159 6341
rect 7285 6375 7343 6381
rect 7285 6341 7297 6375
rect 7331 6372 7343 6375
rect 7374 6372 7380 6384
rect 7331 6344 7380 6372
rect 7331 6341 7343 6344
rect 7285 6335 7343 6341
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 7668 6245 7696 6412
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 8168 6412 8309 6440
rect 8168 6400 8174 6412
rect 8297 6409 8309 6412
rect 8343 6409 8355 6443
rect 8297 6403 8355 6409
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 8720 6412 9045 6440
rect 8720 6400 8726 6412
rect 9033 6409 9045 6412
rect 9079 6409 9091 6443
rect 9398 6440 9404 6452
rect 9359 6412 9404 6440
rect 9033 6403 9091 6409
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 9677 6443 9735 6449
rect 9677 6409 9689 6443
rect 9723 6440 9735 6443
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 9723 6412 9873 6440
rect 9723 6409 9735 6412
rect 9677 6403 9735 6409
rect 9861 6409 9873 6412
rect 9907 6440 9919 6443
rect 10229 6443 10287 6449
rect 10229 6440 10241 6443
rect 9907 6412 10241 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10229 6409 10241 6412
rect 10275 6440 10287 6443
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 10275 6412 10609 6440
rect 10275 6409 10287 6412
rect 10229 6403 10287 6409
rect 10597 6409 10609 6412
rect 10643 6440 10655 6443
rect 10686 6440 10692 6452
rect 10643 6412 10692 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 12710 6440 12716 6452
rect 12623 6412 12716 6440
rect 12710 6400 12716 6412
rect 12768 6440 12774 6452
rect 13538 6440 13544 6452
rect 12768 6412 13544 6440
rect 12768 6400 12774 6412
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 19610 6440 19616 6452
rect 19571 6412 19616 6440
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 20073 6443 20131 6449
rect 20073 6409 20085 6443
rect 20119 6440 20131 6443
rect 20714 6440 20720 6452
rect 20119 6412 20720 6440
rect 20119 6409 20131 6412
rect 20073 6403 20131 6409
rect 20714 6400 20720 6412
rect 20772 6400 20778 6452
rect 7926 6332 7932 6384
rect 7984 6372 7990 6384
rect 10134 6372 10140 6384
rect 7984 6344 10140 6372
rect 7984 6332 7990 6344
rect 10134 6332 10140 6344
rect 10192 6332 10198 6384
rect 11333 6375 11391 6381
rect 11333 6341 11345 6375
rect 11379 6372 11391 6375
rect 11793 6375 11851 6381
rect 11793 6372 11805 6375
rect 11379 6344 11805 6372
rect 11379 6341 11391 6344
rect 11333 6335 11391 6341
rect 11793 6341 11805 6344
rect 11839 6372 11851 6375
rect 12161 6375 12219 6381
rect 12161 6372 12173 6375
rect 11839 6344 12173 6372
rect 11839 6341 11851 6344
rect 11793 6335 11851 6341
rect 12161 6341 12173 6344
rect 12207 6372 12219 6375
rect 13446 6372 13452 6384
rect 12207 6344 13452 6372
rect 12207 6341 12219 6344
rect 12161 6335 12219 6341
rect 13446 6332 13452 6344
rect 13504 6332 13510 6384
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7800 6276 7849 6304
rect 7800 6264 7806 6276
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 8444 6276 9689 6304
rect 8444 6264 8450 6276
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 3881 6239 3939 6245
rect 3881 6236 3893 6239
rect 3016 6208 3893 6236
rect 3016 6196 3022 6208
rect 3881 6205 3893 6208
rect 3927 6205 3939 6239
rect 3881 6199 3939 6205
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6205 7711 6239
rect 7653 6199 7711 6205
rect 9306 6196 9312 6248
rect 9364 6236 9370 6248
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 9364 6208 10885 6236
rect 9364 6196 9370 6208
rect 10873 6205 10885 6208
rect 10919 6236 10931 6239
rect 11606 6236 11612 6248
rect 10919 6208 11612 6236
rect 10919 6205 10931 6208
rect 10873 6199 10931 6205
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 12158 6196 12164 6248
rect 12216 6236 12222 6248
rect 19889 6239 19947 6245
rect 19889 6236 19901 6239
rect 12216 6208 19901 6236
rect 12216 6196 12222 6208
rect 19889 6205 19901 6208
rect 19935 6236 19947 6239
rect 20441 6239 20499 6245
rect 20441 6236 20453 6239
rect 19935 6208 20453 6236
rect 19935 6205 19947 6208
rect 19889 6199 19947 6205
rect 20441 6205 20453 6208
rect 20487 6205 20499 6239
rect 20441 6199 20499 6205
rect 6454 6128 6460 6180
rect 6512 6168 6518 6180
rect 8478 6168 8484 6180
rect 6512 6140 8484 6168
rect 6512 6128 6518 6140
rect 8478 6128 8484 6140
rect 8536 6168 8542 6180
rect 8665 6171 8723 6177
rect 8665 6168 8677 6171
rect 8536 6140 8677 6168
rect 8536 6128 8542 6140
rect 8665 6137 8677 6140
rect 8711 6137 8723 6171
rect 8665 6131 8723 6137
rect 4246 6060 4252 6112
rect 4304 6100 4310 6112
rect 4709 6103 4767 6109
rect 4709 6100 4721 6103
rect 4304 6072 4721 6100
rect 4304 6060 4310 6072
rect 4709 6069 4721 6072
rect 4755 6069 4767 6103
rect 5074 6100 5080 6112
rect 5035 6072 5080 6100
rect 4709 6063 4767 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 7432 6072 7757 6100
rect 7432 6060 7438 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 19058 6100 19064 6112
rect 8352 6072 19064 6100
rect 8352 6060 8358 6072
rect 19058 6060 19064 6072
rect 19116 6060 19122 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 2832 5868 2877 5896
rect 2832 5856 2838 5868
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3016 5868 3433 5896
rect 3016 5856 3022 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 3421 5859 3479 5865
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 4154 5896 4160 5908
rect 3927 5868 4160 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 4154 5856 4160 5868
rect 4212 5856 4218 5908
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 5169 5899 5227 5905
rect 5169 5896 5181 5899
rect 4856 5868 5181 5896
rect 4856 5856 4862 5868
rect 5169 5865 5181 5868
rect 5215 5865 5227 5899
rect 5626 5896 5632 5908
rect 5587 5868 5632 5896
rect 5169 5859 5227 5865
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 6178 5896 6184 5908
rect 6139 5868 6184 5896
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 6546 5896 6552 5908
rect 6507 5868 6552 5896
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7282 5896 7288 5908
rect 7243 5868 7288 5896
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 8113 5899 8171 5905
rect 8113 5865 8125 5899
rect 8159 5896 8171 5899
rect 8202 5896 8208 5908
rect 8159 5868 8208 5896
rect 8159 5865 8171 5868
rect 8113 5859 8171 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8754 5896 8760 5908
rect 8715 5868 8760 5896
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 10594 5856 10600 5908
rect 10652 5896 10658 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10652 5868 10701 5896
rect 10652 5856 10658 5868
rect 10689 5865 10701 5868
rect 10735 5896 10747 5899
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 10735 5868 11069 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 11057 5865 11069 5868
rect 11103 5896 11115 5899
rect 11425 5899 11483 5905
rect 11425 5896 11437 5899
rect 11103 5868 11437 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 11425 5865 11437 5868
rect 11471 5896 11483 5899
rect 12710 5896 12716 5908
rect 11471 5868 12716 5896
rect 11471 5865 11483 5868
rect 11425 5859 11483 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 20441 5899 20499 5905
rect 20441 5865 20453 5899
rect 20487 5896 20499 5899
rect 21174 5896 21180 5908
rect 20487 5868 21180 5896
rect 20487 5865 20499 5868
rect 20441 5859 20499 5865
rect 21174 5856 21180 5868
rect 21232 5856 21238 5908
rect 1394 5788 1400 5840
rect 1452 5828 1458 5840
rect 1949 5831 2007 5837
rect 1949 5828 1961 5831
rect 1452 5800 1961 5828
rect 1452 5788 1458 5800
rect 1949 5797 1961 5800
rect 1995 5797 2007 5831
rect 1949 5791 2007 5797
rect 3145 5831 3203 5837
rect 3145 5797 3157 5831
rect 3191 5828 3203 5831
rect 3602 5828 3608 5840
rect 3191 5800 3608 5828
rect 3191 5797 3203 5800
rect 3145 5791 3203 5797
rect 3602 5788 3608 5800
rect 3660 5788 3666 5840
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 12158 5828 12164 5840
rect 4120 5800 12164 5828
rect 4120 5788 4126 5800
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 5258 5760 5264 5772
rect 4387 5732 5264 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 7190 5760 7196 5772
rect 7055 5732 7196 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 7800 5732 8401 5760
rect 7800 5720 7806 5732
rect 8389 5729 8401 5732
rect 8435 5729 8447 5763
rect 20254 5760 20260 5772
rect 20215 5732 20260 5760
rect 8389 5723 8447 5729
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 4890 5692 4896 5704
rect 4851 5664 4896 5692
rect 4890 5652 4896 5664
rect 4948 5652 4954 5704
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 7616 5664 9137 5692
rect 7616 5652 7622 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 4798 5584 4804 5636
rect 4856 5624 4862 5636
rect 5166 5624 5172 5636
rect 4856 5596 5172 5624
rect 4856 5584 4862 5596
rect 5166 5584 5172 5596
rect 5224 5624 5230 5636
rect 8662 5624 8668 5636
rect 5224 5596 8668 5624
rect 5224 5584 5230 5596
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 5350 5516 5356 5568
rect 5408 5556 5414 5568
rect 7098 5556 7104 5568
rect 5408 5528 7104 5556
rect 5408 5516 5414 5528
rect 7098 5516 7104 5528
rect 7156 5556 7162 5568
rect 7653 5559 7711 5565
rect 7653 5556 7665 5559
rect 7156 5528 7665 5556
rect 7156 5516 7162 5528
rect 7653 5525 7665 5528
rect 7699 5525 7711 5559
rect 7653 5519 7711 5525
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 9364 5528 9873 5556
rect 9364 5516 9370 5528
rect 9861 5525 9873 5528
rect 9907 5556 9919 5559
rect 10229 5559 10287 5565
rect 10229 5556 10241 5559
rect 9907 5528 10241 5556
rect 9907 5525 9919 5528
rect 9861 5519 9919 5525
rect 10229 5525 10241 5528
rect 10275 5525 10287 5559
rect 10229 5519 10287 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 2225 5355 2283 5361
rect 2225 5321 2237 5355
rect 2271 5352 2283 5355
rect 2406 5352 2412 5364
rect 2271 5324 2412 5352
rect 2271 5321 2283 5324
rect 2225 5315 2283 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 2590 5352 2596 5364
rect 2551 5324 2596 5352
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 2961 5355 3019 5361
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 3418 5352 3424 5364
rect 3007 5324 3424 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4706 5352 4712 5364
rect 4571 5324 4712 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6086 5352 6092 5364
rect 6043 5324 6092 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7466 5352 7472 5364
rect 7147 5324 7472 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7466 5312 7472 5324
rect 7524 5312 7530 5364
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 7929 5355 7987 5361
rect 7929 5352 7941 5355
rect 7800 5324 7941 5352
rect 7800 5312 7806 5324
rect 7929 5321 7941 5324
rect 7975 5352 7987 5355
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 7975 5324 8309 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8297 5321 8309 5324
rect 8343 5352 8355 5355
rect 8386 5352 8392 5364
rect 8343 5324 8392 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 8570 5352 8576 5364
rect 8531 5324 8576 5352
rect 8570 5312 8576 5324
rect 8628 5352 8634 5364
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 8628 5324 8953 5352
rect 8628 5312 8634 5324
rect 8941 5321 8953 5324
rect 8987 5352 8999 5355
rect 9306 5352 9312 5364
rect 8987 5324 9312 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 20717 5355 20775 5361
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 20898 5352 20904 5364
rect 20763 5324 20904 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 3329 5287 3387 5293
rect 3329 5253 3341 5287
rect 3375 5284 3387 5287
rect 3694 5284 3700 5296
rect 3375 5256 3700 5284
rect 3375 5253 3387 5256
rect 3329 5247 3387 5253
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 6365 5287 6423 5293
rect 6365 5253 6377 5287
rect 6411 5284 6423 5287
rect 7558 5284 7564 5296
rect 6411 5256 7564 5284
rect 6411 5253 6423 5256
rect 6365 5247 6423 5253
rect 7558 5244 7564 5256
rect 7616 5244 7622 5296
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 3142 5216 3148 5228
rect 1719 5188 3148 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 3292 5188 3617 5216
rect 3292 5176 3298 5188
rect 3605 5185 3617 5188
rect 3651 5216 3663 5219
rect 4157 5219 4215 5225
rect 4157 5216 4169 5219
rect 3651 5188 4169 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 4157 5185 4169 5188
rect 4203 5216 4215 5219
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4203 5188 4813 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 4801 5185 4813 5188
rect 4847 5216 4859 5219
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4847 5188 5181 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 5169 5185 5181 5188
rect 5215 5216 5227 5219
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 5215 5188 5549 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5537 5185 5549 5188
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 7650 5216 7656 5228
rect 7515 5188 7656 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 4120 5120 20545 5148
rect 4120 5108 4126 5120
rect 20533 5117 20545 5120
rect 20579 5148 20591 5151
rect 21085 5151 21143 5157
rect 21085 5148 21097 5151
rect 20579 5120 21097 5148
rect 20579 5117 20591 5120
rect 20533 5111 20591 5117
rect 21085 5117 21097 5120
rect 21131 5117 21143 5151
rect 21085 5111 21143 5117
rect 3970 5040 3976 5092
rect 4028 5080 4034 5092
rect 20254 5080 20260 5092
rect 4028 5052 20260 5080
rect 4028 5040 4034 5052
rect 20254 5040 20260 5052
rect 20312 5040 20318 5092
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 2130 4808 2136 4820
rect 1903 4780 2136 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 2225 4811 2283 4817
rect 2225 4777 2237 4811
rect 2271 4808 2283 4811
rect 2498 4808 2504 4820
rect 2271 4780 2504 4808
rect 2271 4777 2283 4780
rect 2225 4771 2283 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 2593 4811 2651 4817
rect 2593 4777 2605 4811
rect 2639 4808 2651 4811
rect 2682 4808 2688 4820
rect 2639 4780 2688 4808
rect 2639 4777 2651 4780
rect 2593 4771 2651 4777
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 2961 4811 3019 4817
rect 2961 4777 2973 4811
rect 3007 4808 3019 4811
rect 3234 4808 3240 4820
rect 3007 4780 3240 4808
rect 3007 4777 3019 4780
rect 2961 4771 3019 4777
rect 3234 4768 3240 4780
rect 3292 4808 3298 4820
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 3292 4780 4905 4808
rect 3292 4768 3298 4780
rect 4893 4777 4905 4780
rect 4939 4808 4951 4811
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 4939 4780 5273 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 5261 4777 5273 4780
rect 5307 4808 5319 4811
rect 5629 4811 5687 4817
rect 5629 4808 5641 4811
rect 5307 4780 5641 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5629 4777 5641 4780
rect 5675 4777 5687 4811
rect 5629 4771 5687 4777
rect 6549 4811 6607 4817
rect 6549 4777 6561 4811
rect 6595 4808 6607 4811
rect 6730 4808 6736 4820
rect 6595 4780 6736 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 6917 4811 6975 4817
rect 6917 4777 6929 4811
rect 6963 4808 6975 4811
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 6963 4780 7297 4808
rect 6963 4777 6975 4780
rect 6917 4771 6975 4777
rect 7285 4777 7297 4780
rect 7331 4808 7343 4811
rect 7653 4811 7711 4817
rect 7653 4808 7665 4811
rect 7331 4780 7665 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 7653 4777 7665 4780
rect 7699 4808 7711 4811
rect 7742 4808 7748 4820
rect 7699 4780 7748 4808
rect 7699 4777 7711 4780
rect 7653 4771 7711 4777
rect 6089 4743 6147 4749
rect 6089 4709 6101 4743
rect 6135 4740 6147 4743
rect 6932 4740 6960 4771
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 8021 4811 8079 4817
rect 8021 4777 8033 4811
rect 8067 4808 8079 4811
rect 8570 4808 8576 4820
rect 8067 4780 8576 4808
rect 8067 4777 8079 4780
rect 8021 4771 8079 4777
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 6135 4712 6960 4740
rect 6135 4709 6147 4712
rect 6089 4703 6147 4709
rect 3697 4471 3755 4477
rect 3697 4437 3709 4471
rect 3743 4468 3755 4471
rect 4062 4468 4068 4480
rect 3743 4440 4068 4468
rect 3743 4437 3755 4440
rect 3697 4431 3755 4437
rect 4062 4428 4068 4440
rect 4120 4468 4126 4480
rect 4525 4471 4583 4477
rect 4525 4468 4537 4471
rect 4120 4440 4537 4468
rect 4120 4428 4126 4440
rect 4525 4437 4537 4440
rect 4571 4437 4583 4471
rect 4525 4431 4583 4437
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 7469 4267 7527 4273
rect 7469 4233 7481 4267
rect 7515 4264 7527 4267
rect 7837 4267 7895 4273
rect 7837 4264 7849 4267
rect 7515 4236 7849 4264
rect 7515 4233 7527 4236
rect 7469 4227 7527 4233
rect 7837 4233 7849 4236
rect 7883 4264 7895 4267
rect 8570 4264 8576 4276
rect 7883 4236 8576 4264
rect 7883 4233 7895 4236
rect 7837 4227 7895 4233
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 2777 4199 2835 4205
rect 2777 4165 2789 4199
rect 2823 4196 2835 4199
rect 2958 4196 2964 4208
rect 2823 4168 2964 4196
rect 2823 4165 2835 4168
rect 2777 4159 2835 4165
rect 2958 4156 2964 4168
rect 3016 4196 3022 4208
rect 3145 4199 3203 4205
rect 3145 4196 3157 4199
rect 3016 4168 3157 4196
rect 3016 4156 3022 4168
rect 3145 4165 3157 4168
rect 3191 4196 3203 4199
rect 3191 4168 3556 4196
rect 3191 4165 3203 4168
rect 3145 4159 3203 4165
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1452 4100 1593 4128
rect 1452 4088 1458 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 3234 4128 3240 4140
rect 2363 4100 3240 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3528 4137 3556 4168
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3559 4100 3985 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3973 4097 3985 4100
rect 4019 4128 4031 4131
rect 4062 4128 4068 4140
rect 4019 4100 4068 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 4062 4088 4068 4100
rect 4120 4128 4126 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4120 4100 4997 4128
rect 4120 4088 4126 4100
rect 4985 4097 4997 4100
rect 5031 4128 5043 4131
rect 5353 4131 5411 4137
rect 5353 4128 5365 4131
rect 5031 4100 5365 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5353 4097 5365 4100
rect 5399 4128 5411 4131
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5399 4100 5733 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 5721 4097 5733 4100
rect 5767 4128 5779 4131
rect 6730 4128 6736 4140
rect 5767 4100 6736 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 6730 4088 6736 4100
rect 6788 4128 6794 4140
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6788 4100 7021 4128
rect 6788 4088 6794 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 11146 4060 11152 4072
rect 5500 4032 11152 4060
rect 5500 4020 5506 4032
rect 11146 4020 11152 4032
rect 11204 4020 11210 4072
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 5350 3992 5356 4004
rect 4028 3964 5356 3992
rect 4028 3952 4034 3964
rect 5350 3952 5356 3964
rect 5408 3952 5414 4004
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 2958 3720 2964 3732
rect 2919 3692 2964 3720
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 5077 3723 5135 3729
rect 5077 3720 5089 3723
rect 4120 3692 5089 3720
rect 4120 3680 4126 3692
rect 5077 3689 5089 3692
rect 5123 3689 5135 3723
rect 5077 3683 5135 3689
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
<< via1 >>
rect 4068 20340 4120 20392
rect 20076 20340 20128 20392
rect 8208 20272 8260 20324
rect 15292 20272 15344 20324
rect 7196 20204 7248 20256
rect 15108 20204 15160 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 1676 20043 1728 20052
rect 1676 20009 1685 20043
rect 1685 20009 1719 20043
rect 1719 20009 1728 20043
rect 1676 20000 1728 20009
rect 2320 19932 2372 19984
rect 5632 20000 5684 20052
rect 8392 20043 8444 20052
rect 8392 20009 8401 20043
rect 8401 20009 8435 20043
rect 8435 20009 8444 20043
rect 8392 20000 8444 20009
rect 8852 20000 8904 20052
rect 9312 20043 9364 20052
rect 9312 20009 9321 20043
rect 9321 20009 9355 20043
rect 9355 20009 9364 20043
rect 9312 20000 9364 20009
rect 9680 20000 9732 20052
rect 13360 20000 13412 20052
rect 14280 20000 14332 20052
rect 15108 20043 15160 20052
rect 15108 20009 15117 20043
rect 15117 20009 15151 20043
rect 15151 20009 15160 20043
rect 15108 20000 15160 20009
rect 15292 20000 15344 20052
rect 16580 20000 16632 20052
rect 17040 20000 17092 20052
rect 17960 20000 18012 20052
rect 20076 20043 20128 20052
rect 20076 20009 20085 20043
rect 20085 20009 20119 20043
rect 20119 20009 20128 20043
rect 20076 20000 20128 20009
rect 2872 19864 2924 19916
rect 4068 19864 4120 19916
rect 4252 19864 4304 19916
rect 1400 19796 1452 19848
rect 4988 19796 5040 19848
rect 4896 19728 4948 19780
rect 11060 19932 11112 19984
rect 9680 19864 9732 19916
rect 9128 19796 9180 19848
rect 12624 19796 12676 19848
rect 13360 19864 13412 19916
rect 14464 19864 14516 19916
rect 15108 19864 15160 19916
rect 16580 19864 16632 19916
rect 17316 19932 17368 19984
rect 18696 19864 18748 19916
rect 18972 19864 19024 19916
rect 9864 19728 9916 19780
rect 18420 19728 18472 19780
rect 3608 19660 3660 19712
rect 4068 19703 4120 19712
rect 4068 19669 4077 19703
rect 4077 19669 4111 19703
rect 4111 19669 4120 19703
rect 4068 19660 4120 19669
rect 6736 19703 6788 19712
rect 6736 19669 6745 19703
rect 6745 19669 6779 19703
rect 6779 19669 6788 19703
rect 6736 19660 6788 19669
rect 7104 19703 7156 19712
rect 7104 19669 7113 19703
rect 7113 19669 7147 19703
rect 7147 19669 7156 19703
rect 7104 19660 7156 19669
rect 7288 19660 7340 19712
rect 8576 19660 8628 19712
rect 8760 19703 8812 19712
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 9404 19660 9456 19712
rect 10140 19660 10192 19712
rect 10416 19660 10468 19712
rect 11796 19660 11848 19712
rect 12624 19660 12676 19712
rect 14372 19703 14424 19712
rect 14372 19669 14381 19703
rect 14381 19669 14415 19703
rect 14415 19669 14424 19703
rect 14372 19660 14424 19669
rect 16672 19703 16724 19712
rect 16672 19669 16681 19703
rect 16681 19669 16715 19703
rect 16715 19669 16724 19703
rect 16672 19660 16724 19669
rect 17040 19703 17092 19712
rect 17040 19669 17049 19703
rect 17049 19669 17083 19703
rect 17083 19669 17092 19703
rect 17040 19660 17092 19669
rect 19800 19703 19852 19712
rect 19800 19669 19809 19703
rect 19809 19669 19843 19703
rect 19843 19669 19852 19703
rect 19800 19660 19852 19669
rect 20444 19703 20496 19712
rect 20444 19669 20453 19703
rect 20453 19669 20487 19703
rect 20487 19669 20496 19703
rect 20444 19660 20496 19669
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 2228 19456 2280 19508
rect 17040 19456 17092 19508
rect 9680 19388 9732 19440
rect 19064 19456 19116 19508
rect 2228 19320 2280 19372
rect 4896 19320 4948 19372
rect 8392 19363 8444 19372
rect 2320 19227 2372 19236
rect 2320 19193 2329 19227
rect 2329 19193 2363 19227
rect 2363 19193 2372 19227
rect 2320 19184 2372 19193
rect 2596 19252 2648 19304
rect 4068 19252 4120 19304
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 8392 19329 8401 19363
rect 8401 19329 8435 19363
rect 8435 19329 8444 19363
rect 8392 19320 8444 19329
rect 6736 19184 6788 19236
rect 7656 19252 7708 19304
rect 9312 19320 9364 19372
rect 9864 19320 9916 19372
rect 9312 19227 9364 19236
rect 9312 19193 9321 19227
rect 9321 19193 9355 19227
rect 9355 19193 9364 19227
rect 9312 19184 9364 19193
rect 1584 19116 1636 19168
rect 2136 19116 2188 19168
rect 4528 19116 4580 19168
rect 4896 19159 4948 19168
rect 4896 19125 4905 19159
rect 4905 19125 4939 19159
rect 4939 19125 4948 19159
rect 4896 19116 4948 19125
rect 4988 19116 5040 19168
rect 6644 19116 6696 19168
rect 8208 19116 8260 19168
rect 8760 19116 8812 19168
rect 8944 19159 8996 19168
rect 8944 19125 8953 19159
rect 8953 19125 8987 19159
rect 8987 19125 8996 19159
rect 8944 19116 8996 19125
rect 9496 19252 9548 19304
rect 11152 19252 11204 19304
rect 12072 19252 12124 19304
rect 12992 19252 13044 19304
rect 13636 19295 13688 19304
rect 13636 19261 13645 19295
rect 13645 19261 13679 19295
rect 13679 19261 13688 19295
rect 13636 19252 13688 19261
rect 14004 19252 14056 19304
rect 14096 19252 14148 19304
rect 14280 19252 14332 19304
rect 15844 19295 15896 19304
rect 9680 19184 9732 19236
rect 10140 19184 10192 19236
rect 11888 19227 11940 19236
rect 11888 19193 11897 19227
rect 11897 19193 11931 19227
rect 11931 19193 11940 19227
rect 11888 19184 11940 19193
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 16396 19295 16448 19304
rect 16396 19261 16405 19295
rect 16405 19261 16439 19295
rect 16439 19261 16448 19295
rect 16396 19252 16448 19261
rect 18696 19388 18748 19440
rect 17592 19252 17644 19304
rect 17776 19252 17828 19304
rect 18144 19252 18196 19304
rect 19800 19295 19852 19304
rect 17500 19184 17552 19236
rect 12900 19116 12952 19168
rect 13912 19116 13964 19168
rect 15016 19116 15068 19168
rect 15200 19116 15252 19168
rect 15660 19116 15712 19168
rect 16120 19116 16172 19168
rect 17684 19159 17736 19168
rect 17684 19125 17693 19159
rect 17693 19125 17727 19159
rect 17727 19125 17736 19159
rect 17684 19116 17736 19125
rect 18328 19227 18380 19236
rect 18328 19193 18337 19227
rect 18337 19193 18371 19227
rect 18371 19193 18380 19227
rect 18328 19184 18380 19193
rect 19800 19261 19809 19295
rect 19809 19261 19843 19295
rect 19843 19261 19852 19295
rect 19800 19252 19852 19261
rect 22100 19252 22152 19304
rect 19340 19227 19392 19236
rect 19340 19193 19349 19227
rect 19349 19193 19383 19227
rect 19383 19193 19392 19227
rect 19340 19184 19392 19193
rect 19616 19184 19668 19236
rect 20812 19116 20864 19168
rect 20904 19159 20956 19168
rect 20904 19125 20913 19159
rect 20913 19125 20947 19159
rect 20947 19125 20956 19159
rect 20904 19116 20956 19125
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 2780 18912 2832 18964
rect 2872 18955 2924 18964
rect 2872 18921 2881 18955
rect 2881 18921 2915 18955
rect 2915 18921 2924 18955
rect 2872 18912 2924 18921
rect 5172 18912 5224 18964
rect 6736 18955 6788 18964
rect 6736 18921 6745 18955
rect 6745 18921 6779 18955
rect 6779 18921 6788 18955
rect 6736 18912 6788 18921
rect 2228 18887 2280 18896
rect 2228 18853 2237 18887
rect 2237 18853 2271 18887
rect 2271 18853 2280 18887
rect 2228 18844 2280 18853
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 2688 18776 2740 18828
rect 204 18708 256 18760
rect 3056 18708 3108 18760
rect 1492 18572 1544 18624
rect 2688 18572 2740 18624
rect 3240 18572 3292 18624
rect 5080 18776 5132 18828
rect 5632 18819 5684 18828
rect 5632 18785 5666 18819
rect 5666 18785 5684 18819
rect 5632 18776 5684 18785
rect 5816 18844 5868 18896
rect 10324 18912 10376 18964
rect 7656 18776 7708 18828
rect 8024 18844 8076 18896
rect 8760 18844 8812 18896
rect 9312 18887 9364 18896
rect 9312 18853 9321 18887
rect 9321 18853 9355 18887
rect 9355 18853 9364 18887
rect 9312 18844 9364 18853
rect 9864 18844 9916 18896
rect 10968 18844 11020 18896
rect 10508 18776 10560 18828
rect 11612 18776 11664 18828
rect 13636 18912 13688 18964
rect 12164 18776 12216 18828
rect 12900 18776 12952 18828
rect 13268 18819 13320 18828
rect 13268 18785 13277 18819
rect 13277 18785 13311 18819
rect 13311 18785 13320 18819
rect 13268 18776 13320 18785
rect 14004 18844 14056 18896
rect 14280 18844 14332 18896
rect 15844 18844 15896 18896
rect 14096 18776 14148 18828
rect 15476 18776 15528 18828
rect 16488 18776 16540 18828
rect 16764 18819 16816 18828
rect 16764 18785 16773 18819
rect 16773 18785 16807 18819
rect 16807 18785 16816 18819
rect 16764 18776 16816 18785
rect 17868 18776 17920 18828
rect 18144 18776 18196 18828
rect 18420 18819 18472 18828
rect 18420 18785 18429 18819
rect 18429 18785 18463 18819
rect 18463 18785 18472 18819
rect 18420 18776 18472 18785
rect 4528 18708 4580 18760
rect 4804 18708 4856 18760
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 7380 18708 7432 18760
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 9588 18708 9640 18760
rect 13360 18708 13412 18760
rect 16120 18708 16172 18760
rect 4068 18683 4120 18692
rect 4068 18649 4077 18683
rect 4077 18649 4111 18683
rect 4111 18649 4120 18683
rect 4068 18640 4120 18649
rect 10876 18640 10928 18692
rect 16396 18708 16448 18760
rect 16580 18708 16632 18760
rect 18972 18708 19024 18760
rect 19156 18751 19208 18760
rect 19156 18717 19165 18751
rect 19165 18717 19199 18751
rect 19199 18717 19208 18751
rect 19156 18708 19208 18717
rect 3976 18572 4028 18624
rect 5724 18572 5776 18624
rect 8208 18572 8260 18624
rect 9680 18572 9732 18624
rect 14004 18615 14056 18624
rect 14004 18581 14013 18615
rect 14013 18581 14047 18615
rect 14047 18581 14056 18615
rect 14004 18572 14056 18581
rect 15016 18572 15068 18624
rect 15568 18572 15620 18624
rect 20444 18640 20496 18692
rect 16672 18572 16724 18624
rect 16856 18572 16908 18624
rect 17592 18572 17644 18624
rect 19984 18572 20036 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 3056 18368 3108 18420
rect 3976 18368 4028 18420
rect 5172 18368 5224 18420
rect 6276 18368 6328 18420
rect 10876 18368 10928 18420
rect 10968 18368 11020 18420
rect 13728 18368 13780 18420
rect 15384 18368 15436 18420
rect 2688 18300 2740 18352
rect 3700 18300 3752 18352
rect 1952 18232 2004 18284
rect 2228 18232 2280 18284
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 2688 18207 2740 18216
rect 2688 18173 2697 18207
rect 2697 18173 2731 18207
rect 2731 18173 2740 18207
rect 2688 18164 2740 18173
rect 4252 18232 4304 18284
rect 5080 18300 5132 18352
rect 5448 18232 5500 18284
rect 5908 18232 5960 18284
rect 6644 18232 6696 18284
rect 5540 18164 5592 18216
rect 8484 18300 8536 18352
rect 9404 18300 9456 18352
rect 10784 18300 10836 18352
rect 12348 18300 12400 18352
rect 8024 18232 8076 18284
rect 8208 18275 8260 18284
rect 8208 18241 8217 18275
rect 8217 18241 8251 18275
rect 8251 18241 8260 18275
rect 8208 18232 8260 18241
rect 8392 18232 8444 18284
rect 9680 18232 9732 18284
rect 10876 18232 10928 18284
rect 13820 18300 13872 18352
rect 15016 18300 15068 18352
rect 18880 18368 18932 18420
rect 19432 18411 19484 18420
rect 19432 18377 19441 18411
rect 19441 18377 19475 18411
rect 19475 18377 19484 18411
rect 19432 18368 19484 18377
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 4068 18096 4120 18148
rect 4252 18028 4304 18080
rect 4804 18028 4856 18080
rect 5172 18028 5224 18080
rect 5356 18028 5408 18080
rect 5816 18028 5868 18080
rect 6092 18096 6144 18148
rect 7196 18096 7248 18148
rect 7380 18096 7432 18148
rect 8116 18096 8168 18148
rect 9128 18207 9180 18216
rect 9128 18173 9137 18207
rect 9137 18173 9171 18207
rect 9171 18173 9180 18207
rect 9128 18164 9180 18173
rect 9588 18164 9640 18216
rect 8944 18096 8996 18148
rect 14372 18164 14424 18216
rect 15384 18232 15436 18284
rect 15568 18232 15620 18284
rect 18788 18300 18840 18352
rect 14556 18164 14608 18216
rect 16028 18164 16080 18216
rect 16120 18164 16172 18216
rect 17408 18232 17460 18284
rect 7564 18028 7616 18080
rect 9588 18028 9640 18080
rect 9680 18028 9732 18080
rect 10876 18028 10928 18080
rect 10968 18028 11020 18080
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 12900 18028 12952 18080
rect 13728 18028 13780 18080
rect 13912 18071 13964 18080
rect 13912 18037 13921 18071
rect 13921 18037 13955 18071
rect 13955 18037 13964 18071
rect 14464 18071 14516 18080
rect 13912 18028 13964 18037
rect 14464 18037 14473 18071
rect 14473 18037 14507 18071
rect 14507 18037 14516 18071
rect 14464 18028 14516 18037
rect 15108 18028 15160 18080
rect 15292 18096 15344 18148
rect 16488 18139 16540 18148
rect 16488 18105 16497 18139
rect 16497 18105 16531 18139
rect 16531 18105 16540 18139
rect 16488 18096 16540 18105
rect 15384 18071 15436 18080
rect 15384 18037 15393 18071
rect 15393 18037 15427 18071
rect 15427 18037 15436 18071
rect 15384 18028 15436 18037
rect 16028 18071 16080 18080
rect 16028 18037 16037 18071
rect 16037 18037 16071 18071
rect 16071 18037 16080 18071
rect 16028 18028 16080 18037
rect 16120 18028 16172 18080
rect 18512 18164 18564 18216
rect 18788 18164 18840 18216
rect 19064 18207 19116 18216
rect 19064 18173 19073 18207
rect 19073 18173 19107 18207
rect 19107 18173 19116 18207
rect 19064 18164 19116 18173
rect 19984 18164 20036 18216
rect 20904 18164 20956 18216
rect 21640 18164 21692 18216
rect 17316 18096 17368 18148
rect 19708 18096 19760 18148
rect 19892 18096 19944 18148
rect 20260 18096 20312 18148
rect 19248 18028 19300 18080
rect 19984 18028 20036 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 2780 17824 2832 17876
rect 3056 17824 3108 17876
rect 4252 17867 4304 17876
rect 4252 17833 4261 17867
rect 4261 17833 4295 17867
rect 4295 17833 4304 17867
rect 4252 17824 4304 17833
rect 5632 17824 5684 17876
rect 7564 17824 7616 17876
rect 8208 17824 8260 17876
rect 8392 17867 8444 17876
rect 8392 17833 8401 17867
rect 8401 17833 8435 17867
rect 8435 17833 8444 17867
rect 8392 17824 8444 17833
rect 9128 17824 9180 17876
rect 9312 17824 9364 17876
rect 9680 17824 9732 17876
rect 9772 17824 9824 17876
rect 11152 17824 11204 17876
rect 12716 17824 12768 17876
rect 12808 17824 12860 17876
rect 13912 17824 13964 17876
rect 2872 17731 2924 17740
rect 1032 17620 1084 17672
rect 2872 17697 2881 17731
rect 2881 17697 2915 17731
rect 2915 17697 2924 17731
rect 2872 17688 2924 17697
rect 6092 17756 6144 17808
rect 14464 17756 14516 17808
rect 16948 17756 17000 17808
rect 20444 17756 20496 17808
rect 1492 17552 1544 17604
rect 2780 17620 2832 17672
rect 4252 17620 4304 17672
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 5172 17620 5224 17672
rect 7656 17688 7708 17740
rect 8484 17731 8536 17740
rect 8484 17697 8493 17731
rect 8493 17697 8527 17731
rect 8527 17697 8536 17731
rect 8484 17688 8536 17697
rect 8668 17688 8720 17740
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 11704 17688 11756 17740
rect 11888 17688 11940 17740
rect 13820 17688 13872 17740
rect 14556 17731 14608 17740
rect 14556 17697 14565 17731
rect 14565 17697 14599 17731
rect 14599 17697 14608 17731
rect 14556 17688 14608 17697
rect 15108 17688 15160 17740
rect 15568 17731 15620 17740
rect 15568 17697 15602 17731
rect 15602 17697 15620 17731
rect 15568 17688 15620 17697
rect 16764 17688 16816 17740
rect 17684 17688 17736 17740
rect 10600 17620 10652 17672
rect 11796 17620 11848 17672
rect 12992 17620 13044 17672
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 3332 17552 3384 17604
rect 6276 17552 6328 17604
rect 4068 17484 4120 17536
rect 6000 17484 6052 17536
rect 6644 17527 6696 17536
rect 6644 17493 6653 17527
rect 6653 17493 6687 17527
rect 6687 17493 6696 17527
rect 6644 17484 6696 17493
rect 7288 17552 7340 17604
rect 9312 17552 9364 17604
rect 10416 17552 10468 17604
rect 13360 17595 13412 17604
rect 11704 17484 11756 17536
rect 11888 17527 11940 17536
rect 11888 17493 11897 17527
rect 11897 17493 11931 17527
rect 11931 17493 11940 17527
rect 11888 17484 11940 17493
rect 13360 17561 13369 17595
rect 13369 17561 13403 17595
rect 13403 17561 13412 17595
rect 13360 17552 13412 17561
rect 14004 17552 14056 17604
rect 15016 17620 15068 17672
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 16488 17620 16540 17672
rect 17316 17620 17368 17672
rect 17868 17620 17920 17672
rect 19064 17688 19116 17740
rect 15200 17552 15252 17604
rect 17408 17595 17460 17604
rect 17408 17561 17417 17595
rect 17417 17561 17451 17595
rect 17451 17561 17460 17595
rect 17408 17552 17460 17561
rect 17592 17552 17644 17604
rect 16212 17484 16264 17536
rect 16304 17484 16356 17536
rect 17500 17484 17552 17536
rect 19340 17484 19392 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1492 17119 1544 17128
rect 1492 17085 1501 17119
rect 1501 17085 1535 17119
rect 1535 17085 1544 17119
rect 1492 17076 1544 17085
rect 2780 17280 2832 17332
rect 3240 17280 3292 17332
rect 4068 17280 4120 17332
rect 10968 17323 11020 17332
rect 5908 17212 5960 17264
rect 10968 17289 10977 17323
rect 10977 17289 11011 17323
rect 11011 17289 11020 17323
rect 10968 17280 11020 17289
rect 11888 17323 11940 17332
rect 11888 17289 11897 17323
rect 11897 17289 11931 17323
rect 11931 17289 11940 17323
rect 11888 17280 11940 17289
rect 19248 17280 19300 17332
rect 20444 17323 20496 17332
rect 20444 17289 20453 17323
rect 20453 17289 20487 17323
rect 20487 17289 20496 17323
rect 20444 17280 20496 17289
rect 14280 17212 14332 17264
rect 15660 17212 15712 17264
rect 16488 17255 16540 17264
rect 16488 17221 16497 17255
rect 16497 17221 16531 17255
rect 16531 17221 16540 17255
rect 16488 17212 16540 17221
rect 16948 17255 17000 17264
rect 16948 17221 16957 17255
rect 16957 17221 16991 17255
rect 16991 17221 17000 17255
rect 16948 17212 17000 17221
rect 2320 17187 2372 17196
rect 2320 17153 2329 17187
rect 2329 17153 2363 17187
rect 2363 17153 2372 17187
rect 2320 17144 2372 17153
rect 2688 17144 2740 17196
rect 6644 17144 6696 17196
rect 8484 17144 8536 17196
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 10600 17144 10652 17196
rect 3240 17119 3292 17128
rect 3240 17085 3274 17119
rect 3274 17085 3292 17119
rect 3240 17076 3292 17085
rect 4804 17076 4856 17128
rect 7104 17076 7156 17128
rect 7564 17119 7616 17128
rect 7564 17085 7598 17119
rect 7598 17085 7616 17119
rect 7564 17076 7616 17085
rect 4252 17008 4304 17060
rect 11888 17076 11940 17128
rect 16212 17144 16264 17196
rect 17316 17144 17368 17196
rect 17592 17187 17644 17196
rect 17592 17153 17601 17187
rect 17601 17153 17635 17187
rect 17635 17153 17644 17187
rect 17592 17144 17644 17153
rect 17776 17212 17828 17264
rect 13360 17076 13412 17128
rect 14464 17076 14516 17128
rect 19064 17144 19116 17196
rect 2964 16940 3016 16992
rect 4344 16983 4396 16992
rect 4344 16949 4353 16983
rect 4353 16949 4387 16983
rect 4387 16949 4396 16983
rect 4344 16940 4396 16949
rect 5264 16940 5316 16992
rect 6276 16940 6328 16992
rect 6368 16940 6420 16992
rect 7380 16940 7432 16992
rect 8208 16940 8260 16992
rect 9404 16940 9456 16992
rect 13820 17008 13872 17060
rect 15016 17008 15068 17060
rect 16212 17008 16264 17060
rect 10508 16940 10560 16992
rect 13912 16940 13964 16992
rect 14556 16983 14608 16992
rect 14556 16949 14565 16983
rect 14565 16949 14599 16983
rect 14599 16949 14608 16983
rect 14556 16940 14608 16949
rect 15108 16940 15160 16992
rect 16672 16940 16724 16992
rect 17868 17008 17920 17060
rect 19616 17008 19668 17060
rect 19340 16940 19392 16992
rect 19432 16983 19484 16992
rect 19432 16949 19441 16983
rect 19441 16949 19475 16983
rect 19475 16949 19484 16983
rect 19432 16940 19484 16949
rect 19984 16940 20036 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 2320 16736 2372 16788
rect 4712 16736 4764 16788
rect 3056 16668 3108 16720
rect 6644 16736 6696 16788
rect 7564 16736 7616 16788
rect 8300 16736 8352 16788
rect 9404 16779 9456 16788
rect 9404 16745 9413 16779
rect 9413 16745 9447 16779
rect 9447 16745 9456 16779
rect 9404 16736 9456 16745
rect 10416 16736 10468 16788
rect 10968 16736 11020 16788
rect 11612 16736 11664 16788
rect 12348 16736 12400 16788
rect 13360 16736 13412 16788
rect 13820 16779 13872 16788
rect 13820 16745 13829 16779
rect 13829 16745 13863 16779
rect 13863 16745 13872 16779
rect 13820 16736 13872 16745
rect 13912 16779 13964 16788
rect 13912 16745 13921 16779
rect 13921 16745 13955 16779
rect 13955 16745 13964 16779
rect 13912 16736 13964 16745
rect 14464 16736 14516 16788
rect 15292 16736 15344 16788
rect 15660 16779 15712 16788
rect 15660 16745 15669 16779
rect 15669 16745 15703 16779
rect 15703 16745 15712 16779
rect 15660 16736 15712 16745
rect 17592 16736 17644 16788
rect 2320 16600 2372 16652
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 2872 16532 2924 16584
rect 5724 16600 5776 16652
rect 6920 16668 6972 16720
rect 9956 16668 10008 16720
rect 4068 16532 4120 16584
rect 4344 16532 4396 16584
rect 5264 16575 5316 16584
rect 5264 16541 5273 16575
rect 5273 16541 5307 16575
rect 5307 16541 5316 16575
rect 5264 16532 5316 16541
rect 6644 16643 6696 16652
rect 6644 16609 6653 16643
rect 6653 16609 6687 16643
rect 6687 16609 6696 16643
rect 6644 16600 6696 16609
rect 7656 16600 7708 16652
rect 7472 16532 7524 16584
rect 8760 16600 8812 16652
rect 17500 16668 17552 16720
rect 19616 16736 19668 16788
rect 19800 16736 19852 16788
rect 20812 16736 20864 16788
rect 8208 16532 8260 16584
rect 10968 16532 11020 16584
rect 2412 16396 2464 16448
rect 4804 16396 4856 16448
rect 5172 16396 5224 16448
rect 6184 16439 6236 16448
rect 6184 16405 6193 16439
rect 6193 16405 6227 16439
rect 6227 16405 6236 16439
rect 6184 16396 6236 16405
rect 7288 16396 7340 16448
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 9312 16396 9364 16448
rect 9956 16396 10008 16448
rect 11704 16464 11756 16516
rect 12164 16396 12216 16448
rect 12348 16600 12400 16652
rect 13544 16600 13596 16652
rect 13636 16600 13688 16652
rect 13912 16600 13964 16652
rect 16028 16600 16080 16652
rect 12716 16532 12768 16584
rect 14004 16532 14056 16584
rect 14280 16532 14332 16584
rect 17132 16600 17184 16652
rect 17684 16600 17736 16652
rect 18052 16668 18104 16720
rect 16304 16532 16356 16584
rect 19340 16600 19392 16652
rect 12624 16396 12676 16448
rect 15200 16396 15252 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2136 16192 2188 16244
rect 4068 16235 4120 16244
rect 4068 16201 4077 16235
rect 4077 16201 4111 16235
rect 4111 16201 4120 16235
rect 4068 16192 4120 16201
rect 4712 16192 4764 16244
rect 5908 16192 5960 16244
rect 8300 16192 8352 16244
rect 10600 16192 10652 16244
rect 2320 16124 2372 16176
rect 1492 16056 1544 16108
rect 2688 16031 2740 16040
rect 2688 15997 2697 16031
rect 2697 15997 2731 16031
rect 2731 15997 2740 16031
rect 2688 15988 2740 15997
rect 2964 16031 3016 16040
rect 2964 15997 2998 16031
rect 2998 15997 3016 16031
rect 2964 15988 3016 15997
rect 4252 15988 4304 16040
rect 4804 15988 4856 16040
rect 7104 16031 7156 16040
rect 7104 15997 7113 16031
rect 7113 15997 7147 16031
rect 7147 15997 7156 16031
rect 7104 15988 7156 15997
rect 7380 16031 7432 16040
rect 7380 15997 7414 16031
rect 7414 15997 7432 16031
rect 7380 15988 7432 15997
rect 8484 15988 8536 16040
rect 10600 15988 10652 16040
rect 11704 16192 11756 16244
rect 12164 16192 12216 16244
rect 17868 16235 17920 16244
rect 11888 16124 11940 16176
rect 12992 16056 13044 16108
rect 12716 15988 12768 16040
rect 15292 16124 15344 16176
rect 16396 16124 16448 16176
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 17960 16192 18012 16244
rect 19340 16192 19392 16244
rect 19248 16056 19300 16108
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 17868 15988 17920 16040
rect 2136 15920 2188 15972
rect 6184 15920 6236 15972
rect 9128 15920 9180 15972
rect 9588 15920 9640 15972
rect 2228 15852 2280 15904
rect 3976 15852 4028 15904
rect 7472 15852 7524 15904
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 14280 15920 14332 15972
rect 13912 15852 13964 15904
rect 14004 15852 14056 15904
rect 15108 15852 15160 15904
rect 15568 15852 15620 15904
rect 16212 15852 16264 15904
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 18880 15920 18932 15972
rect 19248 15920 19300 15972
rect 19616 15852 19668 15904
rect 20168 15895 20220 15904
rect 20168 15861 20177 15895
rect 20177 15861 20211 15895
rect 20211 15861 20220 15895
rect 20168 15852 20220 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 2964 15648 3016 15700
rect 3240 15691 3292 15700
rect 3240 15657 3249 15691
rect 3249 15657 3283 15691
rect 3283 15657 3292 15691
rect 3240 15648 3292 15657
rect 4712 15648 4764 15700
rect 5264 15648 5316 15700
rect 6552 15648 6604 15700
rect 6920 15691 6972 15700
rect 6920 15657 6929 15691
rect 6929 15657 6963 15691
rect 6963 15657 6972 15691
rect 6920 15648 6972 15657
rect 8576 15648 8628 15700
rect 10232 15648 10284 15700
rect 12072 15648 12124 15700
rect 12348 15648 12400 15700
rect 13176 15648 13228 15700
rect 13912 15691 13964 15700
rect 13912 15657 13921 15691
rect 13921 15657 13955 15691
rect 13955 15657 13964 15691
rect 13912 15648 13964 15657
rect 16212 15691 16264 15700
rect 3976 15580 4028 15632
rect 14924 15623 14976 15632
rect 14924 15589 14933 15623
rect 14933 15589 14967 15623
rect 14967 15589 14976 15623
rect 14924 15580 14976 15589
rect 16212 15657 16221 15691
rect 16221 15657 16255 15691
rect 16255 15657 16264 15691
rect 16212 15648 16264 15657
rect 17868 15691 17920 15700
rect 17868 15657 17877 15691
rect 17877 15657 17911 15691
rect 17911 15657 17920 15691
rect 17868 15648 17920 15657
rect 17960 15648 18012 15700
rect 18880 15691 18932 15700
rect 18880 15657 18889 15691
rect 18889 15657 18923 15691
rect 18923 15657 18932 15691
rect 18880 15648 18932 15657
rect 19432 15691 19484 15700
rect 19432 15657 19441 15691
rect 19441 15657 19475 15691
rect 19475 15657 19484 15691
rect 19432 15648 19484 15657
rect 19616 15648 19668 15700
rect 16764 15580 16816 15632
rect 3148 15555 3200 15564
rect 3148 15521 3157 15555
rect 3157 15521 3191 15555
rect 3191 15521 3200 15555
rect 3148 15512 3200 15521
rect 4068 15512 4120 15564
rect 5816 15512 5868 15564
rect 7932 15555 7984 15564
rect 6092 15444 6144 15496
rect 6368 15444 6420 15496
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 8944 15555 8996 15564
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 7472 15487 7524 15496
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 10508 15512 10560 15564
rect 11612 15512 11664 15564
rect 13912 15512 13964 15564
rect 14740 15512 14792 15564
rect 15108 15512 15160 15564
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 10140 15444 10192 15496
rect 10600 15444 10652 15496
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 12992 15444 13044 15453
rect 14280 15444 14332 15496
rect 16304 15487 16356 15496
rect 8576 15419 8628 15428
rect 8576 15385 8585 15419
rect 8585 15385 8619 15419
rect 8619 15385 8628 15419
rect 8576 15376 8628 15385
rect 13820 15376 13872 15428
rect 16304 15453 16313 15487
rect 16313 15453 16347 15487
rect 16347 15453 16356 15487
rect 16304 15444 16356 15453
rect 17132 15444 17184 15496
rect 17960 15512 18012 15564
rect 18696 15512 18748 15564
rect 18420 15444 18472 15496
rect 19432 15444 19484 15496
rect 20168 15376 20220 15428
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 2136 15308 2188 15360
rect 5632 15351 5684 15360
rect 5632 15317 5641 15351
rect 5641 15317 5675 15351
rect 5675 15317 5684 15351
rect 5632 15308 5684 15317
rect 5724 15308 5776 15360
rect 6644 15308 6696 15360
rect 7564 15308 7616 15360
rect 11060 15308 11112 15360
rect 12348 15308 12400 15360
rect 13084 15308 13136 15360
rect 13544 15351 13596 15360
rect 13544 15317 13553 15351
rect 13553 15317 13587 15351
rect 13587 15317 13596 15351
rect 13544 15308 13596 15317
rect 15752 15308 15804 15360
rect 16396 15308 16448 15360
rect 16764 15308 16816 15360
rect 17500 15308 17552 15360
rect 17776 15351 17828 15360
rect 17776 15317 17785 15351
rect 17785 15317 17819 15351
rect 17819 15317 17828 15351
rect 17776 15308 17828 15317
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 4712 15147 4764 15156
rect 4712 15113 4721 15147
rect 4721 15113 4755 15147
rect 4755 15113 4764 15147
rect 4712 15104 4764 15113
rect 6184 15147 6236 15156
rect 6184 15113 6193 15147
rect 6193 15113 6227 15147
rect 6227 15113 6236 15147
rect 6184 15104 6236 15113
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 7932 15147 7984 15156
rect 7932 15113 7941 15147
rect 7941 15113 7975 15147
rect 7975 15113 7984 15147
rect 7932 15104 7984 15113
rect 8944 15104 8996 15156
rect 10232 15104 10284 15156
rect 10508 15104 10560 15156
rect 11152 15147 11204 15156
rect 11152 15113 11161 15147
rect 11161 15113 11195 15147
rect 11195 15113 11204 15147
rect 11152 15104 11204 15113
rect 1308 15036 1360 15088
rect 7656 15036 7708 15088
rect 2320 14968 2372 15020
rect 12348 14968 12400 15020
rect 1492 14900 1544 14952
rect 1952 14943 2004 14952
rect 1952 14909 1961 14943
rect 1961 14909 1995 14943
rect 1995 14909 2004 14943
rect 1952 14900 2004 14909
rect 2596 14832 2648 14884
rect 3148 14943 3200 14952
rect 3148 14909 3182 14943
rect 3182 14909 3200 14943
rect 4804 14943 4856 14952
rect 3148 14900 3200 14909
rect 4804 14909 4813 14943
rect 4813 14909 4847 14943
rect 4847 14909 4856 14943
rect 4804 14900 4856 14909
rect 4896 14900 4948 14952
rect 6368 14900 6420 14952
rect 7288 14943 7340 14952
rect 7288 14909 7297 14943
rect 7297 14909 7331 14943
rect 7331 14909 7340 14943
rect 7288 14900 7340 14909
rect 8484 14900 8536 14952
rect 12900 15036 12952 15088
rect 13268 15036 13320 15088
rect 16120 15104 16172 15156
rect 16396 15104 16448 15156
rect 17132 15147 17184 15156
rect 15660 15036 15712 15088
rect 17132 15113 17141 15147
rect 17141 15113 17175 15147
rect 17175 15113 17184 15147
rect 17132 15104 17184 15113
rect 19340 15104 19392 15156
rect 20168 15104 20220 15156
rect 19248 15036 19300 15088
rect 12716 14968 12768 15020
rect 12808 14900 12860 14952
rect 13084 14943 13136 14952
rect 13084 14909 13093 14943
rect 13093 14909 13127 14943
rect 13127 14909 13136 14943
rect 14004 14968 14056 15020
rect 14832 15011 14884 15020
rect 14832 14977 14841 15011
rect 14841 14977 14875 15011
rect 14875 14977 14884 15011
rect 14832 14968 14884 14977
rect 15200 14968 15252 15020
rect 15752 15011 15804 15020
rect 15752 14977 15761 15011
rect 15761 14977 15795 15011
rect 15795 14977 15804 15011
rect 15752 14968 15804 14977
rect 16856 14968 16908 15020
rect 17684 14968 17736 15020
rect 13084 14900 13136 14909
rect 13912 14900 13964 14952
rect 14280 14900 14332 14952
rect 14740 14943 14792 14952
rect 8852 14832 8904 14884
rect 9312 14832 9364 14884
rect 9404 14832 9456 14884
rect 10140 14832 10192 14884
rect 3056 14764 3108 14816
rect 4068 14764 4120 14816
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 9128 14764 9180 14816
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 11704 14764 11756 14773
rect 12532 14764 12584 14816
rect 12624 14807 12676 14816
rect 12624 14773 12633 14807
rect 12633 14773 12667 14807
rect 12667 14773 12676 14807
rect 12624 14764 12676 14773
rect 12992 14764 13044 14816
rect 13084 14764 13136 14816
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 14740 14909 14749 14943
rect 14749 14909 14783 14943
rect 14783 14909 14792 14943
rect 14740 14900 14792 14909
rect 15384 14943 15436 14952
rect 15384 14909 15393 14943
rect 15393 14909 15427 14943
rect 15427 14909 15436 14943
rect 15384 14900 15436 14909
rect 16304 14900 16356 14952
rect 16764 14832 16816 14884
rect 17316 14832 17368 14884
rect 17960 14832 18012 14884
rect 18328 14900 18380 14952
rect 19432 14900 19484 14952
rect 19616 14900 19668 14952
rect 17500 14764 17552 14816
rect 19432 14764 19484 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 2044 14560 2096 14612
rect 4160 14560 4212 14612
rect 7748 14560 7800 14612
rect 8944 14560 8996 14612
rect 10140 14603 10192 14612
rect 10140 14569 10149 14603
rect 10149 14569 10183 14603
rect 10183 14569 10192 14603
rect 10140 14560 10192 14569
rect 12808 14560 12860 14612
rect 5724 14492 5776 14544
rect 7380 14492 7432 14544
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 2228 14424 2280 14476
rect 3332 14467 3384 14476
rect 3332 14433 3341 14467
rect 3341 14433 3375 14467
rect 3375 14433 3384 14467
rect 3332 14424 3384 14433
rect 3608 14424 3660 14476
rect 4712 14424 4764 14476
rect 6920 14467 6972 14476
rect 6920 14433 6954 14467
rect 6954 14433 6972 14467
rect 6920 14424 6972 14433
rect 7472 14424 7524 14476
rect 9128 14492 9180 14544
rect 15660 14560 15712 14612
rect 18512 14560 18564 14612
rect 18972 14560 19024 14612
rect 10324 14424 10376 14476
rect 1492 14356 1544 14408
rect 2320 14356 2372 14408
rect 4160 14356 4212 14408
rect 2596 14288 2648 14340
rect 2872 14263 2924 14272
rect 2872 14229 2881 14263
rect 2881 14229 2915 14263
rect 2915 14229 2924 14263
rect 3976 14288 4028 14340
rect 4804 14356 4856 14408
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 11704 14356 11756 14408
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 12348 14424 12400 14476
rect 13728 14424 13780 14476
rect 13820 14424 13872 14476
rect 14096 14424 14148 14476
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 13268 14399 13320 14408
rect 12440 14356 12492 14365
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 14556 14424 14608 14476
rect 6276 14288 6328 14340
rect 12624 14288 12676 14340
rect 12900 14288 12952 14340
rect 15200 14356 15252 14408
rect 15384 14424 15436 14476
rect 15936 14424 15988 14476
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 18420 14492 18472 14544
rect 18788 14492 18840 14544
rect 19248 14492 19300 14544
rect 19340 14492 19392 14544
rect 16764 14356 16816 14408
rect 16856 14356 16908 14408
rect 15384 14288 15436 14340
rect 16304 14288 16356 14340
rect 16580 14288 16632 14340
rect 17960 14356 18012 14408
rect 18420 14399 18472 14408
rect 18420 14365 18429 14399
rect 18429 14365 18463 14399
rect 18463 14365 18472 14399
rect 18420 14356 18472 14365
rect 17776 14288 17828 14340
rect 2872 14220 2924 14229
rect 3608 14220 3660 14272
rect 6092 14263 6144 14272
rect 6092 14229 6101 14263
rect 6101 14229 6135 14263
rect 6135 14229 6144 14263
rect 6092 14220 6144 14229
rect 7380 14220 7432 14272
rect 8668 14263 8720 14272
rect 8668 14229 8677 14263
rect 8677 14229 8711 14263
rect 8711 14229 8720 14263
rect 8668 14220 8720 14229
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 14280 14220 14332 14272
rect 14464 14220 14516 14272
rect 19800 14263 19852 14272
rect 19800 14229 19809 14263
rect 19809 14229 19843 14263
rect 19843 14229 19852 14263
rect 19800 14220 19852 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2780 14016 2832 14068
rect 1400 13880 1452 13932
rect 3332 14016 3384 14068
rect 4160 14016 4212 14068
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 5264 13991 5316 14000
rect 5264 13957 5273 13991
rect 5273 13957 5307 13991
rect 5307 13957 5316 13991
rect 5264 13948 5316 13957
rect 6920 14016 6972 14068
rect 10140 14016 10192 14068
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 2596 13812 2648 13864
rect 3700 13812 3752 13864
rect 4160 13855 4212 13864
rect 4160 13821 4194 13855
rect 4194 13821 4212 13855
rect 4160 13812 4212 13821
rect 5908 13812 5960 13864
rect 13820 14016 13872 14068
rect 6276 13923 6328 13932
rect 6276 13889 6285 13923
rect 6285 13889 6319 13923
rect 6319 13889 6328 13923
rect 7380 13923 7432 13932
rect 6276 13880 6328 13889
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 15660 13948 15712 14000
rect 18604 13948 18656 14000
rect 19432 13991 19484 14000
rect 7196 13855 7248 13864
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 7564 13812 7616 13864
rect 8484 13812 8536 13864
rect 8668 13855 8720 13864
rect 8668 13821 8702 13855
rect 8702 13821 8720 13855
rect 8668 13812 8720 13821
rect 9588 13812 9640 13864
rect 10600 13855 10652 13864
rect 10600 13821 10609 13855
rect 10609 13821 10643 13855
rect 10643 13821 10652 13855
rect 10600 13812 10652 13821
rect 11152 13812 11204 13864
rect 12348 13812 12400 13864
rect 4804 13744 4856 13796
rect 6092 13787 6144 13796
rect 6092 13753 6101 13787
rect 6101 13753 6135 13787
rect 6135 13753 6144 13787
rect 6092 13744 6144 13753
rect 9772 13744 9824 13796
rect 10692 13744 10744 13796
rect 13820 13812 13872 13864
rect 16396 13812 16448 13864
rect 16580 13855 16632 13864
rect 16580 13821 16614 13855
rect 16614 13821 16632 13855
rect 16580 13812 16632 13821
rect 14372 13744 14424 13796
rect 7748 13676 7800 13728
rect 9680 13676 9732 13728
rect 11980 13719 12032 13728
rect 11980 13685 11989 13719
rect 11989 13685 12023 13719
rect 12023 13685 12032 13719
rect 11980 13676 12032 13685
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 13268 13676 13320 13728
rect 13728 13676 13780 13728
rect 15384 13719 15436 13728
rect 15384 13685 15393 13719
rect 15393 13685 15427 13719
rect 15427 13685 15436 13719
rect 15384 13676 15436 13685
rect 17684 13719 17736 13728
rect 17684 13685 17693 13719
rect 17693 13685 17727 13719
rect 17727 13685 17736 13719
rect 18972 13880 19024 13932
rect 17960 13812 18012 13864
rect 19432 13957 19441 13991
rect 19441 13957 19475 13991
rect 19475 13957 19484 13991
rect 19432 13948 19484 13957
rect 19800 13991 19852 14000
rect 19800 13957 19809 13991
rect 19809 13957 19843 13991
rect 19843 13957 19852 13991
rect 19800 13948 19852 13957
rect 19248 13880 19300 13932
rect 18512 13787 18564 13796
rect 18512 13753 18521 13787
rect 18521 13753 18555 13787
rect 18555 13753 18564 13787
rect 18512 13744 18564 13753
rect 17684 13676 17736 13685
rect 19156 13676 19208 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 2872 13472 2924 13524
rect 4712 13472 4764 13524
rect 5356 13472 5408 13524
rect 7196 13472 7248 13524
rect 7288 13472 7340 13524
rect 8208 13472 8260 13524
rect 9772 13472 9824 13524
rect 1584 13404 1636 13456
rect 13452 13472 13504 13524
rect 13636 13472 13688 13524
rect 1400 13379 1452 13388
rect 1400 13345 1409 13379
rect 1409 13345 1443 13379
rect 1443 13345 1452 13379
rect 1400 13336 1452 13345
rect 1676 13336 1728 13388
rect 1952 13379 2004 13388
rect 1952 13345 1961 13379
rect 1961 13345 1995 13379
rect 1995 13345 2004 13379
rect 1952 13336 2004 13345
rect 4160 13336 4212 13388
rect 5172 13379 5224 13388
rect 5172 13345 5206 13379
rect 5206 13345 5224 13379
rect 5172 13336 5224 13345
rect 3424 13268 3476 13320
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 4804 13200 4856 13252
rect 6092 13132 6144 13184
rect 7380 13336 7432 13388
rect 6368 13268 6420 13320
rect 6644 13311 6696 13320
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 8852 13336 8904 13388
rect 9496 13336 9548 13388
rect 13084 13404 13136 13456
rect 13728 13404 13780 13456
rect 12532 13336 12584 13388
rect 13176 13336 13228 13388
rect 13820 13336 13872 13388
rect 14372 13472 14424 13524
rect 15384 13472 15436 13524
rect 16948 13515 17000 13524
rect 16948 13481 16957 13515
rect 16957 13481 16991 13515
rect 16991 13481 17000 13515
rect 16948 13472 17000 13481
rect 18788 13515 18840 13524
rect 18788 13481 18797 13515
rect 18797 13481 18831 13515
rect 18831 13481 18840 13515
rect 18788 13472 18840 13481
rect 18880 13472 18932 13524
rect 15568 13404 15620 13456
rect 15936 13447 15988 13456
rect 15936 13413 15945 13447
rect 15945 13413 15979 13447
rect 15979 13413 15988 13447
rect 15936 13404 15988 13413
rect 17684 13404 17736 13456
rect 18512 13404 18564 13456
rect 9680 13268 9732 13320
rect 10140 13268 10192 13320
rect 12624 13268 12676 13320
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 11980 13200 12032 13252
rect 13084 13268 13136 13320
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 14464 13268 14516 13320
rect 15660 13268 15712 13320
rect 18696 13268 18748 13320
rect 19156 13268 19208 13320
rect 6368 13132 6420 13184
rect 8668 13132 8720 13184
rect 8760 13132 8812 13184
rect 12716 13132 12768 13184
rect 13636 13132 13688 13184
rect 16580 13200 16632 13252
rect 16948 13200 17000 13252
rect 18052 13200 18104 13252
rect 14832 13132 14884 13184
rect 18604 13132 18656 13184
rect 19064 13175 19116 13184
rect 19064 13141 19073 13175
rect 19073 13141 19107 13175
rect 19107 13141 19116 13175
rect 19064 13132 19116 13141
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1860 12928 1912 12980
rect 1400 12792 1452 12844
rect 1584 12792 1636 12844
rect 4160 12835 4212 12844
rect 4160 12801 4169 12835
rect 4169 12801 4203 12835
rect 4203 12801 4212 12835
rect 4160 12792 4212 12801
rect 4252 12792 4304 12844
rect 4712 12928 4764 12980
rect 4896 12928 4948 12980
rect 5172 12928 5224 12980
rect 5540 12860 5592 12912
rect 9220 12928 9272 12980
rect 9588 12971 9640 12980
rect 9588 12937 9597 12971
rect 9597 12937 9631 12971
rect 9631 12937 9640 12971
rect 9588 12928 9640 12937
rect 11796 12928 11848 12980
rect 14280 12928 14332 12980
rect 15568 12928 15620 12980
rect 18512 12928 18564 12980
rect 19064 12971 19116 12980
rect 19064 12937 19073 12971
rect 19073 12937 19107 12971
rect 19107 12937 19116 12971
rect 19064 12928 19116 12937
rect 9496 12860 9548 12912
rect 13912 12860 13964 12912
rect 1492 12767 1544 12776
rect 1492 12733 1501 12767
rect 1501 12733 1535 12767
rect 1535 12733 1544 12767
rect 1492 12724 1544 12733
rect 2044 12767 2096 12776
rect 2044 12733 2053 12767
rect 2053 12733 2087 12767
rect 2087 12733 2096 12767
rect 2044 12724 2096 12733
rect 1400 12656 1452 12708
rect 2136 12656 2188 12708
rect 7564 12724 7616 12776
rect 10140 12792 10192 12844
rect 9680 12724 9732 12776
rect 11796 12792 11848 12844
rect 12440 12792 12492 12844
rect 13084 12835 13136 12844
rect 13084 12801 13093 12835
rect 13093 12801 13127 12835
rect 13127 12801 13136 12835
rect 14280 12835 14332 12844
rect 13084 12792 13136 12801
rect 4804 12699 4856 12708
rect 4804 12665 4838 12699
rect 4838 12665 4856 12699
rect 4804 12656 4856 12665
rect 5540 12656 5592 12708
rect 2044 12588 2096 12640
rect 5080 12588 5132 12640
rect 7196 12631 7248 12640
rect 7196 12597 7205 12631
rect 7205 12597 7239 12631
rect 7239 12597 7248 12631
rect 7196 12588 7248 12597
rect 8576 12588 8628 12640
rect 11980 12656 12032 12708
rect 11704 12588 11756 12640
rect 12256 12588 12308 12640
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12900 12631 12952 12640
rect 12440 12588 12492 12597
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 14372 12835 14424 12844
rect 14372 12801 14381 12835
rect 14381 12801 14415 12835
rect 14415 12801 14424 12835
rect 14832 12835 14884 12844
rect 14372 12792 14424 12801
rect 14832 12801 14841 12835
rect 14841 12801 14875 12835
rect 14875 12801 14884 12835
rect 14832 12792 14884 12801
rect 19432 12835 19484 12844
rect 19432 12801 19441 12835
rect 19441 12801 19475 12835
rect 19475 12801 19484 12835
rect 19432 12792 19484 12801
rect 15200 12724 15252 12776
rect 17592 12724 17644 12776
rect 17960 12724 18012 12776
rect 13912 12656 13964 12708
rect 14556 12656 14608 12708
rect 18512 12699 18564 12708
rect 15016 12588 15068 12640
rect 17132 12588 17184 12640
rect 17592 12631 17644 12640
rect 17592 12597 17601 12631
rect 17601 12597 17635 12631
rect 17635 12597 17644 12631
rect 17592 12588 17644 12597
rect 18512 12665 18521 12699
rect 18521 12665 18555 12699
rect 18555 12665 18564 12699
rect 18512 12656 18564 12665
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 1768 12427 1820 12436
rect 1768 12393 1777 12427
rect 1777 12393 1811 12427
rect 1811 12393 1820 12427
rect 1768 12384 1820 12393
rect 2964 12384 3016 12436
rect 1952 12316 2004 12368
rect 6276 12384 6328 12436
rect 6368 12384 6420 12436
rect 8852 12384 8904 12436
rect 9772 12384 9824 12436
rect 11060 12384 11112 12436
rect 11888 12384 11940 12436
rect 14280 12384 14332 12436
rect 16764 12384 16816 12436
rect 17132 12384 17184 12436
rect 4068 12316 4120 12368
rect 12900 12316 12952 12368
rect 13636 12316 13688 12368
rect 15200 12316 15252 12368
rect 18512 12384 18564 12436
rect 21364 12384 21416 12436
rect 1676 12248 1728 12300
rect 2228 12248 2280 12300
rect 3240 12248 3292 12300
rect 1492 12180 1544 12232
rect 1768 12180 1820 12232
rect 4712 12248 4764 12300
rect 5448 12248 5500 12300
rect 6184 12291 6236 12300
rect 6184 12257 6218 12291
rect 6218 12257 6236 12291
rect 6184 12248 6236 12257
rect 7564 12248 7616 12300
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 8208 12248 8260 12300
rect 8576 12291 8628 12300
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 9496 12248 9548 12300
rect 10140 12248 10192 12300
rect 11704 12248 11756 12300
rect 12256 12248 12308 12300
rect 12440 12248 12492 12300
rect 12808 12248 12860 12300
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 5540 12180 5592 12232
rect 7840 12180 7892 12232
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 8852 12223 8904 12232
rect 8852 12189 8861 12223
rect 8861 12189 8895 12223
rect 8895 12189 8904 12223
rect 8852 12180 8904 12189
rect 9588 12180 9640 12232
rect 10048 12180 10100 12232
rect 5724 12112 5776 12164
rect 3792 12087 3844 12096
rect 3792 12053 3801 12087
rect 3801 12053 3835 12087
rect 3835 12053 3844 12087
rect 3792 12044 3844 12053
rect 11060 12180 11112 12232
rect 12716 12180 12768 12232
rect 12900 12180 12952 12232
rect 13452 12180 13504 12232
rect 14372 12248 14424 12300
rect 14556 12248 14608 12300
rect 15568 12248 15620 12300
rect 16304 12248 16356 12300
rect 17684 12248 17736 12300
rect 15016 12180 15068 12232
rect 15200 12180 15252 12232
rect 17776 12180 17828 12232
rect 18604 12248 18656 12300
rect 19800 12248 19852 12300
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 16672 12112 16724 12164
rect 16948 12112 17000 12164
rect 17592 12112 17644 12164
rect 7380 12044 7432 12096
rect 7472 12044 7524 12096
rect 7656 12044 7708 12096
rect 8944 12044 8996 12096
rect 11796 12044 11848 12096
rect 12716 12044 12768 12096
rect 13452 12044 13504 12096
rect 16212 12044 16264 12096
rect 17684 12044 17736 12096
rect 20444 12044 20496 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 4896 11840 4948 11892
rect 3792 11772 3844 11824
rect 6828 11840 6880 11892
rect 9680 11840 9732 11892
rect 10140 11883 10192 11892
rect 10140 11849 10149 11883
rect 10149 11849 10183 11883
rect 10183 11849 10192 11883
rect 10140 11840 10192 11849
rect 11704 11840 11756 11892
rect 12164 11840 12216 11892
rect 9496 11815 9548 11824
rect 9496 11781 9505 11815
rect 9505 11781 9539 11815
rect 9539 11781 9548 11815
rect 9496 11772 9548 11781
rect 11888 11815 11940 11824
rect 11888 11781 11897 11815
rect 11897 11781 11931 11815
rect 11931 11781 11940 11815
rect 11888 11772 11940 11781
rect 13452 11840 13504 11892
rect 19432 11883 19484 11892
rect 2504 11636 2556 11688
rect 2872 11636 2924 11688
rect 4160 11636 4212 11688
rect 5264 11636 5316 11688
rect 5540 11636 5592 11688
rect 5724 11636 5776 11688
rect 6368 11704 6420 11756
rect 6460 11704 6512 11756
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 7012 11636 7064 11688
rect 7656 11636 7708 11688
rect 3056 11611 3108 11620
rect 3056 11577 3090 11611
rect 3090 11577 3108 11611
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 3056 11568 3108 11577
rect 4068 11568 4120 11620
rect 10048 11636 10100 11688
rect 8944 11568 8996 11620
rect 11060 11636 11112 11688
rect 12716 11772 12768 11824
rect 13268 11772 13320 11824
rect 14096 11772 14148 11824
rect 16304 11815 16356 11824
rect 16304 11781 16313 11815
rect 16313 11781 16347 11815
rect 16347 11781 16356 11815
rect 16304 11772 16356 11781
rect 17592 11772 17644 11824
rect 17776 11815 17828 11824
rect 17776 11781 17785 11815
rect 17785 11781 17819 11815
rect 17819 11781 17828 11815
rect 17776 11772 17828 11781
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 12808 11679 12860 11688
rect 12164 11568 12216 11620
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 13268 11636 13320 11688
rect 13452 11636 13504 11688
rect 18052 11679 18104 11688
rect 12532 11568 12584 11620
rect 13636 11611 13688 11620
rect 3240 11500 3292 11552
rect 3700 11500 3752 11552
rect 4436 11543 4488 11552
rect 4436 11509 4445 11543
rect 4445 11509 4479 11543
rect 4479 11509 4488 11543
rect 4436 11500 4488 11509
rect 4804 11543 4856 11552
rect 4804 11509 4813 11543
rect 4813 11509 4847 11543
rect 4847 11509 4856 11543
rect 4804 11500 4856 11509
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 5264 11500 5316 11552
rect 6276 11500 6328 11552
rect 7196 11543 7248 11552
rect 7196 11509 7205 11543
rect 7205 11509 7239 11543
rect 7239 11509 7248 11543
rect 7196 11500 7248 11509
rect 7656 11500 7708 11552
rect 10048 11500 10100 11552
rect 10692 11500 10744 11552
rect 11888 11500 11940 11552
rect 12716 11500 12768 11552
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 13636 11577 13645 11611
rect 13645 11577 13679 11611
rect 13679 11577 13688 11611
rect 13636 11568 13688 11577
rect 13728 11611 13780 11620
rect 13728 11577 13737 11611
rect 13737 11577 13771 11611
rect 13771 11577 13780 11611
rect 13728 11568 13780 11577
rect 14188 11568 14240 11620
rect 14372 11611 14424 11620
rect 14372 11577 14381 11611
rect 14381 11577 14415 11611
rect 14415 11577 14424 11611
rect 14372 11568 14424 11577
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 15476 11568 15528 11620
rect 15660 11568 15712 11620
rect 15568 11500 15620 11552
rect 16672 11500 16724 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 18144 11568 18196 11620
rect 18604 11568 18656 11620
rect 19248 11568 19300 11620
rect 19616 11500 19668 11552
rect 19800 11543 19852 11552
rect 19800 11509 19809 11543
rect 19809 11509 19843 11543
rect 19843 11509 19852 11543
rect 19800 11500 19852 11509
rect 20444 11500 20496 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2504 11296 2556 11348
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 4528 11296 4580 11348
rect 5172 11296 5224 11348
rect 5448 11296 5500 11348
rect 7196 11296 7248 11348
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 9404 11296 9456 11348
rect 10140 11296 10192 11348
rect 10876 11296 10928 11348
rect 13452 11296 13504 11348
rect 13820 11296 13872 11348
rect 1676 11228 1728 11280
rect 1952 11160 2004 11212
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 2504 11160 2556 11169
rect 2044 11092 2096 11144
rect 2228 11092 2280 11144
rect 4712 11203 4764 11212
rect 4712 11169 4721 11203
rect 4721 11169 4755 11203
rect 4755 11169 4764 11203
rect 4712 11160 4764 11169
rect 6000 11160 6052 11212
rect 6276 11203 6328 11212
rect 6276 11169 6285 11203
rect 6285 11169 6319 11203
rect 6319 11169 6328 11203
rect 6276 11160 6328 11169
rect 2688 11092 2740 11144
rect 3056 11092 3108 11144
rect 6460 11092 6512 11144
rect 4068 11024 4120 11076
rect 7288 11160 7340 11212
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 6644 11024 6696 11076
rect 2228 10956 2280 11008
rect 2504 10956 2556 11008
rect 2872 10956 2924 11008
rect 3976 10956 4028 11008
rect 6920 10956 6972 11008
rect 7656 11160 7708 11212
rect 8208 11160 8260 11212
rect 8852 11228 8904 11280
rect 11796 11228 11848 11280
rect 12532 11228 12584 11280
rect 12900 11228 12952 11280
rect 13912 11228 13964 11280
rect 15660 11296 15712 11348
rect 16948 11296 17000 11348
rect 17960 11296 18012 11348
rect 19432 11296 19484 11348
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 20444 11339 20496 11348
rect 20444 11305 20453 11339
rect 20453 11305 20487 11339
rect 20487 11305 20496 11339
rect 20444 11296 20496 11305
rect 15384 11228 15436 11280
rect 18512 11228 18564 11280
rect 19248 11271 19300 11280
rect 19248 11237 19257 11271
rect 19257 11237 19291 11271
rect 19291 11237 19300 11271
rect 19248 11228 19300 11237
rect 11060 11160 11112 11212
rect 14556 11203 14608 11212
rect 10692 11092 10744 11144
rect 8576 11024 8628 11076
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 14648 11203 14700 11212
rect 14648 11169 14657 11203
rect 14657 11169 14691 11203
rect 14691 11169 14700 11203
rect 14648 11160 14700 11169
rect 15016 11160 15068 11212
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 16212 11160 16264 11212
rect 17776 11160 17828 11212
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 15108 11092 15160 11144
rect 15292 11092 15344 11144
rect 14648 11024 14700 11076
rect 15476 11024 15528 11076
rect 16672 11092 16724 11144
rect 18144 11135 18196 11144
rect 18144 11101 18153 11135
rect 18153 11101 18187 11135
rect 18187 11101 18196 11135
rect 18144 11092 18196 11101
rect 19340 11092 19392 11144
rect 16120 11024 16172 11076
rect 18788 11024 18840 11076
rect 20536 11024 20588 11076
rect 8208 10956 8260 11008
rect 8944 10956 8996 11008
rect 9864 10999 9916 11008
rect 9864 10965 9873 10999
rect 9873 10965 9907 10999
rect 9907 10965 9916 10999
rect 9864 10956 9916 10965
rect 12900 10956 12952 11008
rect 13084 10956 13136 11008
rect 16396 10956 16448 11008
rect 17960 10956 18012 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 4068 10752 4120 10804
rect 5172 10795 5224 10804
rect 5172 10761 5181 10795
rect 5181 10761 5215 10795
rect 5215 10761 5224 10795
rect 5172 10752 5224 10761
rect 6092 10752 6144 10804
rect 8576 10752 8628 10804
rect 8760 10752 8812 10804
rect 12716 10752 12768 10804
rect 15476 10795 15528 10804
rect 15476 10761 15485 10795
rect 15485 10761 15519 10795
rect 15519 10761 15528 10795
rect 15476 10752 15528 10761
rect 17960 10752 18012 10804
rect 20536 10795 20588 10804
rect 6644 10727 6696 10736
rect 6644 10693 6653 10727
rect 6653 10693 6687 10727
rect 6687 10693 6696 10727
rect 6644 10684 6696 10693
rect 8208 10727 8260 10736
rect 8208 10693 8217 10727
rect 8217 10693 8251 10727
rect 8251 10693 8260 10727
rect 8208 10684 8260 10693
rect 8944 10684 8996 10736
rect 2504 10616 2556 10668
rect 3240 10616 3292 10668
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 5724 10616 5776 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 10876 10616 10928 10668
rect 11980 10616 12032 10668
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 20536 10761 20545 10795
rect 20545 10761 20579 10795
rect 20579 10761 20588 10795
rect 20536 10752 20588 10761
rect 19616 10684 19668 10736
rect 20444 10684 20496 10736
rect 1308 10548 1360 10600
rect 1492 10548 1544 10600
rect 2320 10548 2372 10600
rect 5540 10548 5592 10600
rect 8852 10591 8904 10600
rect 3056 10480 3108 10532
rect 4712 10480 4764 10532
rect 7104 10523 7156 10532
rect 7104 10489 7138 10523
rect 7138 10489 7156 10523
rect 7104 10480 7156 10489
rect 1952 10412 2004 10464
rect 2320 10412 2372 10464
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 3332 10412 3384 10464
rect 3976 10412 4028 10464
rect 5724 10412 5776 10464
rect 7012 10412 7064 10464
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 9404 10548 9456 10600
rect 11060 10548 11112 10600
rect 11704 10548 11756 10600
rect 13452 10548 13504 10600
rect 15568 10548 15620 10600
rect 16396 10548 16448 10600
rect 19432 10548 19484 10600
rect 10784 10480 10836 10532
rect 11520 10480 11572 10532
rect 13084 10480 13136 10532
rect 15108 10480 15160 10532
rect 16028 10523 16080 10532
rect 16028 10489 16062 10523
rect 16062 10489 16080 10523
rect 16028 10480 16080 10489
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 12808 10412 12860 10464
rect 13728 10412 13780 10464
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 2228 10208 2280 10260
rect 2504 10208 2556 10260
rect 6184 10208 6236 10260
rect 10324 10208 10376 10260
rect 13084 10251 13136 10260
rect 1768 10183 1820 10192
rect 1768 10149 1777 10183
rect 1777 10149 1811 10183
rect 1811 10149 1820 10183
rect 1768 10140 1820 10149
rect 2228 10115 2280 10124
rect 2228 10081 2237 10115
rect 2237 10081 2271 10115
rect 2271 10081 2280 10115
rect 2228 10072 2280 10081
rect 2688 10140 2740 10192
rect 2964 10140 3016 10192
rect 3516 10072 3568 10124
rect 5724 10140 5776 10192
rect 13084 10217 13093 10251
rect 13093 10217 13127 10251
rect 13127 10217 13136 10251
rect 13084 10208 13136 10217
rect 18512 10208 18564 10260
rect 18788 10251 18840 10260
rect 18788 10217 18797 10251
rect 18797 10217 18831 10251
rect 18831 10217 18840 10251
rect 18788 10208 18840 10217
rect 19616 10251 19668 10260
rect 19616 10217 19625 10251
rect 19625 10217 19659 10251
rect 19659 10217 19668 10251
rect 19616 10208 19668 10217
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 20536 10208 20588 10260
rect 13728 10140 13780 10192
rect 15292 10140 15344 10192
rect 15844 10183 15896 10192
rect 15844 10149 15853 10183
rect 15853 10149 15887 10183
rect 15887 10149 15896 10183
rect 15844 10140 15896 10149
rect 17132 10140 17184 10192
rect 6000 10115 6052 10124
rect 6000 10081 6034 10115
rect 6034 10081 6052 10115
rect 6000 10072 6052 10081
rect 6828 10072 6880 10124
rect 6920 10072 6972 10124
rect 7472 10072 7524 10124
rect 8760 10072 8812 10124
rect 8852 10072 8904 10124
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 10692 10072 10744 10124
rect 11704 10115 11756 10124
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 11704 10072 11756 10081
rect 11980 10115 12032 10124
rect 11980 10081 12014 10115
rect 12014 10081 12032 10115
rect 11980 10072 12032 10081
rect 13452 10072 13504 10124
rect 14096 10072 14148 10124
rect 15936 10072 15988 10124
rect 16396 10115 16448 10124
rect 16396 10081 16405 10115
rect 16405 10081 16439 10115
rect 16439 10081 16448 10115
rect 16396 10072 16448 10081
rect 18604 10072 18656 10124
rect 3332 10047 3384 10056
rect 3056 9936 3108 9988
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 5540 10004 5592 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 7104 9979 7156 9988
rect 2320 9868 2372 9920
rect 7104 9945 7113 9979
rect 7113 9945 7147 9979
rect 7147 9945 7156 9979
rect 7104 9936 7156 9945
rect 15108 9936 15160 9988
rect 3884 9868 3936 9920
rect 6092 9868 6144 9920
rect 6920 9868 6972 9920
rect 7196 9868 7248 9920
rect 7656 9868 7708 9920
rect 10968 9868 11020 9920
rect 11980 9868 12032 9920
rect 17040 9868 17092 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 1768 9707 1820 9716
rect 1768 9673 1777 9707
rect 1777 9673 1811 9707
rect 1811 9673 1820 9707
rect 1768 9664 1820 9673
rect 2504 9664 2556 9716
rect 2872 9664 2924 9716
rect 3424 9664 3476 9716
rect 4068 9664 4120 9716
rect 15660 9664 15712 9716
rect 15844 9664 15896 9716
rect 17408 9664 17460 9716
rect 19616 9664 19668 9716
rect 5080 9596 5132 9648
rect 6552 9596 6604 9648
rect 6920 9596 6972 9648
rect 2688 9460 2740 9512
rect 4068 9528 4120 9580
rect 5724 9528 5776 9580
rect 7104 9528 7156 9580
rect 9956 9596 10008 9648
rect 10140 9596 10192 9648
rect 7656 9528 7708 9580
rect 8208 9528 8260 9580
rect 12440 9596 12492 9648
rect 13820 9596 13872 9648
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 12716 9528 12768 9580
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 14556 9596 14608 9648
rect 19156 9596 19208 9648
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 17776 9528 17828 9580
rect 19340 9528 19392 9580
rect 19984 9528 20036 9580
rect 2504 9392 2556 9444
rect 6552 9460 6604 9512
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 7472 9460 7524 9512
rect 5816 9392 5868 9444
rect 6460 9392 6512 9444
rect 9680 9392 9732 9444
rect 10876 9460 10928 9512
rect 11520 9460 11572 9512
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 15200 9460 15252 9512
rect 17408 9460 17460 9512
rect 16304 9392 16356 9444
rect 17040 9435 17092 9444
rect 17040 9401 17049 9435
rect 17049 9401 17083 9435
rect 17083 9401 17092 9435
rect 17040 9392 17092 9401
rect 3240 9367 3292 9376
rect 3240 9333 3249 9367
rect 3249 9333 3283 9367
rect 3283 9333 3292 9367
rect 3240 9324 3292 9333
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 4068 9324 4120 9376
rect 4712 9324 4764 9376
rect 5080 9324 5132 9376
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 6552 9324 6604 9376
rect 6920 9324 6972 9376
rect 9496 9324 9548 9376
rect 9588 9324 9640 9376
rect 9864 9324 9916 9376
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 10784 9324 10836 9376
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12440 9324 12492 9333
rect 15108 9324 15160 9376
rect 15936 9324 15988 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2228 9120 2280 9172
rect 5724 9163 5776 9172
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 6368 9163 6420 9172
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 7196 9120 7248 9172
rect 7380 9120 7432 9172
rect 8576 9120 8628 9172
rect 10048 9120 10100 9172
rect 10968 9120 11020 9172
rect 11520 9163 11572 9172
rect 11520 9129 11529 9163
rect 11529 9129 11563 9163
rect 11563 9129 11572 9163
rect 11520 9120 11572 9129
rect 12808 9163 12860 9172
rect 12808 9129 12817 9163
rect 12817 9129 12851 9163
rect 12851 9129 12860 9163
rect 12808 9120 12860 9129
rect 13084 9120 13136 9172
rect 15108 9120 15160 9172
rect 15476 9120 15528 9172
rect 17132 9120 17184 9172
rect 17500 9120 17552 9172
rect 19340 9120 19392 9172
rect 3332 9052 3384 9104
rect 4160 9052 4212 9104
rect 2136 8984 2188 9036
rect 2964 8984 3016 9036
rect 5356 8984 5408 9036
rect 6828 8984 6880 9036
rect 9036 8984 9088 9036
rect 9588 8984 9640 9036
rect 15016 9052 15068 9104
rect 16856 9052 16908 9104
rect 16028 8984 16080 9036
rect 17040 8984 17092 9036
rect 2504 8916 2556 8968
rect 6920 8916 6972 8968
rect 8484 8916 8536 8968
rect 1032 8848 1084 8900
rect 4068 8848 4120 8900
rect 4988 8848 5040 8900
rect 9680 8916 9732 8968
rect 10692 8916 10744 8968
rect 3148 8780 3200 8832
rect 4252 8780 4304 8832
rect 4712 8780 4764 8832
rect 5080 8780 5132 8832
rect 5356 8823 5408 8832
rect 5356 8789 5365 8823
rect 5365 8789 5399 8823
rect 5399 8789 5408 8823
rect 5356 8780 5408 8789
rect 6276 8780 6328 8832
rect 8760 8780 8812 8832
rect 9220 8848 9272 8900
rect 10784 8891 10836 8900
rect 10784 8857 10793 8891
rect 10793 8857 10827 8891
rect 10827 8857 10836 8891
rect 10784 8848 10836 8857
rect 10140 8780 10192 8832
rect 11980 8780 12032 8832
rect 13728 8780 13780 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 3516 8576 3568 8628
rect 3884 8619 3936 8628
rect 3884 8585 3893 8619
rect 3893 8585 3927 8619
rect 3927 8585 3936 8619
rect 3884 8576 3936 8585
rect 4252 8576 4304 8628
rect 5172 8576 5224 8628
rect 6920 8619 6972 8628
rect 6920 8585 6929 8619
rect 6929 8585 6963 8619
rect 6963 8585 6972 8619
rect 6920 8576 6972 8585
rect 9680 8576 9732 8628
rect 10968 8576 11020 8628
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 11980 8619 12032 8628
rect 11980 8585 11989 8619
rect 11989 8585 12023 8619
rect 12023 8585 12032 8619
rect 11980 8576 12032 8585
rect 12900 8576 12952 8628
rect 13728 8619 13780 8628
rect 13728 8585 13737 8619
rect 13737 8585 13771 8619
rect 13771 8585 13780 8619
rect 13728 8576 13780 8585
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 16028 8619 16080 8628
rect 16028 8585 16037 8619
rect 16037 8585 16071 8619
rect 16071 8585 16080 8619
rect 16028 8576 16080 8585
rect 16396 8619 16448 8628
rect 16396 8585 16405 8619
rect 16405 8585 16439 8619
rect 16439 8585 16448 8619
rect 16396 8576 16448 8585
rect 16856 8619 16908 8628
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 17500 8576 17552 8628
rect 3332 8440 3384 8492
rect 10140 8508 10192 8560
rect 10692 8551 10744 8560
rect 10692 8517 10701 8551
rect 10701 8517 10735 8551
rect 10735 8517 10744 8551
rect 10692 8508 10744 8517
rect 12164 8508 12216 8560
rect 14004 8508 14056 8560
rect 7104 8440 7156 8492
rect 3240 8372 3292 8424
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 2688 8304 2740 8356
rect 2872 8304 2924 8356
rect 5816 8347 5868 8356
rect 3240 8236 3292 8288
rect 4252 8279 4304 8288
rect 4252 8245 4261 8279
rect 4261 8245 4295 8279
rect 4295 8245 4304 8279
rect 4252 8236 4304 8245
rect 4712 8279 4764 8288
rect 4712 8245 4721 8279
rect 4721 8245 4755 8279
rect 4755 8245 4764 8279
rect 4712 8236 4764 8245
rect 5816 8313 5825 8347
rect 5825 8313 5859 8347
rect 5859 8313 5868 8347
rect 5816 8304 5868 8313
rect 6920 8304 6972 8356
rect 5356 8236 5408 8288
rect 7104 8236 7156 8288
rect 8944 8440 8996 8492
rect 8484 8304 8536 8356
rect 11888 8304 11940 8356
rect 14372 8440 14424 8492
rect 14280 8372 14332 8424
rect 17316 8304 17368 8356
rect 9588 8279 9640 8288
rect 9588 8245 9597 8279
rect 9597 8245 9631 8279
rect 9631 8245 9640 8279
rect 9588 8236 9640 8245
rect 11704 8236 11756 8288
rect 11980 8236 12032 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 2780 8032 2832 8084
rect 4252 8032 4304 8084
rect 5080 8032 5132 8084
rect 7288 8032 7340 8084
rect 7656 8032 7708 8084
rect 8208 8032 8260 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 8668 8032 8720 8084
rect 10324 8032 10376 8084
rect 12072 8075 12124 8084
rect 12072 8041 12081 8075
rect 12081 8041 12115 8075
rect 12115 8041 12124 8075
rect 12072 8032 12124 8041
rect 12992 8032 13044 8084
rect 13360 8032 13412 8084
rect 13544 8075 13596 8084
rect 13544 8041 13553 8075
rect 13553 8041 13587 8075
rect 13587 8041 13596 8075
rect 13544 8032 13596 8041
rect 13912 8075 13964 8084
rect 13912 8041 13921 8075
rect 13921 8041 13955 8075
rect 13955 8041 13964 8075
rect 13912 8032 13964 8041
rect 14280 8032 14332 8084
rect 16856 8032 16908 8084
rect 3148 7964 3200 8016
rect 3792 7964 3844 8016
rect 4068 7964 4120 8016
rect 2780 7896 2832 7948
rect 2964 7896 3016 7948
rect 4160 7896 4212 7948
rect 4712 7896 4764 7948
rect 5356 7939 5408 7948
rect 5356 7905 5390 7939
rect 5390 7905 5408 7939
rect 5356 7896 5408 7905
rect 6828 7896 6880 7948
rect 7104 7939 7156 7948
rect 7104 7905 7113 7939
rect 7113 7905 7147 7939
rect 7147 7905 7156 7939
rect 7104 7896 7156 7905
rect 7748 7896 7800 7948
rect 7840 7896 7892 7948
rect 12164 7896 12216 7948
rect 12716 7896 12768 7948
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 3792 7828 3844 7880
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 8208 7828 8260 7880
rect 10508 7828 10560 7880
rect 11888 7828 11940 7880
rect 11980 7828 12032 7880
rect 1124 7760 1176 7812
rect 3240 7760 3292 7812
rect 8944 7803 8996 7812
rect 8944 7769 8953 7803
rect 8953 7769 8987 7803
rect 8987 7769 8996 7803
rect 8944 7760 8996 7769
rect 10968 7760 11020 7812
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 3976 7692 4028 7744
rect 7012 7692 7064 7744
rect 8852 7692 8904 7744
rect 9956 7692 10008 7744
rect 15936 7760 15988 7812
rect 12900 7692 12952 7744
rect 15016 7735 15068 7744
rect 15016 7701 15025 7735
rect 15025 7701 15059 7735
rect 15059 7701 15068 7735
rect 15016 7692 15068 7701
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 1952 7488 2004 7540
rect 3792 7488 3844 7540
rect 2872 7352 2924 7404
rect 5080 7488 5132 7540
rect 7012 7488 7064 7540
rect 10508 7488 10560 7540
rect 11612 7488 11664 7540
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 12624 7488 12676 7540
rect 13176 7531 13228 7540
rect 13176 7497 13185 7531
rect 13185 7497 13219 7531
rect 13219 7497 13228 7531
rect 13176 7488 13228 7497
rect 13268 7488 13320 7540
rect 19524 7488 19576 7540
rect 12164 7420 12216 7472
rect 2504 7284 2556 7336
rect 2136 7259 2188 7268
rect 2136 7225 2145 7259
rect 2145 7225 2179 7259
rect 2179 7225 2188 7259
rect 2136 7216 2188 7225
rect 3332 7327 3384 7336
rect 3332 7293 3366 7327
rect 3366 7293 3384 7327
rect 3332 7284 3384 7293
rect 3240 7216 3292 7268
rect 5816 7352 5868 7404
rect 6828 7395 6880 7404
rect 5724 7284 5776 7336
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 10048 7352 10100 7404
rect 13452 7352 13504 7404
rect 15016 7352 15068 7404
rect 16672 7284 16724 7336
rect 7104 7259 7156 7268
rect 7104 7225 7138 7259
rect 7138 7225 7156 7259
rect 7104 7216 7156 7225
rect 7380 7216 7432 7268
rect 2872 7191 2924 7200
rect 2872 7157 2881 7191
rect 2881 7157 2915 7191
rect 2915 7157 2924 7191
rect 2872 7148 2924 7157
rect 5356 7148 5408 7200
rect 8300 7148 8352 7200
rect 8852 7191 8904 7200
rect 8852 7157 8861 7191
rect 8861 7157 8895 7191
rect 8895 7157 8904 7191
rect 8852 7148 8904 7157
rect 8944 7191 8996 7200
rect 8944 7157 8953 7191
rect 8953 7157 8987 7191
rect 8987 7157 8996 7191
rect 9864 7191 9916 7200
rect 8944 7148 8996 7157
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 4252 6944 4304 6996
rect 5540 6944 5592 6996
rect 5724 6987 5776 6996
rect 5724 6953 5733 6987
rect 5733 6953 5767 6987
rect 5767 6953 5776 6987
rect 5724 6944 5776 6953
rect 3332 6876 3384 6928
rect 1492 6808 1544 6860
rect 2044 6851 2096 6860
rect 2044 6817 2053 6851
rect 2053 6817 2087 6851
rect 2087 6817 2096 6851
rect 2044 6808 2096 6817
rect 2228 6808 2280 6860
rect 3056 6808 3108 6860
rect 4344 6876 4396 6928
rect 5080 6876 5132 6928
rect 6828 6919 6880 6928
rect 6828 6885 6837 6919
rect 6837 6885 6871 6919
rect 6871 6885 6880 6919
rect 6828 6876 6880 6885
rect 6000 6808 6052 6860
rect 7748 6944 7800 6996
rect 8300 6944 8352 6996
rect 10048 6944 10100 6996
rect 7104 6876 7156 6928
rect 7288 6808 7340 6860
rect 8208 6876 8260 6928
rect 8668 6851 8720 6860
rect 6644 6740 6696 6792
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 4160 6672 4212 6724
rect 8484 6740 8536 6792
rect 9036 6808 9088 6860
rect 9404 6808 9456 6860
rect 11980 6808 12032 6860
rect 12532 6808 12584 6860
rect 14188 6808 14240 6860
rect 19064 6851 19116 6860
rect 19064 6817 19073 6851
rect 19073 6817 19107 6851
rect 19107 6817 19116 6851
rect 19064 6808 19116 6817
rect 11796 6740 11848 6792
rect 8116 6672 8168 6724
rect 9864 6715 9916 6724
rect 9864 6681 9873 6715
rect 9873 6681 9907 6715
rect 9907 6681 9916 6715
rect 9864 6672 9916 6681
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 7840 6604 7892 6656
rect 19616 6672 19668 6724
rect 19892 6672 19944 6724
rect 10140 6604 10192 6656
rect 10692 6604 10744 6656
rect 11612 6604 11664 6656
rect 13544 6647 13596 6656
rect 13544 6613 13553 6647
rect 13553 6613 13587 6647
rect 13587 6613 13596 6647
rect 13544 6604 13596 6613
rect 20076 6604 20128 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 1860 6400 1912 6452
rect 2780 6400 2832 6452
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 5908 6400 5960 6452
rect 6920 6400 6972 6452
rect 1768 6332 1820 6384
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 5356 6332 5408 6384
rect 6828 6332 6880 6384
rect 7380 6332 7432 6384
rect 2964 6196 3016 6248
rect 8116 6400 8168 6452
rect 8668 6400 8720 6452
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 10692 6400 10744 6452
rect 12716 6443 12768 6452
rect 12716 6409 12725 6443
rect 12725 6409 12759 6443
rect 12759 6409 12768 6443
rect 12716 6400 12768 6409
rect 13544 6400 13596 6452
rect 19616 6443 19668 6452
rect 19616 6409 19625 6443
rect 19625 6409 19659 6443
rect 19659 6409 19668 6443
rect 19616 6400 19668 6409
rect 20720 6400 20772 6452
rect 7932 6332 7984 6384
rect 10140 6332 10192 6384
rect 13452 6332 13504 6384
rect 7748 6264 7800 6316
rect 8392 6264 8444 6316
rect 9312 6196 9364 6248
rect 11612 6196 11664 6248
rect 12164 6196 12216 6248
rect 6460 6128 6512 6180
rect 8484 6128 8536 6180
rect 4252 6060 4304 6112
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 7380 6060 7432 6112
rect 8300 6060 8352 6112
rect 19064 6103 19116 6112
rect 19064 6069 19073 6103
rect 19073 6069 19107 6103
rect 19107 6069 19116 6103
rect 19064 6060 19116 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 2780 5899 2832 5908
rect 2780 5865 2789 5899
rect 2789 5865 2823 5899
rect 2823 5865 2832 5899
rect 2780 5856 2832 5865
rect 2964 5856 3016 5908
rect 4160 5856 4212 5908
rect 4804 5856 4856 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 6184 5899 6236 5908
rect 6184 5865 6193 5899
rect 6193 5865 6227 5899
rect 6227 5865 6236 5899
rect 6184 5856 6236 5865
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 7288 5899 7340 5908
rect 7288 5865 7297 5899
rect 7297 5865 7331 5899
rect 7331 5865 7340 5899
rect 7288 5856 7340 5865
rect 8208 5856 8260 5908
rect 8760 5899 8812 5908
rect 8760 5865 8769 5899
rect 8769 5865 8803 5899
rect 8803 5865 8812 5899
rect 8760 5856 8812 5865
rect 10600 5856 10652 5908
rect 12716 5856 12768 5908
rect 21180 5856 21232 5908
rect 1400 5788 1452 5840
rect 3608 5788 3660 5840
rect 4068 5788 4120 5840
rect 12164 5788 12216 5840
rect 5264 5720 5316 5772
rect 7196 5720 7248 5772
rect 7748 5720 7800 5772
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 4896 5695 4948 5704
rect 4896 5661 4905 5695
rect 4905 5661 4939 5695
rect 4939 5661 4948 5695
rect 4896 5652 4948 5661
rect 7564 5652 7616 5704
rect 4804 5584 4856 5636
rect 5172 5584 5224 5636
rect 8668 5584 8720 5636
rect 5356 5516 5408 5568
rect 7104 5516 7156 5568
rect 9312 5516 9364 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 2412 5312 2464 5364
rect 2596 5355 2648 5364
rect 2596 5321 2605 5355
rect 2605 5321 2639 5355
rect 2639 5321 2648 5355
rect 2596 5312 2648 5321
rect 3424 5312 3476 5364
rect 4712 5312 4764 5364
rect 6092 5312 6144 5364
rect 7472 5312 7524 5364
rect 7748 5312 7800 5364
rect 8392 5312 8444 5364
rect 8576 5355 8628 5364
rect 8576 5321 8585 5355
rect 8585 5321 8619 5355
rect 8619 5321 8628 5355
rect 8576 5312 8628 5321
rect 9312 5355 9364 5364
rect 9312 5321 9321 5355
rect 9321 5321 9355 5355
rect 9355 5321 9364 5355
rect 9312 5312 9364 5321
rect 20904 5312 20956 5364
rect 3700 5244 3752 5296
rect 7564 5244 7616 5296
rect 3148 5176 3200 5228
rect 3240 5176 3292 5228
rect 7656 5176 7708 5228
rect 4068 5108 4120 5160
rect 3976 5040 4028 5092
rect 20260 5083 20312 5092
rect 20260 5049 20269 5083
rect 20269 5049 20303 5083
rect 20303 5049 20312 5083
rect 20260 5040 20312 5049
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2136 4768 2188 4820
rect 2504 4768 2556 4820
rect 2688 4768 2740 4820
rect 3240 4811 3292 4820
rect 3240 4777 3249 4811
rect 3249 4777 3283 4811
rect 3283 4777 3292 4811
rect 3240 4768 3292 4777
rect 6736 4768 6788 4820
rect 7748 4768 7800 4820
rect 8576 4768 8628 4820
rect 4068 4428 4120 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 8576 4224 8628 4276
rect 2964 4156 3016 4208
rect 1400 4088 1452 4140
rect 3240 4088 3292 4140
rect 4068 4088 4120 4140
rect 6736 4088 6788 4140
rect 5448 4020 5500 4072
rect 11152 4020 11204 4072
rect 3976 3952 4028 4004
rect 5356 3952 5408 4004
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 2964 3723 3016 3732
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 4068 3680 4120 3732
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
<< metal2 >>
rect 202 22000 258 22800
rect 570 22000 626 22800
rect 1030 22000 1086 22800
rect 1490 22000 1546 22800
rect 1950 22000 2006 22800
rect 2042 22536 2098 22545
rect 2042 22471 2098 22480
rect 216 18766 244 22000
rect 584 19122 612 22000
rect 938 19136 994 19145
rect 584 19094 938 19122
rect 938 19071 994 19080
rect 204 18760 256 18766
rect 204 18702 256 18708
rect 1044 17678 1072 22000
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1306 18864 1362 18873
rect 1412 18834 1440 19790
rect 1306 18799 1362 18808
rect 1400 18828 1452 18834
rect 1032 17672 1084 17678
rect 1032 17614 1084 17620
rect 1320 15094 1348 18799
rect 1400 18770 1452 18776
rect 1412 18465 1440 18770
rect 1504 18630 1532 22000
rect 1674 21176 1730 21185
rect 1674 21111 1730 21120
rect 1582 20632 1638 20641
rect 1582 20567 1638 20576
rect 1596 19174 1624 20567
rect 1688 20058 1716 21111
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1858 19272 1914 19281
rect 1858 19207 1914 19216
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1766 18592 1822 18601
rect 1766 18527 1822 18536
rect 1398 18456 1454 18465
rect 1398 18391 1454 18400
rect 1780 18222 1808 18527
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1492 17604 1544 17610
rect 1492 17546 1544 17552
rect 1504 17134 1532 17546
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 1504 16114 1532 17070
rect 1582 16552 1638 16561
rect 1582 16487 1638 16496
rect 1596 16250 1624 16487
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1308 15088 1360 15094
rect 1308 15030 1360 15036
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1412 13938 1440 14418
rect 1504 14414 1532 14894
rect 1492 14408 1544 14414
rect 1492 14350 1544 14356
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1596 13870 1624 15302
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 13462 1624 13806
rect 1584 13456 1636 13462
rect 1584 13398 1636 13404
rect 1688 13394 1716 17478
rect 1766 16960 1822 16969
rect 1766 16895 1822 16904
rect 1780 16794 1808 16895
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1766 13696 1822 13705
rect 1766 13631 1822 13640
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1412 12850 1440 13330
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1400 12708 1452 12714
rect 1400 12650 1452 12656
rect 1308 10600 1360 10606
rect 1308 10542 1360 10548
rect 1320 9353 1348 10542
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 1214 9208 1270 9217
rect 1214 9143 1270 9152
rect 1032 8900 1084 8906
rect 1032 8842 1084 8848
rect 1044 1057 1072 8842
rect 1124 7812 1176 7818
rect 1124 7754 1176 7760
rect 1030 1048 1086 1057
rect 1030 983 1086 992
rect 1136 649 1164 7754
rect 1228 2961 1256 9143
rect 1320 5658 1348 9279
rect 1412 5846 1440 12650
rect 1504 12238 1532 12718
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1504 6866 1532 10542
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1596 5914 1624 12786
rect 1780 12442 1808 13631
rect 1872 12986 1900 19207
rect 1964 18290 1992 22000
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1964 17921 1992 18022
rect 1950 17912 2006 17921
rect 1950 17847 2006 17856
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17377 1992 17478
rect 1950 17368 2006 17377
rect 1950 17303 2006 17312
rect 1950 15464 2006 15473
rect 1950 15399 2006 15408
rect 1964 14958 1992 15399
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 2056 14618 2084 22471
rect 2410 22000 2466 22800
rect 2870 22000 2926 22800
rect 3238 22128 3294 22137
rect 3238 22063 3294 22072
rect 2320 19984 2372 19990
rect 2320 19926 2372 19932
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 2240 19378 2268 19450
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2148 16250 2176 19110
rect 2240 18902 2268 19314
rect 2332 19242 2360 19926
rect 2320 19236 2372 19242
rect 2320 19178 2372 19184
rect 2228 18896 2280 18902
rect 2332 18873 2360 19178
rect 2228 18838 2280 18844
rect 2318 18864 2374 18873
rect 2318 18799 2374 18808
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2136 15972 2188 15978
rect 2136 15914 2188 15920
rect 2148 15366 2176 15914
rect 2240 15910 2268 18226
rect 2318 18048 2374 18057
rect 2318 17983 2374 17992
rect 2332 17202 2360 17983
rect 2424 17785 2452 22000
rect 2778 21584 2834 21593
rect 2778 21519 2834 21528
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2608 18204 2636 19246
rect 2686 19000 2742 19009
rect 2792 18970 2820 21519
rect 2884 20346 2912 22000
rect 3252 21706 3280 22063
rect 3330 22000 3386 22800
rect 3790 22000 3846 22800
rect 4250 22000 4306 22800
rect 4710 22000 4766 22800
rect 5170 22000 5226 22800
rect 5630 22000 5686 22800
rect 6090 22000 6146 22800
rect 6550 22000 6606 22800
rect 7010 22000 7066 22800
rect 7470 22000 7526 22800
rect 7930 22000 7986 22800
rect 8390 22000 8446 22800
rect 8850 22000 8906 22800
rect 9310 22000 9366 22800
rect 9770 22000 9826 22800
rect 10230 22000 10286 22800
rect 10690 22000 10746 22800
rect 11150 22000 11206 22800
rect 11610 22000 11666 22800
rect 11978 22000 12034 22800
rect 12438 22000 12494 22800
rect 12898 22000 12954 22800
rect 13358 22000 13414 22800
rect 13818 22000 13874 22800
rect 14278 22000 14334 22800
rect 14738 22000 14794 22800
rect 15198 22000 15254 22800
rect 15658 22000 15714 22800
rect 16118 22000 16174 22800
rect 16578 22000 16634 22800
rect 17038 22000 17094 22800
rect 17498 22000 17554 22800
rect 17958 22000 18014 22800
rect 18418 22000 18474 22800
rect 18878 22000 18934 22800
rect 19338 22000 19394 22800
rect 19798 22000 19854 22800
rect 20258 22000 20314 22800
rect 20718 22000 20774 22800
rect 21178 22000 21234 22800
rect 21638 22000 21694 22800
rect 22098 22000 22154 22800
rect 22558 22000 22614 22800
rect 3344 21842 3372 22000
rect 3344 21814 3740 21842
rect 3252 21678 3372 21706
rect 2884 20318 3188 20346
rect 2962 20224 3018 20233
rect 2962 20159 3018 20168
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 2884 18970 2912 19858
rect 2686 18935 2742 18944
rect 2780 18964 2832 18970
rect 2700 18834 2728 18935
rect 2780 18906 2832 18912
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2700 18358 2728 18566
rect 2688 18352 2740 18358
rect 2688 18294 2740 18300
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 2688 18216 2740 18222
rect 2608 18176 2688 18204
rect 2688 18158 2740 18164
rect 2410 17776 2466 17785
rect 2410 17711 2466 17720
rect 2700 17202 2728 18158
rect 2792 17882 2820 18255
rect 2870 17912 2926 17921
rect 2780 17876 2832 17882
rect 2870 17847 2926 17856
rect 2780 17818 2832 17824
rect 2884 17746 2912 17847
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2780 17672 2832 17678
rect 2778 17640 2780 17649
rect 2832 17640 2834 17649
rect 2778 17575 2834 17584
rect 2778 17504 2834 17513
rect 2778 17439 2834 17448
rect 2792 17338 2820 17439
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2332 16794 2360 17138
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2320 16652 2372 16658
rect 2372 16612 2452 16640
rect 2320 16594 2372 16600
rect 2424 16454 2452 16612
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 2228 15904 2280 15910
rect 2228 15846 2280 15852
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 2044 14612 2096 14618
rect 2044 14554 2096 14560
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1964 12374 1992 13330
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2056 12646 2084 12718
rect 2148 12714 2176 15302
rect 2332 15026 2360 16118
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2136 12708 2188 12714
rect 2136 12650 2188 12656
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1952 12368 2004 12374
rect 1952 12310 2004 12316
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1688 11558 1716 12242
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11286 1716 11494
rect 1676 11280 1728 11286
rect 1676 11222 1728 11228
rect 1780 10282 1808 12174
rect 2056 11336 2084 12582
rect 2240 12424 2268 14418
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 1688 10254 1808 10282
rect 1872 11308 2084 11336
rect 2148 12396 2268 12424
rect 1688 6458 1716 10254
rect 1768 10192 1820 10198
rect 1768 10134 1820 10140
rect 1780 9722 1808 10134
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1766 9616 1822 9625
rect 1766 9551 1822 9560
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1780 6390 1808 9551
rect 1872 6458 1900 11308
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1964 10470 1992 11154
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 7546 1992 10406
rect 2056 9761 2084 11086
rect 2042 9752 2098 9761
rect 2042 9687 2098 9696
rect 2148 9602 2176 12396
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2240 11529 2268 12242
rect 2226 11520 2282 11529
rect 2226 11455 2282 11464
rect 2240 11150 2268 11455
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2240 10266 2268 10950
rect 2332 10606 2360 14350
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2056 9574 2176 9602
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2056 6866 2084 9574
rect 2240 9178 2268 10066
rect 2332 9926 2360 10406
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2332 9058 2360 9862
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2240 9030 2360 9058
rect 2148 7274 2176 8978
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1400 5840 1452 5846
rect 1400 5782 1452 5788
rect 1320 5630 1440 5658
rect 1412 4146 1440 5630
rect 2148 4826 2176 7210
rect 2240 6866 2268 9030
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2332 5914 2360 7822
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2424 5370 2452 16390
rect 2700 16153 2728 17138
rect 2884 16590 2912 17682
rect 2976 16998 3004 20159
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 3068 18426 3096 18702
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3068 17882 3096 18362
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3054 17640 3110 17649
rect 3054 17575 3110 17584
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 3068 16726 3096 17575
rect 3160 17105 3188 20318
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 17338 3280 18566
rect 3344 17610 3372 21678
rect 3514 19816 3570 19825
rect 3514 19751 3570 19760
rect 3332 17604 3384 17610
rect 3332 17546 3384 17552
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3252 17134 3280 17274
rect 3240 17128 3292 17134
rect 3146 17096 3202 17105
rect 3240 17070 3292 17076
rect 3146 17031 3202 17040
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2686 16144 2742 16153
rect 2686 16079 2742 16088
rect 3054 16144 3110 16153
rect 3054 16079 3110 16088
rect 2700 16046 2728 16079
rect 2688 16040 2740 16046
rect 2964 16040 3016 16046
rect 2688 15982 2740 15988
rect 2778 16008 2834 16017
rect 2964 15982 3016 15988
rect 2778 15943 2834 15952
rect 2686 15056 2742 15065
rect 2686 14991 2742 15000
rect 2594 14920 2650 14929
rect 2594 14855 2596 14864
rect 2648 14855 2650 14864
rect 2596 14826 2648 14832
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2608 13870 2636 14282
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2516 11354 2544 11630
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2516 11014 2544 11154
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2516 10674 2544 10950
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2516 9722 2544 10202
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2516 9353 2544 9386
rect 2502 9344 2558 9353
rect 2502 9279 2558 9288
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2516 7342 2544 8910
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2516 4826 2544 7278
rect 2608 5370 2636 13806
rect 2700 11354 2728 14991
rect 2792 14074 2820 15943
rect 2976 15706 3004 15982
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2962 15600 3018 15609
rect 2962 15535 3018 15544
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2778 13968 2834 13977
rect 2778 13903 2834 13912
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2700 10305 2728 11086
rect 2686 10296 2742 10305
rect 2686 10231 2742 10240
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2700 9518 2728 10134
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2700 8362 2728 9454
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2686 8256 2742 8265
rect 2686 8191 2742 8200
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2700 4826 2728 8191
rect 2792 8090 2820 13903
rect 2884 13530 2912 14214
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2976 12442 3004 15535
rect 3068 14822 3096 16079
rect 3252 15706 3280 16594
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 3160 14958 3188 15506
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 3146 14648 3202 14657
rect 3146 14583 3202 14592
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2872 11688 2924 11694
rect 2924 11648 3004 11676
rect 2872 11630 2924 11636
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2884 9722 2912 10950
rect 2976 10198 3004 11648
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 3068 11150 3096 11562
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 3068 9994 3096 10474
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2792 6458 2820 7890
rect 2884 7410 2912 8298
rect 2976 7954 3004 8978
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7857 3004 7890
rect 2962 7848 3018 7857
rect 2962 7783 3018 7792
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2870 7304 2926 7313
rect 2870 7239 2926 7248
rect 2884 7206 2912 7239
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2792 5914 2820 6394
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 2884 3505 2912 7142
rect 2976 6254 3004 7686
rect 3068 6866 3096 9930
rect 3160 8838 3188 14583
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3344 14074 3372 14418
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3424 13320 3476 13326
rect 3528 13308 3556 19751
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3620 15473 3648 19654
rect 3712 18358 3740 21814
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 3606 15464 3662 15473
rect 3606 15399 3662 15408
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3620 14278 3648 14418
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3476 13280 3556 13308
rect 3424 13262 3476 13268
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 3252 11558 3280 12242
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3252 10470 3280 10610
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3252 9382 3280 10406
rect 3344 10062 3372 10406
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3252 8430 3280 9318
rect 3344 9110 3372 9998
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2976 5914 3004 6190
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 3160 5234 3188 7958
rect 3252 7818 3280 8230
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3344 7342 3372 8434
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 5234 3280 7210
rect 3344 6934 3372 7278
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3436 5370 3464 9658
rect 3528 9382 3556 10066
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 8634 3556 9318
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3620 5846 3648 14214
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3712 11642 3740 13806
rect 3804 12220 3832 22000
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4080 19922 4108 20334
rect 4264 20074 4292 22000
rect 4172 20046 4292 20074
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 19310 4108 19654
rect 4068 19304 4120 19310
rect 4066 19272 4068 19281
rect 4120 19272 4122 19281
rect 4066 19207 4122 19216
rect 4080 19181 4108 19207
rect 4066 18728 4122 18737
rect 4066 18663 4068 18672
rect 4120 18663 4122 18672
rect 4068 18634 4120 18640
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 4066 18592 4122 18601
rect 3988 18426 4016 18566
rect 4066 18527 4122 18536
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 4080 18154 4108 18527
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 17338 4108 17478
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4080 16250 4108 16526
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3988 15638 4016 15846
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 4080 15570 4108 16186
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3976 14340 4028 14346
rect 4080 14328 4108 14758
rect 4172 14618 4200 20046
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 4264 18290 4292 19858
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4434 19408 4490 19417
rect 4434 19343 4490 19352
rect 4448 19145 4476 19343
rect 4528 19168 4580 19174
rect 4434 19136 4490 19145
rect 4528 19110 4580 19116
rect 4434 19071 4490 19080
rect 4540 18766 4568 19110
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4264 17882 4292 18022
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4264 17066 4292 17614
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4356 16590 4384 16934
rect 4724 16794 4752 22000
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4908 19378 4936 19722
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4908 19174 4936 19314
rect 5000 19174 5028 19790
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4988 19168 5040 19174
rect 5092 19145 5120 19246
rect 4988 19110 5040 19116
rect 5078 19136 5134 19145
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4816 18086 4844 18702
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4908 18034 4936 19110
rect 5078 19071 5134 19080
rect 5184 18970 5212 22000
rect 5644 20058 5672 22000
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5354 19136 5410 19145
rect 5354 19071 5410 19080
rect 5262 19000 5318 19009
rect 5172 18964 5224 18970
rect 5262 18935 5318 18944
rect 5172 18906 5224 18912
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 5092 18358 5120 18770
rect 5184 18426 5212 18906
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5080 18352 5132 18358
rect 5080 18294 5132 18300
rect 5276 18193 5304 18935
rect 5368 18766 5396 19071
rect 5552 18958 5856 18986
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5262 18184 5318 18193
rect 5262 18119 5318 18128
rect 5172 18080 5224 18086
rect 4908 18006 5028 18034
rect 5172 18022 5224 18028
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4816 17134 4844 17614
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4356 16436 4384 16526
rect 4264 16408 4384 16436
rect 4264 16046 4292 16408
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4724 16250 4752 16730
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4816 16153 4844 16390
rect 4802 16144 4858 16153
rect 4802 16079 4858 16088
rect 4816 16046 4844 16079
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4724 15162 4752 15642
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4816 14958 4844 15982
rect 4804 14952 4856 14958
rect 4896 14952 4948 14958
rect 4804 14894 4856 14900
rect 4894 14920 4896 14929
rect 4948 14920 4950 14929
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4028 14300 4108 14328
rect 3976 14282 4028 14288
rect 4080 13954 4108 14300
rect 4172 14074 4200 14350
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4080 13926 4200 13954
rect 4172 13870 4200 13926
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4724 13530 4752 14418
rect 4816 14414 4844 14894
rect 4894 14855 4950 14864
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4816 13802 4844 14350
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4172 12850 4200 13330
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4068 12368 4120 12374
rect 4066 12336 4068 12345
rect 4120 12336 4122 12345
rect 4066 12271 4122 12280
rect 4068 12232 4120 12238
rect 3804 12192 3924 12220
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11830 3832 12038
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3712 11614 3832 11642
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3608 5840 3660 5846
rect 3608 5782 3660 5788
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3712 5302 3740 11494
rect 3804 8022 3832 11614
rect 3896 10674 3924 12192
rect 4264 12186 4292 12786
rect 4724 12306 4752 12922
rect 4816 12714 4844 13194
rect 4908 12986 4936 13262
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4120 12180 4292 12186
rect 4068 12174 4292 12180
rect 4080 12158 4292 12174
rect 4066 11792 4122 11801
rect 4066 11727 4122 11736
rect 4080 11626 4108 11727
rect 4172 11694 4200 12158
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4908 11558 4936 11834
rect 4436 11552 4488 11558
rect 4434 11520 4436 11529
rect 4804 11552 4856 11558
rect 4488 11520 4490 11529
rect 4804 11494 4856 11500
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4434 11455 4490 11464
rect 4066 11384 4122 11393
rect 4066 11319 4122 11328
rect 4528 11348 4580 11354
rect 4080 11082 4108 11319
rect 4816 11336 4844 11494
rect 4580 11308 4844 11336
rect 4528 11290 4580 11296
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3988 10470 4016 10950
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4066 10840 4122 10849
rect 4388 10832 4684 10852
rect 4066 10775 4068 10784
rect 4120 10775 4122 10784
rect 4068 10746 4120 10752
rect 4724 10538 4752 11154
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 4066 10432 4122 10441
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 8634 3924 9862
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3792 7880 3844 7886
rect 3988 7834 4016 10406
rect 4066 10367 4122 10376
rect 4080 9722 4108 10367
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4068 9580 4120 9586
rect 4120 9540 4292 9568
rect 4068 9522 4120 9528
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 8906 4108 9318
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4172 8537 4200 9046
rect 4264 8838 4292 9540
rect 4724 9382 4752 10474
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 8838 4752 9318
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4264 8634 4292 8774
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4158 8528 4214 8537
rect 4158 8463 4214 8472
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4264 8090 4292 8230
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 3792 7822 3844 7828
rect 3804 7546 3832 7822
rect 3896 7806 4016 7834
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3252 4826 3280 5170
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2976 3738 3004 4150
rect 3252 4146 3280 4762
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2870 3496 2926 3505
rect 2870 3431 2926 3440
rect 1214 2952 1270 2961
rect 1214 2887 1270 2896
rect 1122 640 1178 649
rect 1122 575 1178 584
rect 3896 241 3924 7806
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 6322 4016 7686
rect 4080 7585 4108 7958
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 4172 6730 4200 7890
rect 4264 7002 4292 8026
rect 4724 7954 4752 8230
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4342 7304 4398 7313
rect 4342 7239 4398 7248
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4356 6934 4384 7239
rect 4344 6928 4396 6934
rect 4264 6876 4344 6882
rect 4264 6870 4396 6876
rect 4264 6854 4384 6870
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4172 5914 4200 6666
rect 4264 6118 4292 6854
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4068 5840 4120 5846
rect 4066 5808 4068 5817
rect 4120 5808 4122 5817
rect 4066 5743 4122 5752
rect 3974 5264 4030 5273
rect 3974 5199 4030 5208
rect 3988 5098 4016 5199
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 4080 4865 4108 5102
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4080 4146 4108 4422
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3988 3913 4016 3946
rect 3974 3904 4030 3913
rect 3974 3839 4030 3848
rect 4080 3738 4108 4082
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4264 2553 4292 6054
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4724 5370 4752 7890
rect 4816 5914 4844 11308
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4908 5710 4936 11494
rect 5000 9058 5028 18006
rect 5184 17678 5212 18022
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5184 16454 5212 17614
rect 5276 16998 5304 18119
rect 5368 18086 5396 18702
rect 5446 18456 5502 18465
rect 5446 18391 5502 18400
rect 5460 18290 5488 18391
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5552 18222 5580 18958
rect 5828 18902 5856 18958
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5644 18714 5672 18770
rect 5644 18686 6040 18714
rect 5724 18624 5776 18630
rect 5776 18601 5856 18612
rect 5776 18592 5870 18601
rect 5776 18584 5814 18592
rect 5724 18566 5776 18572
rect 5814 18527 5870 18536
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5828 18086 5856 18527
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5920 17898 5948 18226
rect 5644 17882 5948 17898
rect 5632 17876 5948 17882
rect 5684 17870 5948 17876
rect 5632 17818 5684 17824
rect 5920 17270 5948 17870
rect 6012 17542 6040 18686
rect 6104 18154 6132 22000
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6090 17912 6146 17921
rect 6090 17847 6146 17856
rect 6104 17814 6132 17847
rect 6092 17808 6144 17814
rect 6092 17750 6144 17756
rect 6288 17610 6316 18362
rect 6276 17604 6328 17610
rect 6276 17546 6328 17552
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5276 15706 5304 16526
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5736 15366 5764 16594
rect 5920 16250 5948 17206
rect 6288 16998 6316 17546
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 6196 15978 6224 16390
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5184 12986 5212 13330
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5092 11540 5120 12582
rect 5276 11694 5304 13942
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5264 11552 5316 11558
rect 5092 11512 5264 11540
rect 5264 11494 5316 11500
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5184 10810 5212 11290
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5092 9382 5120 9590
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5092 9217 5120 9318
rect 5078 9208 5134 9217
rect 5078 9143 5134 9152
rect 5000 9030 5212 9058
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 5000 6916 5028 8842
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 8090 5120 8774
rect 5184 8634 5212 9030
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5092 7546 5120 7822
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5080 6928 5132 6934
rect 5000 6888 5080 6916
rect 5080 6870 5132 6876
rect 5092 6118 5120 6870
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4250 2544 4306 2553
rect 4250 2479 4306 2488
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4816 2009 4844 5578
rect 4802 2000 4858 2009
rect 4802 1935 4858 1944
rect 5092 1601 5120 6054
rect 5184 5642 5212 8570
rect 5276 5778 5304 11494
rect 5368 9042 5396 13466
rect 5538 13288 5594 13297
rect 5538 13223 5594 13232
rect 5552 12918 5580 13223
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5460 11354 5488 12242
rect 5552 12238 5580 12650
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 11234 5580 11630
rect 5460 11206 5580 11234
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8294 5396 8774
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5368 7206 5396 7890
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 6662 5396 7142
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6390 5396 6598
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 4010 5396 5510
rect 5460 4078 5488 11206
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5552 10062 5580 10542
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5552 6458 5580 6938
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5644 5914 5672 15302
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 5736 14074 5764 14486
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11694 5764 12106
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5736 10470 5764 10610
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10198 5764 10406
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5736 9586 5764 10134
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 9178 5764 9522
rect 5828 9450 5856 15506
rect 6092 15496 6144 15502
rect 6196 15484 6224 15914
rect 6380 15502 6408 16934
rect 6564 15706 6592 22000
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6748 19242 6776 19654
rect 6736 19236 6788 19242
rect 6736 19178 6788 19184
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6656 18290 6684 19110
rect 6748 18970 6776 19178
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 7024 18034 7052 22000
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7116 18057 7144 19654
rect 7208 18154 7236 20198
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 6840 18006 7052 18034
rect 7102 18048 7158 18057
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6656 17202 6684 17478
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6656 16697 6684 16730
rect 6642 16688 6698 16697
rect 6642 16623 6644 16632
rect 6696 16623 6698 16632
rect 6644 16594 6696 16600
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6144 15456 6224 15484
rect 6092 15438 6144 15444
rect 6196 15162 6224 15456
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6380 14958 6408 15438
rect 6564 15162 6592 15642
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6656 15042 6684 15302
rect 6564 15014 6684 15042
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5814 8392 5870 8401
rect 5814 8327 5816 8336
rect 5868 8327 5870 8336
rect 5816 8298 5868 8304
rect 5814 8120 5870 8129
rect 5814 8055 5870 8064
rect 5828 7410 5856 8055
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5736 7002 5764 7278
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5920 6458 5948 13806
rect 6104 13802 6132 14214
rect 6288 13938 6316 14282
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6288 13172 6316 13874
rect 6380 13326 6408 14894
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6368 13184 6420 13190
rect 6288 13144 6368 13172
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6012 10690 6040 11154
rect 6104 10810 6132 13126
rect 6288 12442 6316 13144
rect 6368 13126 6420 13132
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6184 12300 6236 12306
rect 6288 12288 6316 12378
rect 6236 12260 6316 12288
rect 6184 12242 6236 12248
rect 6380 12220 6408 12378
rect 6288 12192 6408 12220
rect 6288 11558 6316 12192
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11218 6316 11494
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6012 10662 6132 10690
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 6866 6040 10066
rect 6104 9926 6132 10662
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6104 6361 6132 9862
rect 6196 9382 6224 10202
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6090 6352 6146 6361
rect 6090 6287 6146 6296
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 6104 5370 6132 6287
rect 6196 5914 6224 9318
rect 6288 8945 6316 11154
rect 6380 9178 6408 11698
rect 6472 11150 6500 11698
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6564 9654 6592 15014
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6656 13326 6684 14350
rect 6644 13320 6696 13326
rect 6696 13280 6776 13308
rect 6644 13262 6696 13268
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6656 10742 6684 11018
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6552 9648 6604 9654
rect 6604 9608 6684 9636
rect 6552 9590 6604 9596
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6274 8936 6330 8945
rect 6274 8871 6330 8880
rect 6288 8838 6316 8871
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6472 6186 6500 9386
rect 6564 9382 6592 9454
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 6564 5914 6592 9318
rect 6656 6798 6684 9608
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6748 4826 6776 13280
rect 6840 11898 6868 18006
rect 7102 17983 7158 17992
rect 7300 17649 7328 19654
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7392 18154 7420 18702
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7286 17640 7342 17649
rect 7286 17575 7288 17584
rect 7340 17575 7342 17584
rect 7288 17546 7340 17552
rect 7300 17515 7328 17546
rect 7484 17218 7512 22000
rect 7944 20346 7972 22000
rect 7760 20318 7972 20346
rect 8208 20324 8260 20330
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7668 18834 7696 19246
rect 7656 18828 7708 18834
rect 7656 18770 7708 18776
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7576 18086 7604 18702
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7024 17190 7512 17218
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6932 15706 6960 16662
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6932 14074 6960 14418
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 7024 11694 7052 17190
rect 7576 17134 7604 17818
rect 7668 17746 7696 18770
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7116 16046 7144 17070
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7300 15484 7328 16390
rect 7392 16046 7420 16934
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7484 15910 7512 16526
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7484 15502 7512 15846
rect 7380 15496 7432 15502
rect 7300 15456 7380 15484
rect 7380 15438 7432 15444
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7208 13530 7236 13806
rect 7300 13530 7328 14894
rect 7392 14550 7420 15438
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7484 14482 7512 15438
rect 7576 15366 7604 16730
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7668 15094 7696 16594
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 13938 7420 14214
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7392 13394 7420 13874
rect 7576 13870 7604 14758
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7208 11558 7236 12582
rect 7576 12306 7604 12718
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7668 12186 7696 15030
rect 7760 14618 7788 20318
rect 8208 20266 8260 20272
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 8220 19174 8248 20266
rect 8404 20210 8432 22000
rect 8312 20182 8432 20210
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8024 18896 8076 18902
rect 8024 18838 8076 18844
rect 8036 18290 8064 18838
rect 8220 18714 8248 19110
rect 8128 18686 8248 18714
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8128 18154 8156 18686
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18290 8248 18566
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8116 18148 8168 18154
rect 8116 18090 8168 18096
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17882 8248 18226
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8220 16590 8248 16934
rect 8312 16794 8340 20182
rect 8864 20058 8892 22000
rect 9324 20058 9352 22000
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 8404 19378 8432 19994
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8484 18352 8536 18358
rect 8484 18294 8536 18300
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8404 17882 8432 18226
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8496 17746 8524 18294
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8312 16250 8340 16730
rect 8496 16454 8524 17138
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8496 16046 8524 16390
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7944 15162 7972 15506
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 8496 14958 8524 15982
rect 8588 15706 8616 19654
rect 8772 19174 8800 19654
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8772 18902 8800 19110
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 8666 18592 8722 18601
rect 8666 18527 8722 18536
rect 8680 17746 8708 18527
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8772 17626 8800 18838
rect 8956 18154 8984 19110
rect 9140 18222 9168 19790
rect 9324 19378 9352 19994
rect 9692 19922 9720 19994
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9312 19236 9364 19242
rect 9312 19178 9364 19184
rect 9324 18902 9352 19178
rect 9312 18896 9364 18902
rect 9312 18838 9364 18844
rect 9416 18358 9444 19654
rect 9680 19440 9732 19446
rect 9600 19388 9680 19394
rect 9600 19382 9732 19388
rect 9600 19366 9720 19382
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9404 18352 9456 18358
rect 9404 18294 9456 18300
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 9140 17882 9168 18158
rect 9128 17876 9180 17882
rect 9312 17876 9364 17882
rect 9128 17818 9180 17824
rect 9232 17836 9312 17864
rect 8772 17598 9076 17626
rect 8758 16688 8814 16697
rect 8758 16623 8760 16632
rect 8812 16623 8814 16632
rect 8760 16594 8812 16600
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8574 15464 8630 15473
rect 8574 15399 8576 15408
rect 8628 15399 8630 15408
rect 8576 15370 8628 15376
rect 8956 15162 8984 15506
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8850 14920 8906 14929
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7760 13734 7788 14554
rect 8496 13870 8524 14894
rect 8850 14855 8852 14864
rect 8904 14855 8906 14864
rect 8852 14826 8904 14832
rect 8956 14618 8984 15098
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 13870 8708 14214
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8220 12306 8248 13466
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7576 12158 7696 12186
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7392 11762 7420 12038
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7208 11354 7236 11494
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6828 10668 6880 10674
rect 6932 10656 6960 10950
rect 6880 10628 6960 10656
rect 6828 10610 6880 10616
rect 7024 10470 7052 11086
rect 7208 10713 7236 11290
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7300 10849 7328 11154
rect 7286 10840 7342 10849
rect 7286 10775 7342 10784
rect 7194 10704 7250 10713
rect 7194 10639 7250 10648
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6840 9636 6868 10066
rect 6932 9926 6960 10066
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6920 9648 6972 9654
rect 6840 9608 6920 9636
rect 6920 9590 6972 9596
rect 6920 9376 6972 9382
rect 6840 9336 6920 9364
rect 6840 9042 6868 9336
rect 6920 9318 6972 9324
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8634 6960 8910
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7024 8378 7052 10406
rect 7116 9994 7144 10474
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7116 9586 7144 9930
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7116 8498 7144 9522
rect 7208 9518 7236 9862
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7208 9178 7236 9454
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7300 9058 7328 10775
rect 7392 9178 7420 11698
rect 7484 10130 7512 12038
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7472 9512 7524 9518
rect 7470 9480 7472 9489
rect 7524 9480 7526 9489
rect 7470 9415 7526 9424
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7300 9030 7512 9058
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7288 8424 7340 8430
rect 6920 8356 6972 8362
rect 7024 8350 7236 8378
rect 7340 8384 7420 8412
rect 7288 8366 7340 8372
rect 6920 8298 6972 8304
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6840 7410 6868 7890
rect 6932 7528 6960 8298
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7116 7954 7144 8230
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7012 7744 7064 7750
rect 7064 7704 7144 7732
rect 7012 7686 7064 7692
rect 7012 7540 7064 7546
rect 6932 7500 7012 7528
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6840 6390 6868 6870
rect 6932 6458 6960 7500
rect 7012 7482 7064 7488
rect 7116 7274 7144 7704
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7116 6934 7144 7210
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 7116 5574 7144 6598
rect 7208 5778 7236 8350
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7300 6866 7328 8026
rect 7392 7274 7420 8384
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6066 7328 6598
rect 7392 6390 7420 7210
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7380 6112 7432 6118
rect 7300 6060 7380 6066
rect 7300 6054 7432 6060
rect 7300 6038 7420 6054
rect 7300 5914 7328 6038
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7484 5370 7512 9030
rect 7576 5710 7604 12158
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11694 7696 12038
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11218 7696 11494
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7668 9926 7696 11154
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7668 9586 7696 9862
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7760 9194 7788 12242
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7852 11762 7880 12174
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 11014 8248 11154
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10742 8248 10950
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7668 9166 7788 9194
rect 7668 8090 7696 9166
rect 8220 8514 8248 9522
rect 8496 9058 8524 13806
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8588 12306 8616 12582
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8680 12238 8708 13126
rect 8772 12753 8800 13126
rect 8758 12744 8814 12753
rect 8758 12679 8814 12688
rect 8864 12442 8892 13330
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8588 10810 8616 11018
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9178 8616 9998
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8496 9030 8616 9058
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 7944 8486 8248 8514
rect 7944 8430 7972 8486
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 8220 8242 8248 8486
rect 8496 8362 8524 8910
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8220 8214 8432 8242
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7576 5302 7604 5646
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7668 5234 7696 8026
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7760 7002 7788 7890
rect 7852 7449 7880 7890
rect 8220 7886 8248 8026
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 7838 7440 7894 7449
rect 7838 7375 7894 7384
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8312 7002 8340 7142
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 7760 6322 7788 6938
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7760 5778 7788 6258
rect 7852 6225 7880 6598
rect 8128 6458 8156 6666
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7932 6384 7984 6390
rect 7930 6352 7932 6361
rect 7984 6352 7986 6361
rect 7930 6287 7986 6296
rect 7838 6216 7894 6225
rect 7838 6151 7894 6160
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8220 5914 8248 6870
rect 8298 6760 8354 6769
rect 8298 6695 8354 6704
rect 8312 6118 8340 6695
rect 8404 6322 8432 8214
rect 8496 8090 8524 8298
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 8404 5370 8432 6258
rect 8496 6186 8524 6734
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 8588 5370 8616 9030
rect 8680 8090 8708 12174
rect 8864 11286 8892 12174
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8956 11626 8984 12038
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8956 11354 8984 11562
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8758 10840 8814 10849
rect 8758 10775 8760 10784
rect 8812 10775 8814 10784
rect 8760 10746 8812 10752
rect 8956 10742 8984 10950
rect 8944 10736 8996 10742
rect 8850 10704 8906 10713
rect 8944 10678 8996 10684
rect 8850 10639 8906 10648
rect 8864 10606 8892 10639
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8864 10130 8892 10542
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8772 8838 8800 10066
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8680 6458 8708 6802
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8680 5642 8708 6394
rect 8772 5914 8800 8774
rect 8864 7750 8892 10066
rect 8942 9072 8998 9081
rect 9048 9042 9076 17598
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 15978 9168 16390
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9140 15502 9168 15914
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 14822 9168 15438
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9140 14550 9168 14758
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9232 12986 9260 17836
rect 9312 17818 9364 17824
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9324 16454 9352 17546
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9416 16794 9444 16934
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9402 14920 9458 14929
rect 9312 14884 9364 14890
rect 9402 14855 9404 14864
rect 9312 14826 9364 14832
rect 9456 14855 9458 14864
rect 9404 14826 9456 14832
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9324 10033 9352 14826
rect 9508 13546 9536 19246
rect 9600 18766 9628 19366
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9600 18222 9628 18702
rect 9692 18630 9720 19178
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9692 18290 9720 18566
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9600 18086 9628 18158
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9600 17202 9628 18022
rect 9692 17882 9720 18022
rect 9784 17882 9812 22000
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9876 19378 9904 19722
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9876 18902 9904 19314
rect 10152 19242 10180 19654
rect 10140 19236 10192 19242
rect 10140 19178 10192 19184
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9586 17096 9642 17105
rect 9586 17031 9642 17040
rect 9600 15978 9628 17031
rect 9956 16720 10008 16726
rect 9954 16688 9956 16697
rect 10008 16688 10010 16697
rect 9954 16623 10010 16632
rect 9956 16448 10008 16454
rect 10060 16436 10088 17682
rect 10008 16408 10088 16436
rect 9956 16390 10008 16396
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9416 13518 9536 13546
rect 9416 11354 9444 13518
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9508 12918 9536 13330
rect 9600 12986 9628 13806
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9692 13326 9720 13670
rect 9784 13530 9812 13738
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9508 11830 9536 12242
rect 9600 12238 9628 12922
rect 9692 12782 9720 13262
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9692 11898 9720 12718
rect 9784 12442 9812 13466
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9416 10606 9444 11290
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9876 10470 9904 10950
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9310 10024 9366 10033
rect 9310 9959 9366 9968
rect 9692 9450 9812 9466
rect 9680 9444 9812 9450
rect 9732 9438 9812 9444
rect 9680 9386 9732 9392
rect 9496 9376 9548 9382
rect 9588 9376 9640 9382
rect 9548 9336 9588 9364
rect 9496 9318 9548 9324
rect 9588 9318 9640 9324
rect 8942 9007 8998 9016
rect 9036 9036 9088 9042
rect 8956 8498 8984 9007
rect 9036 8978 9088 8984
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9218 8936 9274 8945
rect 9218 8871 9220 8880
rect 9272 8871 9274 8880
rect 9220 8842 9272 8848
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 9600 8294 9628 8978
rect 9680 8968 9732 8974
rect 9784 8956 9812 9438
rect 9876 9382 9904 10406
rect 9968 9654 9996 16390
rect 10244 15706 10272 22000
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10322 19408 10378 19417
rect 10322 19343 10378 19352
rect 10336 19145 10364 19343
rect 10322 19136 10378 19145
rect 10322 19071 10378 19080
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10152 14890 10180 15438
rect 10244 15162 10272 15642
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10152 14618 10180 14826
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10152 14074 10180 14554
rect 10336 14482 10364 18906
rect 10428 17610 10456 19654
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10416 17604 10468 17610
rect 10416 17546 10468 17552
rect 10428 16794 10456 17546
rect 10520 16998 10548 18770
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10612 17202 10640 17614
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10612 16250 10640 17138
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10520 15162 10548 15506
rect 10612 15502 10640 15982
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10612 13870 10640 15438
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10152 12850 10180 13262
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10060 11694 10088 12174
rect 10152 11898 10180 12242
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 10130 10088 11494
rect 10152 11354 10180 11834
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 9178 10088 9318
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9732 8928 9812 8956
rect 9680 8910 9732 8916
rect 9692 8634 9720 8910
rect 10152 8838 10180 9590
rect 10336 9382 10364 10202
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 10152 8566 10180 8774
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8864 7206 8892 7686
rect 8956 7206 8984 7754
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 9048 6866 9076 7346
rect 9600 7313 9628 8230
rect 10336 8090 10364 9318
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9968 7410 9996 7686
rect 10520 7546 10548 7822
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9586 7304 9642 7313
rect 9586 7239 9642 7248
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9416 6458 9444 6802
rect 9876 6730 9904 7142
rect 10060 7002 10088 7346
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 10152 6390 10180 6598
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 9324 5574 9352 6190
rect 10612 5914 10640 13806
rect 10704 13802 10732 22000
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 10782 18456 10838 18465
rect 10888 18426 10916 18634
rect 10980 18426 11008 18838
rect 10782 18391 10838 18400
rect 10876 18420 10928 18426
rect 10796 18358 10824 18391
rect 10876 18362 10928 18368
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10888 18086 10916 18226
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 17338 11008 18022
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10980 16794 11008 17274
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10980 16590 11008 16730
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 11072 15366 11100 19926
rect 11164 19310 11192 22000
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 11624 19009 11652 22000
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11610 19000 11666 19009
rect 11610 18935 11666 18944
rect 11702 18864 11758 18873
rect 11612 18828 11664 18834
rect 11702 18799 11758 18808
rect 11612 18770 11664 18776
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11164 17785 11192 17818
rect 11150 17776 11206 17785
rect 11150 17711 11206 17720
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11164 15162 11192 17711
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11624 16794 11652 18770
rect 11716 18601 11744 18799
rect 11702 18592 11758 18601
rect 11702 18527 11758 18536
rect 11808 17762 11836 19654
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11900 19009 11928 19178
rect 11886 19000 11942 19009
rect 11886 18935 11942 18944
rect 11886 18864 11942 18873
rect 11886 18799 11942 18808
rect 11900 18329 11928 18799
rect 11886 18320 11942 18329
rect 11886 18255 11942 18264
rect 11716 17746 11836 17762
rect 11704 17740 11836 17746
rect 11756 17734 11836 17740
rect 11888 17740 11940 17746
rect 11704 17682 11756 17688
rect 11888 17682 11940 17688
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11624 16164 11652 16730
rect 11716 16522 11744 17478
rect 11808 17218 11836 17614
rect 11900 17542 11928 17682
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11900 17338 11928 17478
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11808 17190 11928 17218
rect 11900 17134 11928 17190
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11794 16960 11850 16969
rect 11794 16895 11850 16904
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11716 16250 11744 16458
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11532 16136 11652 16164
rect 11532 15450 11560 16136
rect 11716 15586 11744 16186
rect 11624 15570 11744 15586
rect 11612 15564 11744 15570
rect 11664 15558 11744 15564
rect 11612 15506 11664 15512
rect 11532 15422 11652 15450
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 10874 14376 10930 14385
rect 10874 14311 10930 14320
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10704 11150 10732 11494
rect 10888 11354 10916 14311
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11072 12322 11100 12378
rect 10980 12294 11100 12322
rect 10876 11348 10928 11354
rect 10796 11308 10876 11336
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10704 10130 10732 11086
rect 10796 10538 10824 11308
rect 10876 11290 10928 11296
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10704 8974 10732 10066
rect 10888 9518 10916 10610
rect 10980 10452 11008 12294
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 11694 11100 12174
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 10606 11100 11154
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10980 10424 11100 10452
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9586 11008 9862
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10704 8566 10732 8910
rect 10796 8906 10824 9318
rect 10980 9178 11008 9522
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10980 8634 11008 9114
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 11072 7834 11100 10424
rect 11164 8634 11192 13806
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11518 10568 11574 10577
rect 11518 10503 11520 10512
rect 11572 10503 11574 10512
rect 11520 10474 11572 10480
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11532 9178 11560 9454
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10980 7818 11100 7834
rect 10968 7812 11100 7818
rect 11020 7806 11100 7812
rect 10968 7754 11020 7760
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11624 7546 11652 15422
rect 11704 14816 11756 14822
rect 11808 14804 11836 16895
rect 11900 16182 11928 17070
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11756 14776 11836 14804
rect 11704 14758 11756 14764
rect 11716 14414 11744 14758
rect 11704 14408 11756 14414
rect 11888 14408 11940 14414
rect 11704 14350 11756 14356
rect 11886 14376 11888 14385
rect 11940 14376 11942 14385
rect 11886 14311 11942 14320
rect 11992 13818 12020 22000
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12084 15858 12112 19246
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12176 18329 12204 18770
rect 12348 18352 12400 18358
rect 12162 18320 12218 18329
rect 12348 18294 12400 18300
rect 12162 18255 12218 18264
rect 12360 17785 12388 18294
rect 12452 18057 12480 22000
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12636 19718 12664 19790
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12530 19136 12586 19145
rect 12530 19071 12586 19080
rect 12438 18048 12494 18057
rect 12438 17983 12494 17992
rect 12346 17776 12402 17785
rect 12346 17711 12402 17720
rect 12360 16969 12388 17711
rect 12346 16960 12402 16969
rect 12346 16895 12402 16904
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12360 16658 12388 16730
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12176 16250 12204 16390
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12084 15830 12204 15858
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 11900 13790 12020 13818
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11808 13025 11836 13194
rect 11794 13016 11850 13025
rect 11794 12951 11796 12960
rect 11848 12951 11850 12960
rect 11796 12922 11848 12928
rect 11808 12891 11836 12922
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11716 12306 11744 12582
rect 11808 12322 11836 12786
rect 11900 12442 11928 13790
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11992 13258 12020 13670
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 11992 12714 12020 13194
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11704 12300 11756 12306
rect 11808 12294 11928 12322
rect 11704 12242 11756 12248
rect 11716 11898 11744 12242
rect 11796 12096 11848 12102
rect 11900 12073 11928 12294
rect 11796 12038 11848 12044
rect 11886 12064 11942 12073
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11716 10606 11744 11834
rect 11808 11286 11836 12038
rect 11886 11999 11942 12008
rect 11900 11830 11928 11999
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11716 10130 11744 10542
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11702 10024 11758 10033
rect 11702 9959 11758 9968
rect 11716 8294 11744 9959
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11808 6798 11836 11222
rect 11900 8362 11928 11494
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11992 10130 12020 10610
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11992 9926 12020 10066
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 8838 12020 9862
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8634 12020 8774
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11900 7886 11928 8298
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11992 7886 12020 8230
rect 12084 8090 12112 15642
rect 12176 11937 12204 15830
rect 12360 15706 12388 16594
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12360 15026 12388 15302
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12360 14482 12388 14962
rect 12544 14906 12572 19071
rect 12636 16572 12664 19654
rect 12912 19174 12940 22000
rect 13372 20058 13400 22000
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12912 18086 12940 18770
rect 13004 18465 13032 19246
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 12990 18456 13046 18465
rect 12990 18391 13046 18400
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12820 17882 12848 18022
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12728 17762 12756 17818
rect 12728 17734 13032 17762
rect 13004 17678 13032 17734
rect 12992 17672 13044 17678
rect 13280 17649 13308 18770
rect 13372 18766 13400 19858
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13648 18970 13676 19246
rect 13832 19156 13860 22000
rect 14292 20058 14320 22000
rect 14752 20618 14780 22000
rect 14752 20590 15056 20618
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14096 19304 14148 19310
rect 14280 19304 14332 19310
rect 14096 19246 14148 19252
rect 14200 19264 14280 19292
rect 13912 19168 13964 19174
rect 13726 19136 13782 19145
rect 13832 19128 13912 19156
rect 13912 19110 13964 19116
rect 13726 19071 13782 19080
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13740 18426 13768 19071
rect 14016 18902 14044 19246
rect 14108 19145 14136 19246
rect 14094 19136 14150 19145
rect 14094 19071 14150 19080
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 14108 18834 14136 19071
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 12992 17614 13044 17620
rect 13266 17640 13322 17649
rect 13266 17575 13322 17584
rect 13360 17604 13412 17610
rect 12716 16584 12768 16590
rect 12636 16544 12716 16572
rect 12716 16526 12768 16532
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12452 14878 12572 14906
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12360 13870 12388 14418
rect 12452 14414 12480 14878
rect 12636 14822 12664 16390
rect 12728 16046 12756 16526
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12728 15026 12756 15982
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12820 14958 12848 15846
rect 13004 15502 13032 16050
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 12992 15496 13044 15502
rect 12990 15464 12992 15473
rect 13044 15464 13046 15473
rect 12990 15399 13046 15408
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12440 14408 12492 14414
rect 12438 14376 12440 14385
rect 12492 14376 12494 14385
rect 12438 14311 12494 14320
rect 12438 14240 12494 14249
rect 12438 14175 12494 14184
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12452 12850 12480 14175
rect 12544 13394 12572 14758
rect 12820 14618 12848 14894
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12912 14346 12940 15030
rect 13096 14958 13124 15302
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13084 14816 13136 14822
rect 13188 14804 13216 15642
rect 13280 15094 13308 17575
rect 13360 17546 13412 17552
rect 13372 17134 13400 17546
rect 13740 17241 13768 18022
rect 13832 17746 13860 18294
rect 14016 18290 14044 18566
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13924 17882 13952 18022
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 14016 17610 14044 18226
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 13726 17232 13782 17241
rect 13726 17167 13782 17176
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13832 16794 13860 17002
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 16794 13952 16934
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13136 14776 13216 14804
rect 13084 14758 13136 14764
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12636 13326 12664 14282
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12268 12306 12296 12582
rect 12452 12306 12480 12582
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12162 11928 12218 11937
rect 12162 11863 12164 11872
rect 12216 11863 12218 11872
rect 12164 11834 12216 11840
rect 12268 11778 12296 12242
rect 12438 12200 12494 12209
rect 12438 12135 12494 12144
rect 12176 11750 12296 11778
rect 12176 11626 12204 11750
rect 12254 11656 12310 11665
rect 12164 11620 12216 11626
rect 12254 11591 12310 11600
rect 12164 11562 12216 11568
rect 12176 8566 12204 11562
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11992 6866 12020 7822
rect 12176 7478 12204 7890
rect 12268 7546 12296 11591
rect 12452 9654 12480 12135
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12544 11286 12572 11562
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12440 9376 12492 9382
rect 12438 9344 12440 9353
rect 12492 9344 12494 9353
rect 12438 9279 12494 9288
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12544 6866 12572 11222
rect 12636 7546 12664 13262
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12238 12756 13126
rect 12912 12646 12940 13670
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12912 12374 12940 12582
rect 12900 12368 12952 12374
rect 12900 12310 12952 12316
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12728 11830 12756 12038
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12728 11558 12756 11766
rect 12820 11694 12848 12242
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12912 11558 12940 12174
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11286 12940 11494
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12728 9586 12756 10746
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12728 7954 12756 9522
rect 12820 9518 12848 10406
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12820 9178 12848 9454
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12912 8634 12940 10950
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12912 7750 12940 8570
rect 13004 8090 13032 14758
rect 13096 13462 13124 14758
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13280 13734 13308 14350
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13084 13456 13136 13462
rect 13280 13433 13308 13670
rect 13084 13398 13136 13404
rect 13266 13424 13322 13433
rect 13176 13388 13228 13394
rect 13266 13359 13322 13368
rect 13176 13330 13228 13336
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13096 12850 13124 13262
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13096 11014 13124 12786
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13096 10266 13124 10474
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13096 9586 13124 10202
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13096 9178 13124 9522
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 13188 7546 13216 13330
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13280 11830 13308 13262
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13280 7546 13308 11630
rect 13372 8090 13400 16730
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13556 15366 13584 16594
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13450 13832 13506 13841
rect 13450 13767 13506 13776
rect 13464 13530 13492 13767
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13452 12232 13504 12238
rect 13450 12200 13452 12209
rect 13504 12200 13506 12209
rect 13450 12135 13506 12144
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13464 11898 13492 12038
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13464 11354 13492 11630
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 10130 13492 10542
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13464 7410 13492 10066
rect 13556 8090 13584 15302
rect 13648 14249 13676 16594
rect 13832 15434 13860 16730
rect 13924 16658 13952 16730
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 14016 15910 14044 16526
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13924 15706 13952 15846
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13924 15570 13952 15642
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13832 14482 13860 15370
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13634 14240 13690 14249
rect 13634 14175 13690 14184
rect 13740 14090 13768 14418
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13648 14062 13768 14090
rect 13832 14074 13860 14214
rect 13820 14068 13872 14074
rect 13648 13530 13676 14062
rect 13820 14010 13872 14016
rect 13726 13968 13782 13977
rect 13726 13903 13782 13912
rect 13740 13734 13768 13903
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13740 13297 13768 13398
rect 13832 13394 13860 13806
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13726 13288 13782 13297
rect 13726 13223 13782 13232
rect 13636 13184 13688 13190
rect 13688 13132 13860 13138
rect 13636 13126 13860 13132
rect 13648 13110 13860 13126
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13648 11626 13676 12310
rect 13726 12064 13782 12073
rect 13726 11999 13782 12008
rect 13740 11626 13768 11999
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13832 11354 13860 13110
rect 13924 12918 13952 14894
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13924 12714 13952 12854
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10470 13768 11086
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10198 13768 10406
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13740 8838 13768 10134
rect 13832 9654 13860 11290
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13740 8634 13768 8774
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13924 8090 13952 11222
rect 14016 8566 14044 14962
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14108 14113 14136 14418
rect 14094 14104 14150 14113
rect 14094 14039 14150 14048
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14108 10674 14136 11766
rect 14200 11626 14228 19264
rect 14280 19246 14332 19252
rect 14280 18896 14332 18902
rect 14280 18838 14332 18844
rect 14292 17270 14320 18838
rect 14384 18222 14412 19654
rect 14476 19009 14504 19858
rect 15028 19174 15056 20590
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15120 20058 15148 20198
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15016 19168 15068 19174
rect 15120 19145 15148 19858
rect 15212 19174 15240 22000
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15304 20058 15332 20266
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15672 19174 15700 22000
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15200 19168 15252 19174
rect 15016 19110 15068 19116
rect 15106 19136 15162 19145
rect 14684 19068 14980 19088
rect 15200 19110 15252 19116
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15106 19071 15162 19080
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14462 19000 14518 19009
rect 14684 18992 14980 19012
rect 15106 19000 15162 19009
rect 14462 18935 14518 18944
rect 15106 18935 15162 18944
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15028 18358 15056 18566
rect 15120 18465 15148 18935
rect 15856 18902 15884 19246
rect 16132 19174 16160 22000
rect 16592 20058 16620 22000
rect 17052 20058 17080 22000
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15106 18456 15162 18465
rect 15106 18391 15162 18400
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15016 18352 15068 18358
rect 14462 18320 14518 18329
rect 15016 18294 15068 18300
rect 14462 18255 14518 18264
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14476 18086 14504 18255
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14476 17513 14504 17750
rect 14568 17746 14596 18158
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 15028 17678 15056 18294
rect 15396 18290 15424 18362
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 15292 18148 15344 18154
rect 15292 18090 15344 18096
rect 15108 18080 15160 18086
rect 15304 18034 15332 18090
rect 15108 18022 15160 18028
rect 15120 17746 15148 18022
rect 15212 18006 15332 18034
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14462 17504 14518 17513
rect 14462 17439 14518 17448
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14292 16590 14320 17206
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14476 16794 14504 17070
rect 15028 17066 15056 17614
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 15120 16998 15148 17682
rect 15212 17610 15240 18006
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 15978 14320 16526
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14292 15502 14320 15914
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14292 14278 14320 14894
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 12986 14320 14214
rect 14384 13977 14412 14758
rect 14568 14482 14596 16934
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15304 16794 15332 17614
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14924 15632 14976 15638
rect 14844 15592 14924 15620
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14752 14958 14780 15506
rect 14844 15026 14872 15592
rect 14924 15574 14976 15580
rect 15120 15570 15148 15846
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15212 15026 15240 16390
rect 15304 16182 15332 16730
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15396 15042 15424 18022
rect 15488 17921 15516 18770
rect 16408 18766 16436 19246
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 18290 15608 18566
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15474 17912 15530 17921
rect 15474 17847 15530 17856
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15304 15014 15424 15042
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 15212 14414 15240 14962
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 14464 14272 14516 14278
rect 14462 14240 14464 14249
rect 14516 14240 14518 14249
rect 14462 14175 14518 14184
rect 14462 14104 14518 14113
rect 14462 14039 14518 14048
rect 14370 13968 14426 13977
rect 14370 13903 14426 13912
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14384 13530 14412 13738
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14384 12850 14412 13466
rect 14476 13326 14504 14039
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14464 13320 14516 13326
rect 15212 13297 15240 14350
rect 14464 13262 14516 13268
rect 15014 13288 15070 13297
rect 15014 13223 15070 13232
rect 15198 13288 15254 13297
rect 15198 13223 15254 13232
rect 14832 13184 14884 13190
rect 14462 13152 14518 13161
rect 14832 13126 14884 13132
rect 14462 13087 14518 13096
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14292 12442 14320 12786
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14372 12300 14424 12306
rect 14292 12260 14372 12288
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14108 10130 14136 10610
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14186 9752 14242 9761
rect 14186 9687 14242 9696
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 10704 6458 10732 6598
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 11624 6254 11652 6598
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 12176 5846 12204 6190
rect 12728 5914 12756 6394
rect 13464 6390 13492 7346
rect 14200 6866 14228 9687
rect 14292 8430 14320 12260
rect 14372 12242 14424 12248
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14384 8498 14412 11562
rect 14476 8634 14504 13087
rect 14844 12850 14872 13126
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14568 12306 14596 12650
rect 15028 12646 15056 13223
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 15028 12238 15056 12582
rect 15212 12374 15240 12718
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14568 9654 14596 11154
rect 14660 11082 14688 11154
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15028 9110 15056 11154
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15120 10538 15148 11086
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15120 9994 15148 10474
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 15120 9382 15148 9930
rect 15212 9518 15240 12174
rect 15304 11150 15332 15014
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15396 14482 15424 14894
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15396 13734 15424 14282
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15396 13530 15424 13670
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15488 13410 15516 17847
rect 15580 17746 15608 18226
rect 16132 18222 16160 18702
rect 16500 18612 16528 18770
rect 16592 18766 16620 19858
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16684 18630 16712 19654
rect 17052 19514 17080 19654
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16672 18624 16724 18630
rect 16500 18584 16620 18612
rect 16592 18329 16620 18584
rect 16672 18566 16724 18572
rect 16578 18320 16634 18329
rect 16578 18255 16634 18264
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 16040 18086 16068 18158
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15580 17354 15608 17682
rect 15580 17326 15700 17354
rect 15672 17270 15700 17326
rect 15660 17264 15712 17270
rect 15660 17206 15712 17212
rect 15672 16794 15700 17206
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 16040 16658 16068 18022
rect 16132 17785 16160 18022
rect 16118 17776 16174 17785
rect 16118 17711 16174 17720
rect 16500 17678 16528 18090
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16224 17202 16252 17478
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16316 17082 16344 17478
rect 16500 17270 16528 17614
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16224 17066 16344 17082
rect 16212 17060 16344 17066
rect 16264 17054 16344 17060
rect 16212 17002 16264 17008
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16304 16584 16356 16590
rect 16356 16532 16436 16538
rect 16304 16526 16436 16532
rect 16316 16510 16436 16526
rect 16408 16182 16436 16510
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 13462 15608 15846
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15672 14618 15700 15030
rect 15764 15026 15792 15302
rect 16132 15162 16160 15982
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 15706 16252 15846
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15672 14006 15700 14554
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15948 13462 15976 14418
rect 15396 13382 15516 13410
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 15396 11286 15424 13382
rect 15580 12986 15608 13398
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15568 12300 15620 12306
rect 15672 12288 15700 13262
rect 15620 12260 15700 12288
rect 15568 12242 15620 12248
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15304 10198 15332 11086
rect 15488 11082 15516 11562
rect 15580 11558 15608 12242
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15488 10810 15516 11018
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15120 9178 15148 9318
rect 15488 9178 15516 10746
rect 15580 10606 15608 11494
rect 15672 11354 15700 11562
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15672 9722 15700 11154
rect 16132 11082 16160 15098
rect 16316 14958 16344 15438
rect 16408 15366 16436 16118
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16408 15162 16436 15302
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16316 14346 16344 14894
rect 16304 14340 16356 14346
rect 16304 14282 16356 14288
rect 16408 13870 16436 15098
rect 16592 14498 16620 18255
rect 16776 17746 16804 18770
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16868 17785 16896 18566
rect 17328 18154 17356 19926
rect 17512 19242 17540 22000
rect 17972 20058 18000 22000
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 18432 19786 18460 22000
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18708 19446 18736 19858
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 17500 19236 17552 19242
rect 17500 19178 17552 19184
rect 17604 18630 17632 19246
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17592 18624 17644 18630
rect 17696 18601 17724 19110
rect 17592 18566 17644 18572
rect 17682 18592 17738 18601
rect 17682 18527 17738 18536
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 16948 17808 17000 17814
rect 16854 17776 16910 17785
rect 16764 17740 16816 17746
rect 16948 17750 17000 17756
rect 16854 17711 16910 17720
rect 16764 17682 16816 17688
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16500 14470 16620 14498
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16500 13716 16528 14470
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16592 13870 16620 14282
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16500 13688 16620 13716
rect 16592 13258 16620 13688
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16684 13138 16712 16934
rect 16776 15638 16804 17682
rect 16764 15632 16816 15638
rect 16764 15574 16816 15580
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16776 14890 16804 15302
rect 16868 15026 16896 17711
rect 16960 17270 16988 17750
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 16948 17264 17000 17270
rect 16948 17206 17000 17212
rect 17328 17202 17356 17614
rect 17420 17610 17448 18226
rect 17788 18057 17816 19246
rect 18156 18834 18184 19246
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 17868 18828 17920 18834
rect 18144 18828 18196 18834
rect 17920 18788 18000 18816
rect 17868 18770 17920 18776
rect 17774 18048 17830 18057
rect 17774 17983 17830 17992
rect 17682 17776 17738 17785
rect 17682 17711 17684 17720
rect 17736 17711 17738 17720
rect 17684 17682 17736 17688
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17500 17536 17552 17542
rect 17604 17513 17632 17546
rect 17500 17478 17552 17484
rect 17590 17504 17646 17513
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17512 16726 17540 17478
rect 17590 17439 17646 17448
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17604 16794 17632 17138
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17684 16652 17736 16658
rect 17788 16640 17816 17206
rect 17880 17066 17908 17614
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17736 16612 17816 16640
rect 17684 16594 17736 16600
rect 17144 15910 17172 16594
rect 17590 16552 17646 16561
rect 17590 16487 17646 16496
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17144 15502 17172 15846
rect 17132 15496 17184 15502
rect 17604 15473 17632 16487
rect 17132 15438 17184 15444
rect 17590 15464 17646 15473
rect 17144 15162 17172 15438
rect 17590 15399 17646 15408
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16776 14414 16804 14826
rect 16868 14414 16896 14962
rect 17316 14884 17368 14890
rect 17316 14826 17368 14832
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16500 13110 16712 13138
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16224 11218 16252 12038
rect 16316 11830 16344 12242
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16500 11676 16528 13110
rect 16776 12442 16804 14350
rect 16960 13530 16988 14418
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16960 13410 16988 13466
rect 16868 13382 16988 13410
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16316 11648 16528 11676
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 15842 10568 15898 10577
rect 15842 10503 15898 10512
rect 16028 10532 16080 10538
rect 15856 10198 15884 10503
rect 16028 10474 16080 10480
rect 15844 10192 15896 10198
rect 15844 10134 15896 10140
rect 15856 9722 15884 10134
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15948 9382 15976 10066
rect 16040 10062 16068 10474
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15016 9104 15068 9110
rect 15016 9046 15068 9052
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14292 8090 14320 8366
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 15948 7818 15976 9318
rect 16040 9042 16068 9998
rect 16316 9450 16344 11648
rect 16684 11558 16712 12106
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16408 10606 16436 10950
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16408 10130 16436 10542
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16040 8634 16068 8978
rect 16408 8634 16436 10066
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7410 15056 7686
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 16684 7342 16712 11086
rect 16868 9110 16896 13382
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16960 12170 16988 13194
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17144 12442 17172 12582
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11354 16988 11494
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 10198 17172 10406
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17052 9450 17080 9862
rect 17144 9586 17172 10134
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17040 9444 17092 9450
rect 17040 9386 17092 9392
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 17052 9042 17080 9386
rect 17144 9178 17172 9522
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16868 8090 16896 8570
rect 17328 8362 17356 14826
rect 17512 14822 17540 15302
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17604 12782 17632 15399
rect 17696 15026 17724 16594
rect 17880 16250 17908 17002
rect 17972 16250 18000 18788
rect 18144 18770 18196 18776
rect 18340 18612 18368 19178
rect 18420 18828 18472 18834
rect 18472 18788 18644 18816
rect 18420 18770 18472 18776
rect 18340 18584 18552 18612
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18524 18222 18552 18584
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18510 18048 18566 18057
rect 18510 17983 18566 17992
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18052 16720 18104 16726
rect 18050 16688 18052 16697
rect 18104 16688 18106 16697
rect 18050 16623 18106 16632
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17880 15706 17908 15982
rect 17972 15706 18000 16186
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17788 14346 17816 15302
rect 17972 14890 18000 15506
rect 18420 15496 18472 15502
rect 18524 15473 18552 17983
rect 18420 15438 18472 15444
rect 18510 15464 18566 15473
rect 18432 15348 18460 15438
rect 18510 15399 18566 15408
rect 18432 15320 18552 15348
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17960 14408 18012 14414
rect 18340 14396 18368 14894
rect 18524 14770 18552 15320
rect 18432 14742 18552 14770
rect 18432 14550 18460 14742
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18420 14408 18472 14414
rect 18340 14376 18420 14396
rect 18472 14376 18474 14385
rect 18340 14368 18418 14376
rect 17960 14350 18012 14356
rect 17776 14340 17828 14346
rect 17776 14282 17828 14288
rect 17972 13870 18000 14350
rect 18418 14311 18474 14320
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 18524 13802 18552 14554
rect 18616 14006 18644 18788
rect 18708 15570 18736 19382
rect 18892 18426 18920 22000
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18984 18766 19012 19858
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18788 18352 18840 18358
rect 18786 18320 18788 18329
rect 18840 18320 18842 18329
rect 18786 18255 18842 18264
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18800 15586 18828 18158
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 18892 15706 18920 15914
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18696 15564 18748 15570
rect 18800 15558 18920 15586
rect 18696 15506 18748 15512
rect 18694 15464 18750 15473
rect 18694 15399 18750 15408
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17696 13462 17724 13670
rect 18524 13462 18552 13738
rect 17684 13456 17736 13462
rect 18512 13456 18564 13462
rect 17684 13398 17736 13404
rect 18050 13424 18106 13433
rect 18512 13398 18564 13404
rect 18050 13359 18106 13368
rect 18064 13258 18092 13359
rect 18616 13274 18644 13942
rect 18708 13326 18736 15399
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18800 13530 18828 14486
rect 18892 13530 18920 15558
rect 18984 14618 19012 18702
rect 19076 18306 19104 19450
rect 19352 19394 19380 22000
rect 19812 19802 19840 22000
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 20088 20058 20116 20334
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 19812 19774 20116 19802
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19352 19366 19564 19394
rect 19338 19272 19394 19281
rect 19338 19207 19340 19216
rect 19392 19207 19394 19216
rect 19340 19178 19392 19184
rect 19430 18864 19486 18873
rect 19430 18799 19486 18808
rect 19156 18760 19208 18766
rect 19154 18728 19156 18737
rect 19208 18728 19210 18737
rect 19154 18663 19210 18672
rect 19444 18426 19472 18799
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19076 18278 19196 18306
rect 19064 18216 19116 18222
rect 19062 18184 19064 18193
rect 19116 18184 19118 18193
rect 19062 18119 19118 18128
rect 19062 17776 19118 17785
rect 19062 17711 19064 17720
rect 19116 17711 19118 17720
rect 19064 17682 19116 17688
rect 19062 17232 19118 17241
rect 19062 17167 19064 17176
rect 19116 17167 19118 17176
rect 19064 17138 19116 17144
rect 19168 14929 19196 18278
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19260 17649 19288 18022
rect 19246 17640 19302 17649
rect 19246 17575 19302 17584
rect 19340 17536 19392 17542
rect 19260 17484 19340 17490
rect 19260 17478 19392 17484
rect 19260 17462 19380 17478
rect 19260 17338 19288 17462
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19340 16992 19392 16998
rect 19338 16960 19340 16969
rect 19432 16992 19484 16998
rect 19392 16960 19394 16969
rect 19432 16934 19484 16940
rect 19338 16895 19394 16904
rect 19338 16824 19394 16833
rect 19260 16782 19338 16810
rect 19260 16561 19288 16782
rect 19338 16759 19394 16768
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19246 16552 19302 16561
rect 19246 16487 19302 16496
rect 19352 16250 19380 16594
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19260 15978 19288 16050
rect 19248 15972 19300 15978
rect 19248 15914 19300 15920
rect 19260 15094 19288 15914
rect 19444 15706 19472 16934
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19444 15502 19472 15642
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19154 14920 19210 14929
rect 19154 14855 19210 14864
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 18972 13932 19024 13938
rect 19024 13892 19104 13920
rect 18972 13874 19024 13880
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 18524 13246 18644 13274
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18524 12986 18552 13246
rect 19076 13190 19104 13892
rect 19168 13734 19196 14855
rect 19260 14550 19288 15030
rect 19352 14550 19380 15098
rect 19444 14958 19472 15438
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19338 14376 19394 14385
rect 19338 14311 19394 14320
rect 19246 13968 19302 13977
rect 19246 13903 19248 13912
rect 19300 13903 19302 13912
rect 19248 13874 19300 13880
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 17592 12776 17644 12782
rect 17960 12776 18012 12782
rect 17644 12724 17724 12730
rect 17592 12718 17724 12724
rect 17960 12718 18012 12724
rect 17604 12702 17724 12718
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17604 12170 17632 12582
rect 17696 12306 17724 12702
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17604 11830 17632 12106
rect 17696 12102 17724 12242
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17684 12096 17736 12102
rect 17788 12073 17816 12174
rect 17684 12038 17736 12044
rect 17774 12064 17830 12073
rect 17774 11999 17830 12008
rect 17788 11830 17816 11999
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17972 11354 18000 12718
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18524 12442 18552 12650
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18616 12306 18644 13126
rect 19076 12986 19104 13126
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 9722 17448 10406
rect 17788 9761 17816 11154
rect 18064 11132 18092 11630
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 18156 11150 18184 11562
rect 18524 11286 18552 12174
rect 18616 11626 18644 12242
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 17972 11104 18092 11132
rect 18144 11144 18196 11150
rect 17972 11014 18000 11104
rect 18144 11086 18196 11092
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10810 18000 10950
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 18524 10266 18552 11222
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18616 10130 18644 11562
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18800 10266 18828 11018
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 17774 9752 17830 9761
rect 17408 9716 17460 9722
rect 18116 9744 18412 9764
rect 17774 9687 17830 9696
rect 17408 9658 17460 9664
rect 17420 9518 17448 9658
rect 17788 9586 17816 9687
rect 19168 9654 19196 13262
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19260 11286 19288 11562
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19352 11150 19380 14311
rect 19444 14006 19472 14758
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19444 11898 19472 12786
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19444 11354 19472 11834
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19444 10606 19472 11290
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 19352 9178 19380 9522
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 17512 8634 17540 9114
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 19536 7546 19564 19366
rect 19812 19310 19840 19654
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19628 17626 19656 19178
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19996 18222 20024 18566
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19708 18148 19760 18154
rect 19708 18090 19760 18096
rect 19892 18148 19944 18154
rect 19892 18090 19944 18096
rect 19720 18034 19748 18090
rect 19720 18006 19840 18034
rect 19628 17598 19748 17626
rect 19616 17060 19668 17066
rect 19616 17002 19668 17008
rect 19628 16794 19656 17002
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19628 15706 19656 15846
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19616 14952 19668 14958
rect 19614 14920 19616 14929
rect 19668 14920 19670 14929
rect 19614 14855 19670 14864
rect 19720 13841 19748 17598
rect 19812 16794 19840 18006
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19812 14006 19840 14214
rect 19800 14000 19852 14006
rect 19800 13942 19852 13948
rect 19706 13832 19762 13841
rect 19706 13767 19762 13776
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19812 11558 19840 12242
rect 19616 11552 19668 11558
rect 19800 11552 19852 11558
rect 19616 11494 19668 11500
rect 19798 11520 19800 11529
rect 19852 11520 19854 11529
rect 19628 11354 19656 11494
rect 19798 11455 19854 11464
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19628 10266 19656 10678
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19628 9722 19656 10202
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 6458 13584 6598
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 19076 6118 19104 6802
rect 19904 6730 19932 18090
rect 19984 18080 20036 18086
rect 19982 18048 19984 18057
rect 20036 18048 20038 18057
rect 19982 17983 20038 17992
rect 19984 16992 20036 16998
rect 19982 16960 19984 16969
rect 20036 16960 20038 16969
rect 19982 16895 20038 16904
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19996 9586 20024 10202
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19628 6458 19656 6666
rect 20088 6662 20116 19774
rect 20272 18154 20300 22000
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20456 18698 20484 19654
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20260 18148 20312 18154
rect 20260 18090 20312 18096
rect 20444 17808 20496 17814
rect 20444 17750 20496 17756
rect 20456 17338 20484 17750
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20180 15434 20208 15846
rect 20168 15428 20220 15434
rect 20168 15370 20220 15376
rect 20180 15162 20208 15370
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11558 20484 12038
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20456 11354 20484 11494
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20456 10742 20484 11290
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20548 10810 20576 11018
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 20548 10266 20576 10746
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20732 6458 20760 22000
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20824 16794 20852 19110
rect 20916 19009 20944 19110
rect 20902 19000 20958 19009
rect 20902 18935 20958 18944
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5370 9352 5510
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7760 4826 7788 5306
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8588 4826 8616 5306
rect 20272 5098 20300 5714
rect 20916 5370 20944 18158
rect 21192 5914 21220 22000
rect 21362 19136 21418 19145
rect 21362 19071 21418 19080
rect 21376 12442 21404 19071
rect 21652 18222 21680 22000
rect 22112 19310 22140 22000
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 22572 16833 22600 22000
rect 22558 16824 22614 16833
rect 22558 16759 22614 16768
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 6748 4146 6776 4762
rect 8588 4282 8616 4762
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 11164 1986 11192 4014
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 11164 1958 11468 1986
rect 5078 1592 5134 1601
rect 5078 1527 5134 1536
rect 11440 800 11468 1958
rect 3882 232 3938 241
rect 3882 167 3938 176
rect 11426 0 11482 800
<< via2 >>
rect 2042 22480 2098 22536
rect 938 19080 994 19136
rect 1306 18808 1362 18864
rect 1674 21120 1730 21176
rect 1582 20576 1638 20632
rect 1858 19216 1914 19272
rect 1766 18536 1822 18592
rect 1398 18400 1454 18456
rect 1582 16496 1638 16552
rect 1766 16904 1822 16960
rect 1766 13640 1822 13696
rect 1306 9288 1362 9344
rect 1214 9152 1270 9208
rect 1030 992 1086 1048
rect 1950 17856 2006 17912
rect 1950 17312 2006 17368
rect 1950 15408 2006 15464
rect 3238 22072 3294 22128
rect 2318 18808 2374 18864
rect 2318 17992 2374 18048
rect 2778 21528 2834 21584
rect 2686 18944 2742 19000
rect 2962 20168 3018 20224
rect 2778 18264 2834 18320
rect 2410 17720 2466 17776
rect 2870 17856 2926 17912
rect 2778 17620 2780 17640
rect 2780 17620 2832 17640
rect 2832 17620 2834 17640
rect 2778 17584 2834 17620
rect 2778 17448 2834 17504
rect 1766 9560 1822 9616
rect 2042 9696 2098 9752
rect 2226 11464 2282 11520
rect 3054 17584 3110 17640
rect 3514 19760 3570 19816
rect 3146 17040 3202 17096
rect 2686 16088 2742 16144
rect 3054 16088 3110 16144
rect 2778 15952 2834 16008
rect 2686 15000 2742 15056
rect 2594 14884 2650 14920
rect 2594 14864 2596 14884
rect 2596 14864 2648 14884
rect 2648 14864 2650 14884
rect 2502 9288 2558 9344
rect 2962 15544 3018 15600
rect 2778 13912 2834 13968
rect 2686 10240 2742 10296
rect 2686 8200 2742 8256
rect 3146 14592 3202 14648
rect 2962 7792 3018 7848
rect 2870 7248 2926 7304
rect 3606 15408 3662 15464
rect 4066 19252 4068 19272
rect 4068 19252 4120 19272
rect 4120 19252 4122 19272
rect 4066 19216 4122 19252
rect 4066 18692 4122 18728
rect 4066 18672 4068 18692
rect 4068 18672 4120 18692
rect 4120 18672 4122 18692
rect 4066 18536 4122 18592
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4434 19352 4490 19408
rect 4434 19080 4490 19136
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 5078 19080 5134 19136
rect 5354 19080 5410 19136
rect 5262 18944 5318 19000
rect 5262 18128 5318 18184
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4802 16088 4858 16144
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4894 14900 4896 14920
rect 4896 14900 4948 14920
rect 4948 14900 4950 14920
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4894 14864 4950 14900
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4066 12316 4068 12336
rect 4068 12316 4120 12336
rect 4120 12316 4122 12336
rect 4066 12280 4122 12316
rect 4066 11736 4122 11792
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4434 11500 4436 11520
rect 4436 11500 4488 11520
rect 4488 11500 4490 11520
rect 4434 11464 4490 11500
rect 4066 11328 4122 11384
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4066 10804 4122 10840
rect 4066 10784 4068 10804
rect 4068 10784 4120 10804
rect 4120 10784 4122 10804
rect 4066 10376 4122 10432
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4158 8472 4214 8528
rect 2870 3440 2926 3496
rect 1214 2896 1270 2952
rect 1122 584 1178 640
rect 4066 7520 4122 7576
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4342 7248 4398 7304
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4066 5788 4068 5808
rect 4068 5788 4120 5808
rect 4120 5788 4122 5808
rect 4066 5752 4122 5788
rect 3974 5208 4030 5264
rect 4066 4800 4122 4856
rect 3974 3848 4030 3904
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 5446 18400 5502 18456
rect 5814 18536 5870 18592
rect 6090 17856 6146 17912
rect 5078 9152 5134 9208
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4250 2488 4306 2544
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 4802 1944 4858 2000
rect 5538 13232 5594 13288
rect 6642 16652 6698 16688
rect 6642 16632 6644 16652
rect 6644 16632 6696 16652
rect 6696 16632 6698 16652
rect 5814 8356 5870 8392
rect 5814 8336 5816 8356
rect 5816 8336 5868 8356
rect 5868 8336 5870 8356
rect 5814 8064 5870 8120
rect 6090 6296 6146 6352
rect 6274 8880 6330 8936
rect 7102 17992 7158 18048
rect 7286 17604 7342 17640
rect 7286 17584 7288 17604
rect 7288 17584 7340 17604
rect 7340 17584 7342 17604
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 8666 18536 8722 18592
rect 8758 16652 8814 16688
rect 8758 16632 8760 16652
rect 8760 16632 8812 16652
rect 8812 16632 8814 16652
rect 8574 15428 8630 15464
rect 8574 15408 8576 15428
rect 8576 15408 8628 15428
rect 8628 15408 8630 15428
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 8850 14884 8906 14920
rect 8850 14864 8852 14884
rect 8852 14864 8904 14884
rect 8904 14864 8906 14884
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7286 10784 7342 10840
rect 7194 10648 7250 10704
rect 7470 9460 7472 9480
rect 7472 9460 7524 9480
rect 7524 9460 7526 9480
rect 7470 9424 7526 9460
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 8758 12688 8814 12744
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7838 7384 7894 7440
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7930 6332 7932 6352
rect 7932 6332 7984 6352
rect 7984 6332 7986 6352
rect 7930 6296 7986 6332
rect 7838 6160 7894 6216
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 8298 6704 8354 6760
rect 8758 10804 8814 10840
rect 8758 10784 8760 10804
rect 8760 10784 8812 10804
rect 8812 10784 8814 10804
rect 8850 10648 8906 10704
rect 8942 9016 8998 9072
rect 9402 14884 9458 14920
rect 9402 14864 9404 14884
rect 9404 14864 9456 14884
rect 9456 14864 9458 14884
rect 9586 17040 9642 17096
rect 9954 16668 9956 16688
rect 9956 16668 10008 16688
rect 10008 16668 10010 16688
rect 9954 16632 10010 16668
rect 9310 9968 9366 10024
rect 9218 8900 9274 8936
rect 9218 8880 9220 8900
rect 9220 8880 9272 8900
rect 9272 8880 9274 8900
rect 10322 19352 10378 19408
rect 10322 19080 10378 19136
rect 9586 7248 9642 7304
rect 10782 18400 10838 18456
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11610 18944 11666 19000
rect 11702 18808 11758 18864
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11150 17720 11206 17776
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11702 18536 11758 18592
rect 11886 18944 11942 19000
rect 11886 18808 11942 18864
rect 11886 18264 11942 18320
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11794 16904 11850 16960
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 10874 14320 10930 14376
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11518 10532 11574 10568
rect 11518 10512 11520 10532
rect 11520 10512 11572 10532
rect 11572 10512 11574 10532
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11886 14356 11888 14376
rect 11888 14356 11940 14376
rect 11940 14356 11942 14376
rect 11886 14320 11942 14356
rect 12162 18264 12218 18320
rect 12530 19080 12586 19136
rect 12438 17992 12494 18048
rect 12346 17720 12402 17776
rect 12346 16904 12402 16960
rect 11794 12980 11850 13016
rect 11794 12960 11796 12980
rect 11796 12960 11848 12980
rect 11848 12960 11850 12980
rect 11886 12008 11942 12064
rect 11702 9968 11758 10024
rect 12990 18400 13046 18456
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 13726 19080 13782 19136
rect 14094 19080 14150 19136
rect 13266 17584 13322 17640
rect 12990 15444 12992 15464
rect 12992 15444 13044 15464
rect 13044 15444 13046 15464
rect 12990 15408 13046 15444
rect 12438 14356 12440 14376
rect 12440 14356 12492 14376
rect 12492 14356 12494 14376
rect 12438 14320 12494 14356
rect 12438 14184 12494 14240
rect 13726 17176 13782 17232
rect 12162 11892 12218 11928
rect 12162 11872 12164 11892
rect 12164 11872 12216 11892
rect 12216 11872 12218 11892
rect 12438 12144 12494 12200
rect 12254 11600 12310 11656
rect 12438 9324 12440 9344
rect 12440 9324 12492 9344
rect 12492 9324 12494 9344
rect 12438 9288 12494 9324
rect 13266 13368 13322 13424
rect 13450 13776 13506 13832
rect 13450 12180 13452 12200
rect 13452 12180 13504 12200
rect 13504 12180 13506 12200
rect 13450 12144 13506 12180
rect 13634 14184 13690 14240
rect 13726 13912 13782 13968
rect 13726 13232 13782 13288
rect 13726 12008 13782 12064
rect 14094 14048 14150 14104
rect 15106 19080 15162 19136
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14462 18944 14518 19000
rect 15106 18944 15162 19000
rect 15106 18400 15162 18456
rect 14462 18264 14518 18320
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14462 17448 14518 17504
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 15474 17856 15530 17912
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14462 14220 14464 14240
rect 14464 14220 14516 14240
rect 14516 14220 14518 14240
rect 14462 14184 14518 14220
rect 14462 14048 14518 14104
rect 14370 13912 14426 13968
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 15014 13232 15070 13288
rect 15198 13232 15254 13288
rect 14462 13096 14518 13152
rect 14186 9696 14242 9752
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 16578 18264 16634 18320
rect 16118 17720 16174 17776
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 17682 18536 17738 18592
rect 16854 17720 16910 17776
rect 17774 17992 17830 18048
rect 17682 17740 17738 17776
rect 17682 17720 17684 17740
rect 17684 17720 17736 17740
rect 17736 17720 17738 17740
rect 17590 17448 17646 17504
rect 17590 16496 17646 16552
rect 17590 15408 17646 15464
rect 15842 10512 15898 10568
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18510 17992 18566 18048
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18050 16668 18052 16688
rect 18052 16668 18104 16688
rect 18104 16668 18106 16688
rect 18050 16632 18106 16668
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18510 15408 18566 15464
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18418 14356 18420 14376
rect 18420 14356 18472 14376
rect 18472 14356 18474 14376
rect 18418 14320 18474 14356
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18786 18300 18788 18320
rect 18788 18300 18840 18320
rect 18840 18300 18842 18320
rect 18786 18264 18842 18300
rect 18694 15408 18750 15464
rect 18050 13368 18106 13424
rect 19338 19236 19394 19272
rect 19338 19216 19340 19236
rect 19340 19216 19392 19236
rect 19392 19216 19394 19236
rect 19430 18808 19486 18864
rect 19154 18708 19156 18728
rect 19156 18708 19208 18728
rect 19208 18708 19210 18728
rect 19154 18672 19210 18708
rect 19062 18164 19064 18184
rect 19064 18164 19116 18184
rect 19116 18164 19118 18184
rect 19062 18128 19118 18164
rect 19062 17740 19118 17776
rect 19062 17720 19064 17740
rect 19064 17720 19116 17740
rect 19116 17720 19118 17740
rect 19062 17196 19118 17232
rect 19062 17176 19064 17196
rect 19064 17176 19116 17196
rect 19116 17176 19118 17196
rect 19246 17584 19302 17640
rect 19338 16940 19340 16960
rect 19340 16940 19392 16960
rect 19392 16940 19394 16960
rect 19338 16904 19394 16940
rect 19338 16768 19394 16824
rect 19246 16496 19302 16552
rect 19154 14864 19210 14920
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 19338 14320 19394 14376
rect 19246 13932 19302 13968
rect 19246 13912 19248 13932
rect 19248 13912 19300 13932
rect 19300 13912 19302 13932
rect 17774 12008 17830 12064
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17774 9696 17830 9752
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 19614 14900 19616 14920
rect 19616 14900 19668 14920
rect 19668 14900 19670 14920
rect 19614 14864 19670 14900
rect 19706 13776 19762 13832
rect 19798 11500 19800 11520
rect 19800 11500 19852 11520
rect 19852 11500 19854 11520
rect 19798 11464 19854 11500
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 19982 18028 19984 18048
rect 19984 18028 20036 18048
rect 20036 18028 20038 18048
rect 19982 17992 20038 18028
rect 19982 16940 19984 16960
rect 19984 16940 20036 16960
rect 20036 16940 20038 16960
rect 19982 16904 20038 16940
rect 20902 18944 20958 19000
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 21362 19080 21418 19136
rect 22558 16768 22614 16824
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 5078 1536 5134 1592
rect 3882 176 3938 232
<< metal3 >>
rect 0 22538 800 22568
rect 2037 22538 2103 22541
rect 0 22536 2103 22538
rect 0 22480 2042 22536
rect 2098 22480 2103 22536
rect 0 22478 2103 22480
rect 0 22448 800 22478
rect 2037 22475 2103 22478
rect 0 22130 800 22160
rect 3233 22130 3299 22133
rect 0 22128 3299 22130
rect 0 22072 3238 22128
rect 3294 22072 3299 22128
rect 0 22070 3299 22072
rect 0 22040 800 22070
rect 3233 22067 3299 22070
rect 0 21586 800 21616
rect 2773 21586 2839 21589
rect 0 21584 2839 21586
rect 0 21528 2778 21584
rect 2834 21528 2839 21584
rect 0 21526 2839 21528
rect 0 21496 800 21526
rect 2773 21523 2839 21526
rect 0 21178 800 21208
rect 1669 21178 1735 21181
rect 0 21176 1735 21178
rect 0 21120 1674 21176
rect 1730 21120 1735 21176
rect 0 21118 1735 21120
rect 0 21088 800 21118
rect 1669 21115 1735 21118
rect 0 20634 800 20664
rect 1577 20634 1643 20637
rect 0 20632 1643 20634
rect 0 20576 1582 20632
rect 1638 20576 1643 20632
rect 0 20574 1643 20576
rect 0 20544 800 20574
rect 1577 20571 1643 20574
rect 0 20226 800 20256
rect 2957 20226 3023 20229
rect 0 20224 3023 20226
rect 0 20168 2962 20224
rect 3018 20168 3023 20224
rect 0 20166 3023 20168
rect 0 20136 800 20166
rect 2957 20163 3023 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19818 800 19848
rect 3509 19818 3575 19821
rect 0 19816 3575 19818
rect 0 19760 3514 19816
rect 3570 19760 3575 19816
rect 0 19758 3575 19760
rect 0 19728 800 19758
rect 3509 19755 3575 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 4429 19410 4495 19413
rect 10317 19410 10383 19413
rect 4429 19408 10383 19410
rect 4429 19352 4434 19408
rect 4490 19352 10322 19408
rect 10378 19352 10383 19408
rect 4429 19350 10383 19352
rect 4429 19347 4495 19350
rect 10317 19347 10383 19350
rect 0 19274 800 19304
rect 1853 19274 1919 19277
rect 0 19272 1919 19274
rect 0 19216 1858 19272
rect 1914 19216 1919 19272
rect 0 19214 1919 19216
rect 0 19184 800 19214
rect 1853 19211 1919 19214
rect 4061 19274 4127 19277
rect 19333 19274 19399 19277
rect 4061 19272 19399 19274
rect 4061 19216 4066 19272
rect 4122 19216 19338 19272
rect 19394 19216 19399 19272
rect 4061 19214 19399 19216
rect 4061 19211 4127 19214
rect 19333 19211 19399 19214
rect 933 19138 999 19141
rect 4429 19138 4495 19141
rect 933 19136 4495 19138
rect 933 19080 938 19136
rect 994 19080 4434 19136
rect 4490 19080 4495 19136
rect 933 19078 4495 19080
rect 933 19075 999 19078
rect 4429 19075 4495 19078
rect 5073 19138 5139 19141
rect 5349 19138 5415 19141
rect 5073 19136 5415 19138
rect 5073 19080 5078 19136
rect 5134 19080 5354 19136
rect 5410 19080 5415 19136
rect 5073 19078 5415 19080
rect 5073 19075 5139 19078
rect 5349 19075 5415 19078
rect 10317 19138 10383 19141
rect 12525 19138 12591 19141
rect 13721 19138 13787 19141
rect 10317 19136 13787 19138
rect 10317 19080 10322 19136
rect 10378 19080 12530 19136
rect 12586 19080 13726 19136
rect 13782 19080 13787 19136
rect 10317 19078 13787 19080
rect 10317 19075 10383 19078
rect 12525 19075 12591 19078
rect 13721 19075 13787 19078
rect 14089 19138 14155 19141
rect 14222 19138 14228 19140
rect 14089 19136 14228 19138
rect 14089 19080 14094 19136
rect 14150 19080 14228 19136
rect 14089 19078 14228 19080
rect 14089 19075 14155 19078
rect 14222 19076 14228 19078
rect 14292 19076 14298 19140
rect 15101 19138 15167 19141
rect 21357 19138 21423 19141
rect 15101 19136 21423 19138
rect 15101 19080 15106 19136
rect 15162 19080 21362 19136
rect 21418 19080 21423 19136
rect 15101 19078 21423 19080
rect 15101 19075 15167 19078
rect 21357 19075 21423 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 2681 19002 2747 19005
rect 5257 19002 5323 19005
rect 11605 19004 11671 19005
rect 11605 19002 11652 19004
rect 2681 19000 5323 19002
rect 2681 18944 2686 19000
rect 2742 18944 5262 19000
rect 5318 18944 5323 19000
rect 2681 18942 5323 18944
rect 11560 19000 11652 19002
rect 11560 18944 11610 19000
rect 11560 18942 11652 18944
rect 2681 18939 2747 18942
rect 5257 18939 5323 18942
rect 11605 18940 11652 18942
rect 11716 18940 11722 19004
rect 11881 19002 11947 19005
rect 14457 19002 14523 19005
rect 11881 19000 14523 19002
rect 11881 18944 11886 19000
rect 11942 18944 14462 19000
rect 14518 18944 14523 19000
rect 11881 18942 14523 18944
rect 11605 18939 11671 18940
rect 11881 18939 11947 18942
rect 14457 18939 14523 18942
rect 15101 19002 15167 19005
rect 20897 19002 20963 19005
rect 15101 19000 20963 19002
rect 15101 18944 15106 19000
rect 15162 18944 20902 19000
rect 20958 18944 20963 19000
rect 15101 18942 20963 18944
rect 15101 18939 15167 18942
rect 20897 18939 20963 18942
rect 0 18866 800 18896
rect 1301 18866 1367 18869
rect 0 18864 1367 18866
rect 0 18808 1306 18864
rect 1362 18808 1367 18864
rect 0 18806 1367 18808
rect 0 18776 800 18806
rect 1301 18803 1367 18806
rect 2313 18866 2379 18869
rect 11697 18866 11763 18869
rect 2313 18864 11763 18866
rect 2313 18808 2318 18864
rect 2374 18808 11702 18864
rect 11758 18808 11763 18864
rect 2313 18806 11763 18808
rect 2313 18803 2379 18806
rect 11697 18803 11763 18806
rect 11881 18866 11947 18869
rect 19425 18866 19491 18869
rect 11881 18864 19491 18866
rect 11881 18808 11886 18864
rect 11942 18808 19430 18864
rect 19486 18808 19491 18864
rect 11881 18806 19491 18808
rect 11881 18803 11947 18806
rect 19425 18803 19491 18806
rect 4061 18730 4127 18733
rect 19149 18730 19215 18733
rect 4061 18728 19215 18730
rect 4061 18672 4066 18728
rect 4122 18672 19154 18728
rect 19210 18672 19215 18728
rect 4061 18670 19215 18672
rect 4061 18667 4127 18670
rect 19149 18667 19215 18670
rect 1761 18594 1827 18597
rect 4061 18594 4127 18597
rect 1761 18592 4127 18594
rect 1761 18536 1766 18592
rect 1822 18536 4066 18592
rect 4122 18536 4127 18592
rect 1761 18534 4127 18536
rect 1761 18531 1827 18534
rect 4061 18531 4127 18534
rect 5809 18594 5875 18597
rect 8661 18594 8727 18597
rect 5809 18592 8727 18594
rect 5809 18536 5814 18592
rect 5870 18536 8666 18592
rect 8722 18536 8727 18592
rect 5809 18534 8727 18536
rect 5809 18531 5875 18534
rect 8661 18531 8727 18534
rect 11697 18594 11763 18597
rect 17677 18594 17743 18597
rect 11697 18592 17743 18594
rect 11697 18536 11702 18592
rect 11758 18536 17682 18592
rect 17738 18536 17743 18592
rect 11697 18534 17743 18536
rect 11697 18531 11763 18534
rect 17677 18531 17743 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 1393 18458 1459 18461
rect 5441 18458 5507 18461
rect 10777 18458 10843 18461
rect 1393 18456 4170 18458
rect 1393 18400 1398 18456
rect 1454 18400 4170 18456
rect 1393 18398 4170 18400
rect 1393 18395 1459 18398
rect 0 18322 800 18352
rect 2773 18322 2839 18325
rect 0 18320 2839 18322
rect 0 18264 2778 18320
rect 2834 18264 2839 18320
rect 0 18262 2839 18264
rect 4110 18322 4170 18398
rect 5441 18456 10843 18458
rect 5441 18400 5446 18456
rect 5502 18400 10782 18456
rect 10838 18400 10843 18456
rect 5441 18398 10843 18400
rect 5441 18395 5507 18398
rect 10777 18395 10843 18398
rect 12566 18396 12572 18460
rect 12636 18458 12642 18460
rect 12985 18458 13051 18461
rect 15101 18458 15167 18461
rect 12636 18456 15167 18458
rect 12636 18400 12990 18456
rect 13046 18400 15106 18456
rect 15162 18400 15167 18456
rect 12636 18398 15167 18400
rect 12636 18396 12642 18398
rect 12985 18395 13051 18398
rect 15101 18395 15167 18398
rect 11881 18322 11947 18325
rect 4110 18320 11947 18322
rect 4110 18264 11886 18320
rect 11942 18264 11947 18320
rect 4110 18262 11947 18264
rect 0 18232 800 18262
rect 2773 18259 2839 18262
rect 11881 18259 11947 18262
rect 12157 18322 12223 18325
rect 14457 18322 14523 18325
rect 12157 18320 14523 18322
rect 12157 18264 12162 18320
rect 12218 18264 14462 18320
rect 14518 18264 14523 18320
rect 12157 18262 14523 18264
rect 12157 18259 12223 18262
rect 14457 18259 14523 18262
rect 16573 18322 16639 18325
rect 18781 18322 18847 18325
rect 16573 18320 18847 18322
rect 16573 18264 16578 18320
rect 16634 18264 18786 18320
rect 18842 18264 18847 18320
rect 16573 18262 18847 18264
rect 16573 18259 16639 18262
rect 18781 18259 18847 18262
rect 5257 18186 5323 18189
rect 19057 18186 19123 18189
rect 5257 18184 19123 18186
rect 5257 18128 5262 18184
rect 5318 18128 19062 18184
rect 19118 18128 19123 18184
rect 5257 18126 19123 18128
rect 5257 18123 5323 18126
rect 19057 18123 19123 18126
rect 2313 18050 2379 18053
rect 7097 18050 7163 18053
rect 12433 18052 12499 18053
rect 2313 18048 7163 18050
rect 2313 17992 2318 18048
rect 2374 17992 7102 18048
rect 7158 17992 7163 18048
rect 2313 17990 7163 17992
rect 2313 17987 2379 17990
rect 7097 17987 7163 17990
rect 12382 17988 12388 18052
rect 12452 18050 12499 18052
rect 17769 18050 17835 18053
rect 18505 18050 18571 18053
rect 19977 18050 20043 18053
rect 12452 18048 12544 18050
rect 12494 17992 12544 18048
rect 12452 17990 12544 17992
rect 17769 18048 18571 18050
rect 17769 17992 17774 18048
rect 17830 17992 18510 18048
rect 18566 17992 18571 18048
rect 17769 17990 18571 17992
rect 12452 17988 12499 17990
rect 12433 17987 12499 17988
rect 17769 17987 17835 17990
rect 18505 17987 18571 17990
rect 19244 18048 20043 18050
rect 19244 17992 19982 18048
rect 20038 17992 20043 18048
rect 19244 17990 20043 17992
rect 7808 17984 8128 17985
rect 0 17914 800 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1945 17914 2011 17917
rect 0 17912 2011 17914
rect 0 17856 1950 17912
rect 2006 17856 2011 17912
rect 0 17854 2011 17856
rect 0 17824 800 17854
rect 1945 17851 2011 17854
rect 2865 17914 2931 17917
rect 6085 17914 6151 17917
rect 2865 17912 6151 17914
rect 2865 17856 2870 17912
rect 2926 17856 6090 17912
rect 6146 17856 6151 17912
rect 2865 17854 6151 17856
rect 2865 17851 2931 17854
rect 6085 17851 6151 17854
rect 15469 17914 15535 17917
rect 19244 17914 19304 17990
rect 19977 17987 20043 17990
rect 15469 17912 19304 17914
rect 15469 17856 15474 17912
rect 15530 17856 19304 17912
rect 15469 17854 19304 17856
rect 15469 17851 15535 17854
rect 19198 17820 19304 17854
rect 2405 17778 2471 17781
rect 11145 17778 11211 17781
rect 2405 17776 11211 17778
rect 2405 17720 2410 17776
rect 2466 17720 11150 17776
rect 11206 17720 11211 17776
rect 2405 17718 11211 17720
rect 2405 17715 2471 17718
rect 11145 17715 11211 17718
rect 12341 17778 12407 17781
rect 16113 17778 16179 17781
rect 16849 17778 16915 17781
rect 12341 17776 16915 17778
rect 12341 17720 12346 17776
rect 12402 17720 16118 17776
rect 16174 17720 16854 17776
rect 16910 17720 16915 17776
rect 12341 17718 16915 17720
rect 12341 17715 12407 17718
rect 16113 17715 16179 17718
rect 16849 17715 16915 17718
rect 17677 17778 17743 17781
rect 19057 17778 19123 17781
rect 17677 17776 19123 17778
rect 17677 17720 17682 17776
rect 17738 17720 19062 17776
rect 19118 17720 19123 17776
rect 17677 17718 19123 17720
rect 17677 17715 17743 17718
rect 19057 17715 19123 17718
rect 2773 17642 2839 17645
rect 3049 17642 3115 17645
rect 7281 17642 7347 17645
rect 2773 17640 3115 17642
rect 2773 17584 2778 17640
rect 2834 17584 3054 17640
rect 3110 17584 3115 17640
rect 2773 17582 3115 17584
rect 2773 17579 2839 17582
rect 3049 17579 3115 17582
rect 4110 17640 7347 17642
rect 4110 17584 7286 17640
rect 7342 17584 7347 17640
rect 4110 17582 7347 17584
rect 2773 17506 2839 17509
rect 4110 17506 4170 17582
rect 7281 17579 7347 17582
rect 13261 17642 13327 17645
rect 19241 17642 19307 17645
rect 13261 17640 19307 17642
rect 13261 17584 13266 17640
rect 13322 17584 19246 17640
rect 19302 17584 19307 17640
rect 13261 17582 19307 17584
rect 13261 17579 13327 17582
rect 19241 17579 19307 17582
rect 2773 17504 4170 17506
rect 2773 17448 2778 17504
rect 2834 17448 4170 17504
rect 2773 17446 4170 17448
rect 14457 17506 14523 17509
rect 17585 17506 17651 17509
rect 14457 17504 17651 17506
rect 14457 17448 14462 17504
rect 14518 17448 17590 17504
rect 17646 17448 17651 17504
rect 14457 17446 17651 17448
rect 2773 17443 2839 17446
rect 14457 17443 14523 17446
rect 17585 17443 17651 17446
rect 4376 17440 4696 17441
rect 0 17370 800 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1945 17370 2011 17373
rect 0 17368 2011 17370
rect 0 17312 1950 17368
rect 2006 17312 2011 17368
rect 0 17310 2011 17312
rect 0 17280 800 17310
rect 1945 17307 2011 17310
rect 13721 17234 13787 17237
rect 19057 17234 19123 17237
rect 13721 17232 19123 17234
rect 13721 17176 13726 17232
rect 13782 17176 19062 17232
rect 19118 17176 19123 17232
rect 13721 17174 19123 17176
rect 13721 17171 13787 17174
rect 19057 17171 19123 17174
rect 3141 17098 3207 17101
rect 9581 17098 9647 17101
rect 3141 17096 9647 17098
rect 3141 17040 3146 17096
rect 3202 17040 9586 17096
rect 9642 17040 9647 17096
rect 3141 17038 9647 17040
rect 3141 17035 3207 17038
rect 9581 17035 9647 17038
rect 0 16962 800 16992
rect 1761 16962 1827 16965
rect 0 16960 1827 16962
rect 0 16904 1766 16960
rect 1822 16904 1827 16960
rect 0 16902 1827 16904
rect 0 16872 800 16902
rect 1761 16899 1827 16902
rect 11789 16962 11855 16965
rect 12341 16962 12407 16965
rect 11789 16960 12407 16962
rect 11789 16904 11794 16960
rect 11850 16904 12346 16960
rect 12402 16904 12407 16960
rect 11789 16902 12407 16904
rect 11789 16899 11855 16902
rect 12341 16899 12407 16902
rect 19333 16962 19399 16965
rect 19977 16962 20043 16965
rect 19333 16960 20043 16962
rect 19333 16904 19338 16960
rect 19394 16904 19982 16960
rect 20038 16904 20043 16960
rect 19333 16902 20043 16904
rect 19333 16899 19399 16902
rect 19977 16899 20043 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 19333 16826 19399 16829
rect 22553 16826 22619 16829
rect 19333 16824 22619 16826
rect 19333 16768 19338 16824
rect 19394 16768 22558 16824
rect 22614 16768 22619 16824
rect 19333 16766 22619 16768
rect 19333 16763 19399 16766
rect 22553 16763 22619 16766
rect 6637 16690 6703 16693
rect 8753 16690 8819 16693
rect 6637 16688 8819 16690
rect 6637 16632 6642 16688
rect 6698 16632 8758 16688
rect 8814 16632 8819 16688
rect 6637 16630 8819 16632
rect 6637 16627 6703 16630
rect 8753 16627 8819 16630
rect 9949 16690 10015 16693
rect 18045 16690 18111 16693
rect 9949 16688 18111 16690
rect 9949 16632 9954 16688
rect 10010 16632 18050 16688
rect 18106 16632 18111 16688
rect 9949 16630 18111 16632
rect 9949 16627 10015 16630
rect 18045 16627 18111 16630
rect 0 16554 800 16584
rect 1577 16554 1643 16557
rect 0 16552 1643 16554
rect 0 16496 1582 16552
rect 1638 16496 1643 16552
rect 0 16494 1643 16496
rect 0 16464 800 16494
rect 1577 16491 1643 16494
rect 17585 16554 17651 16557
rect 19241 16554 19307 16557
rect 17585 16552 19307 16554
rect 17585 16496 17590 16552
rect 17646 16496 19246 16552
rect 19302 16496 19307 16552
rect 17585 16494 19307 16496
rect 17585 16491 17651 16494
rect 19241 16491 19307 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 2681 16146 2747 16149
rect 3049 16146 3115 16149
rect 4797 16146 4863 16149
rect 2681 16144 4863 16146
rect 2681 16088 2686 16144
rect 2742 16088 3054 16144
rect 3110 16088 4802 16144
rect 4858 16088 4863 16144
rect 2681 16086 4863 16088
rect 2681 16083 2747 16086
rect 3049 16083 3115 16086
rect 4797 16083 4863 16086
rect 0 16010 800 16040
rect 2773 16010 2839 16013
rect 0 16008 2839 16010
rect 0 15952 2778 16008
rect 2834 15952 2839 16008
rect 0 15950 2839 15952
rect 0 15920 800 15950
rect 2773 15947 2839 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 800 15632
rect 2957 15602 3023 15605
rect 0 15600 3023 15602
rect 0 15544 2962 15600
rect 3018 15544 3023 15600
rect 0 15542 3023 15544
rect 0 15512 800 15542
rect 2957 15539 3023 15542
rect 1945 15466 2011 15469
rect 3601 15466 3667 15469
rect 8569 15466 8635 15469
rect 1945 15464 8635 15466
rect 1945 15408 1950 15464
rect 2006 15408 3606 15464
rect 3662 15408 8574 15464
rect 8630 15408 8635 15464
rect 1945 15406 8635 15408
rect 1945 15403 2011 15406
rect 3601 15403 3667 15406
rect 8569 15403 8635 15406
rect 12985 15466 13051 15469
rect 17585 15466 17651 15469
rect 12985 15464 17651 15466
rect 12985 15408 12990 15464
rect 13046 15408 17590 15464
rect 17646 15408 17651 15464
rect 12985 15406 17651 15408
rect 12985 15403 13051 15406
rect 17585 15403 17651 15406
rect 18505 15466 18571 15469
rect 18689 15466 18755 15469
rect 18505 15464 18755 15466
rect 18505 15408 18510 15464
rect 18566 15408 18694 15464
rect 18750 15408 18755 15464
rect 18505 15406 18755 15408
rect 18505 15403 18571 15406
rect 18689 15403 18755 15406
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 800 15088
rect 2681 15058 2747 15061
rect 0 15056 2747 15058
rect 0 15000 2686 15056
rect 2742 15000 2747 15056
rect 0 14998 2747 15000
rect 0 14968 800 14998
rect 2681 14995 2747 14998
rect 2589 14922 2655 14925
rect 4889 14922 4955 14925
rect 2589 14920 4955 14922
rect 2589 14864 2594 14920
rect 2650 14864 4894 14920
rect 4950 14864 4955 14920
rect 2589 14862 4955 14864
rect 2589 14859 2655 14862
rect 4889 14859 4955 14862
rect 8845 14922 8911 14925
rect 9397 14922 9463 14925
rect 8845 14920 9463 14922
rect 8845 14864 8850 14920
rect 8906 14864 9402 14920
rect 9458 14864 9463 14920
rect 8845 14862 9463 14864
rect 8845 14859 8911 14862
rect 9397 14859 9463 14862
rect 19149 14922 19215 14925
rect 19609 14922 19675 14925
rect 19149 14920 19675 14922
rect 19149 14864 19154 14920
rect 19210 14864 19614 14920
rect 19670 14864 19675 14920
rect 19149 14862 19675 14864
rect 19149 14859 19215 14862
rect 19609 14859 19675 14862
rect 7808 14720 8128 14721
rect 0 14650 800 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 3141 14650 3207 14653
rect 0 14648 3207 14650
rect 0 14592 3146 14648
rect 3202 14592 3207 14648
rect 0 14590 3207 14592
rect 0 14560 800 14590
rect 3141 14587 3207 14590
rect 10869 14378 10935 14381
rect 11881 14378 11947 14381
rect 12433 14378 12499 14381
rect 10869 14376 12499 14378
rect 10869 14320 10874 14376
rect 10930 14320 11886 14376
rect 11942 14320 12438 14376
rect 12494 14320 12499 14376
rect 10869 14318 12499 14320
rect 10869 14315 10935 14318
rect 11881 14315 11947 14318
rect 12433 14315 12499 14318
rect 18413 14378 18479 14381
rect 19333 14378 19399 14381
rect 18413 14376 19399 14378
rect 18413 14320 18418 14376
rect 18474 14320 19338 14376
rect 19394 14320 19399 14376
rect 18413 14318 19399 14320
rect 18413 14315 18479 14318
rect 19333 14315 19399 14318
rect 12433 14242 12499 14245
rect 13629 14242 13695 14245
rect 14457 14242 14523 14245
rect 12433 14240 14523 14242
rect 12433 14184 12438 14240
rect 12494 14184 13634 14240
rect 13690 14184 14462 14240
rect 14518 14184 14523 14240
rect 12433 14182 14523 14184
rect 12433 14179 12499 14182
rect 13629 14179 13695 14182
rect 14457 14179 14523 14182
rect 4376 14176 4696 14177
rect 0 14106 800 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 14089 14106 14155 14109
rect 14457 14106 14523 14109
rect 0 14046 1410 14106
rect 0 14016 800 14046
rect 1350 13970 1410 14046
rect 14089 14104 14523 14106
rect 14089 14048 14094 14104
rect 14150 14048 14462 14104
rect 14518 14048 14523 14104
rect 14089 14046 14523 14048
rect 14089 14043 14155 14046
rect 14457 14043 14523 14046
rect 2773 13970 2839 13973
rect 1350 13968 2839 13970
rect 1350 13912 2778 13968
rect 2834 13912 2839 13968
rect 1350 13910 2839 13912
rect 2773 13907 2839 13910
rect 13721 13970 13787 13973
rect 14365 13970 14431 13973
rect 19241 13970 19307 13973
rect 13721 13968 19307 13970
rect 13721 13912 13726 13968
rect 13782 13912 14370 13968
rect 14426 13912 19246 13968
rect 19302 13912 19307 13968
rect 13721 13910 19307 13912
rect 13721 13907 13787 13910
rect 14365 13907 14431 13910
rect 19241 13907 19307 13910
rect 13445 13834 13511 13837
rect 19701 13834 19767 13837
rect 13445 13832 19767 13834
rect 13445 13776 13450 13832
rect 13506 13776 19706 13832
rect 19762 13776 19767 13832
rect 13445 13774 19767 13776
rect 13445 13771 13511 13774
rect 19701 13771 19767 13774
rect 0 13698 800 13728
rect 1761 13698 1827 13701
rect 0 13696 1827 13698
rect 0 13640 1766 13696
rect 1822 13640 1827 13696
rect 0 13638 1827 13640
rect 0 13608 800 13638
rect 1761 13635 1827 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 13261 13426 13327 13429
rect 18045 13426 18111 13429
rect 13261 13424 18111 13426
rect 13261 13368 13266 13424
rect 13322 13368 18050 13424
rect 18106 13368 18111 13424
rect 13261 13366 18111 13368
rect 13261 13363 13327 13366
rect 18045 13363 18111 13366
rect 0 13290 800 13320
rect 5533 13290 5599 13293
rect 0 13288 5599 13290
rect 0 13232 5538 13288
rect 5594 13232 5599 13288
rect 0 13230 5599 13232
rect 0 13200 800 13230
rect 5533 13227 5599 13230
rect 13721 13290 13787 13293
rect 15009 13290 15075 13293
rect 15193 13290 15259 13293
rect 13721 13288 15259 13290
rect 13721 13232 13726 13288
rect 13782 13232 15014 13288
rect 15070 13232 15198 13288
rect 15254 13232 15259 13288
rect 13721 13230 15259 13232
rect 13721 13227 13787 13230
rect 15009 13227 15075 13230
rect 15193 13227 15259 13230
rect 14222 13092 14228 13156
rect 14292 13154 14298 13156
rect 14457 13154 14523 13157
rect 14292 13152 14523 13154
rect 14292 13096 14462 13152
rect 14518 13096 14523 13152
rect 14292 13094 14523 13096
rect 14292 13092 14298 13094
rect 14457 13091 14523 13094
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 11646 12956 11652 13020
rect 11716 13018 11722 13020
rect 11789 13018 11855 13021
rect 11716 13016 11855 13018
rect 11716 12960 11794 13016
rect 11850 12960 11855 13016
rect 11716 12958 11855 12960
rect 11716 12956 11722 12958
rect 11789 12955 11855 12958
rect 0 12746 800 12776
rect 8753 12746 8819 12749
rect 0 12744 8819 12746
rect 0 12688 8758 12744
rect 8814 12688 8819 12744
rect 0 12686 8819 12688
rect 0 12656 800 12686
rect 8753 12683 8819 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 800 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 800 12278
rect 4061 12275 4127 12278
rect 11830 12140 11836 12204
rect 11900 12202 11906 12204
rect 12433 12202 12499 12205
rect 11900 12200 12499 12202
rect 11900 12144 12438 12200
rect 12494 12144 12499 12200
rect 11900 12142 12499 12144
rect 11900 12140 11906 12142
rect 12433 12139 12499 12142
rect 13302 12140 13308 12204
rect 13372 12202 13378 12204
rect 13445 12202 13511 12205
rect 13372 12200 13511 12202
rect 13372 12144 13450 12200
rect 13506 12144 13511 12200
rect 13372 12142 13511 12144
rect 13372 12140 13378 12142
rect 13445 12139 13511 12142
rect 11881 12066 11947 12069
rect 13721 12066 13787 12069
rect 17769 12066 17835 12069
rect 11881 12064 17835 12066
rect 11881 12008 11886 12064
rect 11942 12008 13726 12064
rect 13782 12008 17774 12064
rect 17830 12008 17835 12064
rect 11881 12006 17835 12008
rect 11881 12003 11947 12006
rect 13721 12003 13787 12006
rect 17769 12003 17835 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 12157 11930 12223 11933
rect 12157 11928 12266 11930
rect 12157 11872 12162 11928
rect 12218 11872 12266 11928
rect 12157 11867 12266 11872
rect 0 11794 800 11824
rect 4061 11794 4127 11797
rect 0 11792 4127 11794
rect 0 11736 4066 11792
rect 4122 11736 4127 11792
rect 0 11734 4127 11736
rect 0 11704 800 11734
rect 4061 11731 4127 11734
rect 12206 11661 12266 11867
rect 12206 11656 12315 11661
rect 12206 11600 12254 11656
rect 12310 11600 12315 11656
rect 12206 11598 12315 11600
rect 12249 11595 12315 11598
rect 2221 11522 2287 11525
rect 4429 11522 4495 11525
rect 2221 11520 4495 11522
rect 2221 11464 2226 11520
rect 2282 11464 4434 11520
rect 4490 11464 4495 11520
rect 2221 11462 4495 11464
rect 2221 11459 2287 11462
rect 4429 11459 4495 11462
rect 19793 11522 19859 11525
rect 22000 11522 22800 11552
rect 19793 11520 22800 11522
rect 19793 11464 19798 11520
rect 19854 11464 22800 11520
rect 19793 11462 22800 11464
rect 19793 11459 19859 11462
rect 7808 11456 8128 11457
rect 0 11386 800 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 22000 11432 22800 11462
rect 14672 11391 14992 11392
rect 4061 11386 4127 11389
rect 0 11384 4127 11386
rect 0 11328 4066 11384
rect 4122 11328 4127 11384
rect 0 11326 4127 11328
rect 0 11296 800 11326
rect 4061 11323 4127 11326
rect 4376 10912 4696 10913
rect 0 10842 800 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 0 10752 800 10782
rect 4061 10779 4127 10782
rect 7281 10842 7347 10845
rect 8753 10842 8819 10845
rect 7281 10840 8819 10842
rect 7281 10784 7286 10840
rect 7342 10784 8758 10840
rect 8814 10784 8819 10840
rect 7281 10782 8819 10784
rect 7281 10779 7347 10782
rect 8753 10779 8819 10782
rect 7189 10706 7255 10709
rect 8845 10706 8911 10709
rect 7189 10704 8911 10706
rect 7189 10648 7194 10704
rect 7250 10648 8850 10704
rect 8906 10648 8911 10704
rect 7189 10646 8911 10648
rect 7189 10643 7255 10646
rect 8845 10643 8911 10646
rect 11513 10570 11579 10573
rect 15837 10570 15903 10573
rect 11513 10568 15903 10570
rect 11513 10512 11518 10568
rect 11574 10512 15842 10568
rect 15898 10512 15903 10568
rect 11513 10510 15903 10512
rect 11513 10507 11579 10510
rect 15837 10507 15903 10510
rect 0 10434 800 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 800 10374
rect 4061 10371 4127 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 2681 10300 2747 10301
rect 2630 10298 2636 10300
rect 2590 10238 2636 10298
rect 2700 10296 2747 10300
rect 2742 10240 2747 10296
rect 2630 10236 2636 10238
rect 2700 10236 2747 10240
rect 2681 10235 2747 10236
rect 0 10026 800 10056
rect 9305 10026 9371 10029
rect 11697 10028 11763 10029
rect 0 10024 9371 10026
rect 0 9968 9310 10024
rect 9366 9968 9371 10024
rect 0 9966 9371 9968
rect 0 9936 800 9966
rect 9305 9963 9371 9966
rect 11646 9964 11652 10028
rect 11716 10026 11763 10028
rect 11716 10024 11808 10026
rect 11758 9968 11808 10024
rect 11716 9966 11808 9968
rect 11716 9964 11763 9966
rect 11697 9963 11763 9964
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 2037 9754 2103 9757
rect 1902 9752 2103 9754
rect 1902 9696 2042 9752
rect 2098 9696 2103 9752
rect 1902 9694 2103 9696
rect 1761 9618 1827 9621
rect 1902 9618 1962 9694
rect 2037 9691 2103 9694
rect 14181 9754 14247 9757
rect 17769 9754 17835 9757
rect 14181 9752 17835 9754
rect 14181 9696 14186 9752
rect 14242 9696 17774 9752
rect 17830 9696 17835 9752
rect 14181 9694 17835 9696
rect 14181 9691 14247 9694
rect 17769 9691 17835 9694
rect 1761 9616 1962 9618
rect 1761 9560 1766 9616
rect 1822 9560 1962 9616
rect 1761 9558 1962 9560
rect 1761 9555 1827 9558
rect 0 9482 800 9512
rect 7465 9482 7531 9485
rect 0 9480 7531 9482
rect 0 9424 7470 9480
rect 7526 9424 7531 9480
rect 0 9422 7531 9424
rect 0 9392 800 9422
rect 7465 9419 7531 9422
rect 1301 9346 1367 9349
rect 2497 9346 2563 9349
rect 1301 9344 2563 9346
rect 1301 9288 1306 9344
rect 1362 9288 2502 9344
rect 2558 9288 2563 9344
rect 1301 9286 2563 9288
rect 1301 9283 1367 9286
rect 2497 9283 2563 9286
rect 12433 9346 12499 9349
rect 12566 9346 12572 9348
rect 12433 9344 12572 9346
rect 12433 9288 12438 9344
rect 12494 9288 12572 9344
rect 12433 9286 12572 9288
rect 12433 9283 12499 9286
rect 12566 9284 12572 9286
rect 12636 9284 12642 9348
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 1209 9210 1275 9213
rect 5073 9210 5139 9213
rect 1209 9208 5139 9210
rect 1209 9152 1214 9208
rect 1270 9152 5078 9208
rect 5134 9152 5139 9208
rect 1209 9150 5139 9152
rect 1209 9147 1275 9150
rect 5073 9147 5139 9150
rect 0 9074 800 9104
rect 8937 9074 9003 9077
rect 0 9072 9003 9074
rect 0 9016 8942 9072
rect 8998 9016 9003 9072
rect 0 9014 9003 9016
rect 0 8984 800 9014
rect 8937 9011 9003 9014
rect 6269 8938 6335 8941
rect 9213 8938 9279 8941
rect 6269 8936 9279 8938
rect 6269 8880 6274 8936
rect 6330 8880 9218 8936
rect 9274 8880 9279 8936
rect 6269 8878 9279 8880
rect 6269 8875 6335 8878
rect 9213 8875 9279 8878
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 800 8560
rect 4153 8530 4219 8533
rect 0 8528 4219 8530
rect 0 8472 4158 8528
rect 4214 8472 4219 8528
rect 0 8470 4219 8472
rect 0 8440 800 8470
rect 4153 8467 4219 8470
rect 5809 8394 5875 8397
rect 12382 8394 12388 8396
rect 5809 8392 12388 8394
rect 5809 8336 5814 8392
rect 5870 8336 12388 8392
rect 5809 8334 12388 8336
rect 5809 8331 5875 8334
rect 12382 8332 12388 8334
rect 12452 8332 12458 8396
rect 2681 8260 2747 8261
rect 2630 8258 2636 8260
rect 2590 8198 2636 8258
rect 2700 8256 2747 8260
rect 2742 8200 2747 8256
rect 2630 8196 2636 8198
rect 2700 8196 2747 8200
rect 2681 8195 2747 8196
rect 7808 8192 8128 8193
rect 0 8122 800 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 5809 8122 5875 8125
rect 0 8120 5875 8122
rect 0 8064 5814 8120
rect 5870 8064 5875 8120
rect 0 8062 5875 8064
rect 0 8032 800 8062
rect 5809 8059 5875 8062
rect 2957 7852 3023 7853
rect 2957 7850 3004 7852
rect 2912 7848 3004 7850
rect 2912 7792 2962 7848
rect 2912 7790 3004 7792
rect 2957 7788 3004 7790
rect 3068 7788 3074 7852
rect 2957 7787 3023 7788
rect 4376 7648 4696 7649
rect 0 7578 800 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 4061 7578 4127 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7488 800 7518
rect 4061 7515 4127 7518
rect 7833 7442 7899 7445
rect 4110 7440 7899 7442
rect 4110 7384 7838 7440
rect 7894 7384 7899 7440
rect 4110 7382 7899 7384
rect 2865 7306 2931 7309
rect 2998 7306 3004 7308
rect 2865 7304 3004 7306
rect 2865 7248 2870 7304
rect 2926 7248 3004 7304
rect 2865 7246 3004 7248
rect 2865 7243 2931 7246
rect 2998 7244 3004 7246
rect 3068 7244 3074 7308
rect 0 7170 800 7200
rect 4110 7170 4170 7382
rect 7833 7379 7899 7382
rect 4337 7306 4403 7309
rect 9581 7306 9647 7309
rect 4337 7304 9647 7306
rect 4337 7248 4342 7304
rect 4398 7248 9586 7304
rect 9642 7248 9647 7304
rect 4337 7246 9647 7248
rect 4337 7243 4403 7246
rect 9581 7243 9647 7246
rect 0 7110 4170 7170
rect 0 7080 800 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 0 6762 800 6792
rect 8293 6762 8359 6765
rect 0 6760 8359 6762
rect 0 6704 8298 6760
rect 8354 6704 8359 6760
rect 0 6702 8359 6704
rect 0 6672 800 6702
rect 8293 6699 8359 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 6085 6354 6151 6357
rect 7925 6354 7991 6357
rect 6085 6352 7991 6354
rect 6085 6296 6090 6352
rect 6146 6296 7930 6352
rect 7986 6296 7991 6352
rect 6085 6294 7991 6296
rect 6085 6291 6151 6294
rect 7925 6291 7991 6294
rect 0 6218 800 6248
rect 7833 6218 7899 6221
rect 0 6216 7899 6218
rect 0 6160 7838 6216
rect 7894 6160 7899 6216
rect 0 6158 7899 6160
rect 0 6128 800 6158
rect 7833 6155 7899 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 800 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 800 5750
rect 4061 5747 4127 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 800 5296
rect 3969 5266 4035 5269
rect 0 5264 4035 5266
rect 0 5208 3974 5264
rect 4030 5208 4035 5264
rect 0 5206 4035 5208
rect 0 5176 800 5206
rect 3969 5203 4035 5206
rect 7808 4928 8128 4929
rect 0 4858 800 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 800 4798
rect 4061 4795 4127 4798
rect 4376 4384 4696 4385
rect 0 4314 800 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 0 4254 4308 4314
rect 0 4224 800 4254
rect 4248 4178 4308 4254
rect 13302 4178 13308 4180
rect 4248 4118 13308 4178
rect 13302 4116 13308 4118
rect 13372 4116 13378 4180
rect 0 3906 800 3936
rect 3969 3906 4035 3909
rect 0 3904 4035 3906
rect 0 3848 3974 3904
rect 4030 3848 4035 3904
rect 0 3846 4035 3848
rect 0 3816 800 3846
rect 3969 3843 4035 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 0 3498 800 3528
rect 2865 3498 2931 3501
rect 0 3496 2931 3498
rect 0 3440 2870 3496
rect 2926 3440 2931 3496
rect 0 3438 2931 3440
rect 0 3408 800 3438
rect 2865 3435 2931 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 800 2984
rect 1209 2954 1275 2957
rect 0 2952 1275 2954
rect 0 2896 1214 2952
rect 1270 2896 1275 2952
rect 0 2894 1275 2896
rect 0 2864 800 2894
rect 1209 2891 1275 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 800 2576
rect 4245 2546 4311 2549
rect 0 2544 4311 2546
rect 0 2488 4250 2544
rect 4306 2488 4311 2544
rect 0 2486 4311 2488
rect 0 2456 800 2486
rect 4245 2483 4311 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 800 2032
rect 4797 2002 4863 2005
rect 0 2000 4863 2002
rect 0 1944 4802 2000
rect 4858 1944 4863 2000
rect 0 1942 4863 1944
rect 0 1912 800 1942
rect 4797 1939 4863 1942
rect 0 1594 800 1624
rect 5073 1594 5139 1597
rect 0 1592 5139 1594
rect 0 1536 5078 1592
rect 5134 1536 5139 1592
rect 0 1534 5139 1536
rect 0 1504 800 1534
rect 5073 1531 5139 1534
rect 0 1050 800 1080
rect 1025 1050 1091 1053
rect 0 1048 1091 1050
rect 0 992 1030 1048
rect 1086 992 1091 1048
rect 0 990 1091 992
rect 0 960 800 990
rect 1025 987 1091 990
rect 0 642 800 672
rect 1117 642 1183 645
rect 0 640 1183 642
rect 0 584 1122 640
rect 1178 584 1183 640
rect 0 582 1183 584
rect 0 552 800 582
rect 1117 579 1183 582
rect 0 234 800 264
rect 3877 234 3943 237
rect 0 232 3943 234
rect 0 176 3882 232
rect 3938 176 3943 232
rect 0 174 3943 176
rect 0 144 800 174
rect 3877 171 3943 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 14228 19076 14292 19140
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 11652 19000 11716 19004
rect 11652 18944 11666 19000
rect 11666 18944 11716 19000
rect 11652 18940 11716 18944
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 12572 18396 12636 18460
rect 12388 18048 12452 18052
rect 12388 17992 12438 18048
rect 12438 17992 12452 18048
rect 12388 17988 12452 17992
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 14228 13092 14292 13156
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 11652 12956 11716 13020
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 11836 12140 11900 12204
rect 13308 12140 13372 12204
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 2636 10296 2700 10300
rect 2636 10240 2686 10296
rect 2686 10240 2700 10296
rect 2636 10236 2700 10240
rect 11652 10024 11716 10028
rect 11652 9968 11702 10024
rect 11702 9968 11716 10024
rect 11652 9964 11716 9968
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 12572 9284 12636 9348
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 12388 8332 12452 8396
rect 2636 8256 2700 8260
rect 2636 8200 2686 8256
rect 2686 8200 2700 8256
rect 2636 8196 2700 8200
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 3004 7848 3068 7852
rect 3004 7792 3018 7848
rect 3018 7792 3068 7848
rect 3004 7788 3068 7792
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 3004 7244 3068 7308
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 13308 4116 13372 4180
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 2635 10300 2701 10301
rect 2635 10236 2636 10300
rect 2700 10236 2701 10300
rect 2635 10235 2701 10236
rect 2638 8261 2698 10235
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 2635 8260 2701 8261
rect 2635 8196 2636 8260
rect 2700 8196 2701 8260
rect 2635 8195 2701 8196
rect 3003 7852 3069 7853
rect 3003 7788 3004 7852
rect 3068 7788 3069 7852
rect 3003 7787 3069 7788
rect 3006 7309 3066 7787
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 3003 7308 3069 7309
rect 3003 7244 3004 7308
rect 3068 7244 3069 7308
rect 3003 7243 3069 7244
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14227 19140 14293 19141
rect 14227 19076 14228 19140
rect 14292 19076 14293 19140
rect 14227 19075 14293 19076
rect 11651 19004 11717 19005
rect 11651 18940 11652 19004
rect 11716 18940 11717 19004
rect 11651 18939 11717 18940
rect 11654 18730 11714 18939
rect 11654 18670 11898 18730
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11651 13020 11717 13021
rect 11651 12956 11652 13020
rect 11716 12956 11717 13020
rect 11651 12955 11717 12956
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11654 10029 11714 12955
rect 11838 12205 11898 18670
rect 12571 18460 12637 18461
rect 12571 18396 12572 18460
rect 12636 18396 12637 18460
rect 12571 18395 12637 18396
rect 12387 18052 12453 18053
rect 12387 17988 12388 18052
rect 12452 17988 12453 18052
rect 12387 17987 12453 17988
rect 11835 12204 11901 12205
rect 11835 12140 11836 12204
rect 11900 12140 11901 12204
rect 11835 12139 11901 12140
rect 11651 10028 11717 10029
rect 11651 9964 11652 10028
rect 11716 9964 11717 10028
rect 11651 9963 11717 9964
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 12390 8397 12450 17987
rect 12574 9349 12634 18395
rect 14230 13157 14290 19075
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14227 13156 14293 13157
rect 14227 13092 14228 13156
rect 14292 13092 14293 13156
rect 14227 13091 14293 13092
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 13307 12204 13373 12205
rect 13307 12140 13308 12204
rect 13372 12140 13373 12204
rect 13307 12139 13373 12140
rect 12571 9348 12637 9349
rect 12571 9284 12572 9348
rect 12636 9284 12637 9348
rect 12571 9283 12637 9284
rect 12387 8396 12453 8397
rect 12387 8332 12388 8396
rect 12452 8332 12453 8396
rect 12387 8331 12453 8332
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 13310 4181 13370 12139
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 13307 4180 13373 4181
rect 13307 4116 13308 4180
rect 13372 4116 13373 4180
rect 13307 4115 13373 4116
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608762952
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608762952
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1608762952
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1608762952
transform 1 0 20792 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1608762952
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_216
timestamp 1608762952
transform 1 0 20976 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1608762952
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608762952
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608762952
transform 1 0 19688 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1608762952
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1608762952
transform 1 0 19228 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1608762952
transform 1 0 19596 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_204
timestamp 1608762952
transform 1 0 19872 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_208
timestamp 1608762952
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608762952
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608762952
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_183
timestamp 1608762952
transform 1 0 17940 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 17756 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_179
timestamp 1608762952
transform 1 0 17572 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608762952
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1608762952
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1608762952
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1608762952
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608762952
transform 1 0 16100 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 15640 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_156
timestamp 1608762952
transform 1 0 15456 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_160
timestamp 1608762952
transform 1 0 15824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608762952
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1608762952
transform 1 0 15088 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1608762952
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 14720 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_146
timestamp 1608762952
transform 1 0 14536 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_150
timestamp 1608762952
transform 1 0 14904 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608762952
transform 1 0 13248 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608762952
transform 1 0 13800 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_129
timestamp 1608762952
transform 1 0 12972 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_136
timestamp 1608762952
transform 1 0 13616 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_142
timestamp 1608762952
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608762952
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1608762952
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_121
timestamp 1608762952
transform 1 0 12236 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1608762952
transform 1 0 12052 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1608762952
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 11684 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_113
timestamp 1608762952
transform 1 0 11500 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_109
timestamp 1608762952
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608762952
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_105
timestamp 1608762952
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_101
timestamp 1608762952
transform 1 0 10396 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1608762952
transform 1 0 9752 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1608762952
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608762952
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 9292 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1608762952
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_84
timestamp 1608762952
transform 1 0 8832 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_88
timestamp 1608762952
transform 1 0 9200 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_80
timestamp 1608762952
transform 1 0 8464 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_76
timestamp 1608762952
transform 1 0 8096 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 7912 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_71
timestamp 1608762952
transform 1 0 7636 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_67
timestamp 1608762952
transform 1 0 7268 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1608762952
transform 1 0 7084 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp 1608762952
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608762952
transform 1 0 5244 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608762952
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 6256 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_54
timestamp 1608762952
transform 1 0 6072 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_58
timestamp 1608762952
transform 1 0 6440 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608762952
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608762952
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_26
timestamp 1608762952
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1608762952
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608762952
transform 1 0 1472 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 2024 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608762952
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1608762952
transform 1 0 1380 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_8
timestamp 1608762952
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_16
timestamp 1608762952
transform 1 0 2576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_20
timestamp 1608762952
transform 1 0 2944 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608762952
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_213
timestamp 1608762952
transform 1 0 20700 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_217
timestamp 1608762952
transform 1 0 21068 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608762952
transform 1 0 18768 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608762952
transform 1 0 19596 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_190
timestamp 1608762952
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_196
timestamp 1608762952
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_200
timestamp 1608762952
transform 1 0 19504 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 16928 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608762952
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1608762952
transform 1 0 17664 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_170
timestamp 1608762952
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_178
timestamp 1608762952
transform 1 0 17480 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1608762952
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608762952
transform 1 0 14720 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608762952
transform 1 0 15272 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608762952
transform 1 0 15824 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608762952
transform 1 0 16376 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1608762952
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_152
timestamp 1608762952
transform 1 0 15088 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_158
timestamp 1608762952
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_164
timestamp 1608762952
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608762952
transform 1 0 13616 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608762952
transform 1 0 14168 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 12880 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_134
timestamp 1608762952
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_140
timestamp 1608762952
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 11592 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608762952
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_112
timestamp 1608762952
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1608762952
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_123
timestamp 1608762952
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 9936 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608762952
transform 1 0 8924 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_94
timestamp 1608762952
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1608762952
transform 1 0 7912 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 7728 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1608762952
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1608762952
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_83
timestamp 1608762952
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 5060 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608762952
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608762952
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1608762952
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 3036 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_37
timestamp 1608762952
transform 1 0 4508 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608762952
transform 1 0 1472 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 2024 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608762952
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1608762952
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1608762952
transform 1 0 1380 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_8
timestamp 1608762952
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_16
timestamp 1608762952
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_20
timestamp 1608762952
transform 1 0 2944 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608762952
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608762952
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1608762952
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1608762952
transform 1 0 21068 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_210
timestamp 1608762952
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1608762952
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1608762952
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 18400 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 19136 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1608762952
transform 1 0 19504 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1608762952
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1608762952
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1608762952
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1608762952
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1608762952
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_206
timestamp 1608762952
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 16744 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 17664 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 17480 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_168
timestamp 1608762952
transform 1 0 16560 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1608762952
transform 1 0 17296 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_186
timestamp 1608762952
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 16008 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608762952
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_146
timestamp 1608762952
transform 1 0 14536 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_150
timestamp 1608762952
transform 1 0 14904 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_160
timestamp 1608762952
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 13248 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1608762952
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1608762952
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_130
timestamp 1608762952
transform 1 0 13064 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1608762952
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1608762952
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 12512 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 11776 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_111
timestamp 1608762952
transform 1 0 11316 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1608762952
transform 1 0 11684 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_122
timestamp 1608762952
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 9844 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608762952
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_86
timestamp 1608762952
transform 1 0 9016 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1608762952
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1608762952
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1608762952
transform 1 0 7084 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 7544 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_68
timestamp 1608762952
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 5336 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_62
timestamp 1608762952
transform 1 0 6808 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1608762952
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608762952
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_28
timestamp 1608762952
transform 1 0 3680 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_41
timestamp 1608762952
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608762952
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 1932 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1608762952
transform 1 0 2852 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608762952
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1608762952
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_15
timestamp 1608762952
transform 1 0 2484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608762952
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20516 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1608762952
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_213
timestamp 1608762952
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_217
timestamp 1608762952
transform 1 0 21068 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20148 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_205
timestamp 1608762952
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1608762952
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 1608762952
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1608762952
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1608762952
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 1608762952
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608762952
transform 1 0 18124 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 17112 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608762952
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_171
timestamp 1608762952
transform 1 0 16836 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1608762952
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1608762952
transform 1 0 18032 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608762952
transform 1 0 14996 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1608762952
transform 1 0 16008 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_147
timestamp 1608762952
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1608762952
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608762952
transform 1 0 13432 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1608762952
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1608762952
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608762952
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608762952
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1608762952
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1608762952
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1608762952
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1608762952
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1608762952
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 9752 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_92
timestamp 1608762952
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608762952
transform 1 0 8740 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1608762952
transform 1 0 7544 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_68
timestamp 1608762952
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_79
timestamp 1608762952
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1608762952
transform 1 0 5520 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608762952
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_43
timestamp 1608762952
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_47
timestamp 1608762952
transform 1 0 5428 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1608762952
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608762952
transform 1 0 4416 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_33
timestamp 1608762952
transform 1 0 4140 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_39
timestamp 1608762952
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608762952
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 2668 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608762952
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1608762952
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_11
timestamp 1608762952
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608762952
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608762952
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20332 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1608762952
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1608762952
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1608762952
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1608762952
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_207
timestamp 1608762952
transform 1 0 20148 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1608762952
transform 1 0 19964 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_203
timestamp 1608762952
transform 1 0 19780 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1608762952
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1608762952
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_199
timestamp 1608762952
transform 1 0 19412 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_195
timestamp 1608762952
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608762952
transform 1 0 18400 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_191
timestamp 1608762952
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1608762952
transform 1 0 17388 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 16928 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1608762952
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_174
timestamp 1608762952
transform 1 0 17112 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1608762952
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 15272 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608762952
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1608762952
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608762952
transform 1 0 13616 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608762952
transform 1 0 14168 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_134
timestamp 1608762952
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_139
timestamp 1608762952
transform 1 0 13892 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762952
transform 1 0 11960 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608762952
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1608762952
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_106
timestamp 1608762952
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_110
timestamp 1608762952
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_114
timestamp 1608762952
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1608762952
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608762952
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_86
timestamp 1608762952
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1608762952
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1608762952
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 8464 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1608762952
transform 1 0 7084 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 1608762952
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_72
timestamp 1608762952
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1608762952
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 5244 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_43
timestamp 1608762952
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1608762952
transform 1 0 6716 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608762952
transform 1 0 4784 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608762952
transform 1 0 3404 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608762952
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1608762952
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_28
timestamp 1608762952
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1608762952
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_36
timestamp 1608762952
transform 1 0 4416 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608762952
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608762952
transform 1 0 2300 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608762952
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608762952
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1608762952
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1608762952
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1608762952
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608762952
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608762952
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1608762952
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1608762952
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608762952
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1608762952
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_216
timestamp 1608762952
transform 1 0 20976 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1608762952
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1608762952
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1608762952
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_208
timestamp 1608762952
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1608762952
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_204
timestamp 1608762952
transform 1 0 19872 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_204
timestamp 1608762952
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_200
timestamp 1608762952
transform 1 0 19504 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_200
timestamp 1608762952
transform 1 0 19504 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 18032 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 18032 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1608762952
transform 1 0 16928 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608762952
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_182
timestamp 1608762952
transform 1 0 17848 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_168
timestamp 1608762952
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1608762952
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 16376 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 14628 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 16192 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_159
timestamp 1608762952
transform 1 0 15732 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_163
timestamp 1608762952
transform 1 0 16100 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_163
timestamp 1608762952
transform 1 0 16100 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608762952
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_147
timestamp 1608762952
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1608762952
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1608762952
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 12696 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608762952
transform 1 0 13432 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_132
timestamp 1608762952
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_143
timestamp 1608762952
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_142
timestamp 1608762952
transform 1 0 14168 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608762952
transform 1 0 12420 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608762952
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_121
timestamp 1608762952
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1608762952
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_123
timestamp 1608762952
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608762952
transform 1 0 11408 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_106
timestamp 1608762952
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_110
timestamp 1608762952
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1608762952
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_112
timestamp 1608762952
transform 1 0 11408 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 9568 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1608762952
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1608762952
transform 1 0 9108 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1608762952
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608762952
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1608762952
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1608762952
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 7268 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1608762952
transform 1 0 7452 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 8464 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_63
timestamp 1608762952
transform 1 0 6900 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_78
timestamp 1608762952
transform 1 0 8280 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_83
timestamp 1608762952
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1608762952
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_62
timestamp 1608762952
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 6348 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608762952
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 6164 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_53
timestamp 1608762952
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1608762952
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1608762952
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1608762952
transform 1 0 5244 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1608762952
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 5704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_48
timestamp 1608762952
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1608762952
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608762952
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_28
timestamp 1608762952
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1608762952
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_36
timestamp 1608762952
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_40
timestamp 1608762952
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 2944 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1608762952
transform 1 0 2852 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 2116 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_17
timestamp 1608762952
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1608762952
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608762952
transform 1 0 1564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608762952
transform 1 0 1472 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 2024 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608762952
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608762952
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1608762952
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_9
timestamp 1608762952
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1608762952
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1608762952
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608762952
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1608762952
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_213
timestamp 1608762952
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_217
timestamp 1608762952
transform 1 0 21068 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1608762952
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_197
timestamp 1608762952
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_201
timestamp 1608762952
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_205
timestamp 1608762952
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1608762952
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608762952
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_168
timestamp 1608762952
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1608762952
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1608762952
transform 1 0 17296 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_180
timestamp 1608762952
transform 1 0 17664 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 14904 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 15916 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1608762952
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_153
timestamp 1608762952
transform 1 0 15180 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1608762952
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_164
timestamp 1608762952
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608762952
transform 1 0 12788 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 13248 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_130
timestamp 1608762952
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608762952
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1608762952
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1608762952
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1608762952
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 8924 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762952
transform 1 0 10672 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_101
timestamp 1608762952
transform 1 0 10396 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 7084 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 1608762952
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608762952
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1608762952
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1608762952
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 4876 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_33
timestamp 1608762952
transform 1 0 4140 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_38
timestamp 1608762952
transform 1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608762952
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 2668 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 1932 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608762952
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1608762952
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1608762952
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608762952
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608762952
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1608762952
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1608762952
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1608762952
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608762952
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608762952
transform 1 0 18860 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 19320 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1608762952
transform 1 0 19688 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1608762952
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_191
timestamp 1608762952
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_196
timestamp 1608762952
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_200
timestamp 1608762952
transform 1 0 19504 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_204
timestamp 1608762952
transform 1 0 19872 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_208
timestamp 1608762952
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608762952
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1608762952
transform 1 0 17848 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 17296 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_169
timestamp 1608762952
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_174
timestamp 1608762952
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_178
timestamp 1608762952
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608762952
transform 1 0 15824 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608762952
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 14904 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_148
timestamp 1608762952
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1608762952
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1608762952
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1608762952
transform 1 0 15640 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1608762952
transform 1 0 13524 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1608762952
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 1608762952
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 10764 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1608762952
transform 1 0 12512 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_121
timestamp 1608762952
transform 1 0 12236 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1608762952
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608762952
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1608762952
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_102
timestamp 1608762952
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1608762952
transform 1 0 7912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1608762952
transform 1 0 8556 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1608762952
transform 1 0 6900 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_72
timestamp 1608762952
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_77
timestamp 1608762952
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1608762952
transform 1 0 5612 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_47
timestamp 1608762952
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_58
timestamp 1608762952
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_62
timestamp 1608762952
transform 1 0 6808 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608762952
transform 1 0 3220 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1608762952
transform 1 0 4600 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608762952
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 3680 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1608762952
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1608762952
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1608762952
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1608762952
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 2300 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_15
timestamp 1608762952
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1608762952
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1608762952
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1608762952
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608762952
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1608762952
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608762952
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_210
timestamp 1608762952
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_214
timestamp 1608762952
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1608762952
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 20240 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_202
timestamp 1608762952
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_206
timestamp 1608762952
transform 1 0 20056 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 18216 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608762952
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1608762952
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1608762952
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1608762952
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 15732 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_153
timestamp 1608762952
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1608762952
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1608762952
transform 1 0 14352 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 13984 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1608762952
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_134
timestamp 1608762952
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1608762952
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_143
timestamp 1608762952
transform 1 0 14260 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608762952
transform 1 0 12604 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1608762952
transform 1 0 11316 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608762952
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_106
timestamp 1608762952
transform 1 0 10856 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608762952
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1608762952
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 10672 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1608762952
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_102
timestamp 1608762952
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 8648 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 7084 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_68
timestamp 1608762952
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_72
timestamp 1608762952
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1608762952
transform 1 0 8096 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608762952
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_56
timestamp 1608762952
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1608762952
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1608762952
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 4784 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_35
timestamp 1608762952
transform 1 0 4324 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608762952
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 2852 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 1932 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608762952
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1608762952
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_15
timestamp 1608762952
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608762952
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608762952
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1608762952
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1608762952
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1608762952
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1608762952
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1608762952
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 18400 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_204
timestamp 1608762952
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1608762952
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608762952
transform 1 0 17572 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1608762952
transform 1 0 16560 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_177
timestamp 1608762952
transform 1 0 17388 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_182
timestamp 1608762952
transform 1 0 17848 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608762952
transform 1 0 15548 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608762952
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 1608762952
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1608762952
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1608762952
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_166
timestamp 1608762952
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608762952
transform 1 0 13800 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608762952
transform 1 0 12788 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_136
timestamp 1608762952
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1608762952
transform 1 0 11408 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_108
timestamp 1608762952
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_121
timestamp 1608762952
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_125
timestamp 1608762952
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1608762952
transform 1 0 9016 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608762952
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1608762952
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1608762952
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1608762952
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1608762952
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_99
timestamp 1608762952
transform 1 0 10212 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_104
timestamp 1608762952
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_76
timestamp 1608762952
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1608762952
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 6624 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 5704 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1608762952
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_49
timestamp 1608762952
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1608762952
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1608762952
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1608762952
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608762952
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1608762952
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1608762952
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608762952
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 1932 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1608762952
transform 1 0 2944 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608762952
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1608762952
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_15
timestamp 1608762952
transform 1 0 2484 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608762952
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_209
timestamp 1608762952
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_213
timestamp 1608762952
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1608762952
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20148 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1608762952
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1608762952
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_201
timestamp 1608762952
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_205
timestamp 1608762952
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1608762952
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608762952
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1608762952
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 16284 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_156
timestamp 1608762952
transform 1 0 15456 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_160
timestamp 1608762952
transform 1 0 15824 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_163
timestamp 1608762952
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762952
transform 1 0 13984 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608762952
transform 1 0 12972 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1608762952
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_138
timestamp 1608762952
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608762952
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1608762952
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1608762952
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 10580 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1608762952
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1608762952
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1608762952
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 8372 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1608762952
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_76
timestamp 1608762952
transform 1 0 8096 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1608762952
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1608762952
transform 1 0 5704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608762952
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_46
timestamp 1608762952
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1608762952
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608762952
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 3864 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_26
timestamp 1608762952
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608762952
transform 1 0 1564 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 2116 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608762952
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1608762952
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1608762952
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_17
timestamp 1608762952
transform 1 0 2668 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608762952
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608762952
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1608762952
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608762952
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608762952
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_213
timestamp 1608762952
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1608762952
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1608762952
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1608762952
transform 1 0 20516 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_209
timestamp 1608762952
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_209
timestamp 1608762952
transform 1 0 20332 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1608762952
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 20148 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_205
timestamp 1608762952
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_205
timestamp 1608762952
transform 1 0 19964 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1608762952
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1608762952
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_201
timestamp 1608762952
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_201
timestamp 1608762952
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1608762952
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1608762952
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1608762952
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1608762952
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1608762952
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 17020 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608762952
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608762952
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1608762952
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1608762952
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608762952
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_168
timestamp 1608762952
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1608762952
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_176
timestamp 1608762952
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_167
timestamp 1608762952
transform 1 0 16468 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1608762952
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_164
timestamp 1608762952
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1608762952
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 15916 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1608762952
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1608762952
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_158
timestamp 1608762952
transform 1 0 15640 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1608762952
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1608762952
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1608762952
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608762952
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1608762952
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1608762952
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608762952
transform 1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_147
timestamp 1608762952
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_148
timestamp 1608762952
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 13248 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608762952
transform 1 0 13800 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 13432 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1608762952
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_137
timestamp 1608762952
transform 1 0 13708 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_131
timestamp 1608762952
transform 1 0 13156 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1608762952
transform 1 0 12328 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1608762952
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608762952
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1608762952
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762952
transform 1 0 10672 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 10488 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608762952
transform 1 0 10028 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1608762952
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_97
timestamp 1608762952
transform 1 0 10028 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_101
timestamp 1608762952
transform 1 0 10396 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_100
timestamp 1608762952
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608762952
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1608762952
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1608762952
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1608762952
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1608762952
transform 1 0 7728 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 8188 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1608762952
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 8280 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_68
timestamp 1608762952
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1608762952
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_76
timestamp 1608762952
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1608762952
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 6624 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608762952
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1608762952
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1608762952
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1608762952
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_57
timestamp 1608762952
transform 1 0 6348 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 4508 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 4876 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_35
timestamp 1608762952
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1608762952
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_38
timestamp 1608762952
transform 1 0 4600 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1608762952
transform 1 0 3496 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608762952
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1608762952
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1608762952
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1608762952
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_16
timestamp 1608762952
transform 1 0 2576 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1608762952
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_19
timestamp 1608762952
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 1932 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 2024 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_8
timestamp 1608762952
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1608762952
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608762952
transform 1 0 1472 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608762952
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608762952
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608762952
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1608762952
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608762952
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608762952
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1608762952
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1608762952
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1608762952
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1608762952
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608762952
transform 1 0 18492 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 19136 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1608762952
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608762952
transform 1 0 17480 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_172
timestamp 1608762952
transform 1 0 16928 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1608762952
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 15456 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608762952
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1608762952
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1608762952
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1608762952
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1608762952
transform 1 0 13708 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1608762952
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_130
timestamp 1608762952
transform 1 0 13064 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_134
timestamp 1608762952
transform 1 0 13432 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 11592 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_108
timestamp 1608762952
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_112
timestamp 1608762952
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1608762952
transform 1 0 10212 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608762952
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_86
timestamp 1608762952
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1608762952
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1608762952
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1608762952
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1608762952
transform 1 0 8188 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 7544 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1608762952
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_73
timestamp 1608762952
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 5888 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1608762952
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608762952
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1608762952
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1608762952
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608762952
transform 1 0 1564 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608762952
transform 1 0 2852 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 2116 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608762952
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1608762952
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_9
timestamp 1608762952
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_17
timestamp 1608762952
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608762952
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 20424 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608762952
transform 1 0 20792 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1608762952
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1608762952
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1608762952
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_204
timestamp 1608762952
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_208
timestamp 1608762952
transform 1 0 20240 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 18032 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1608762952
transform 1 0 16560 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608762952
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_177
timestamp 1608762952
transform 1 0 17388 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 14904 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_147
timestamp 1608762952
transform 1 0 14628 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1608762952
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608762952
transform 1 0 13248 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 14076 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1608762952
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608762952
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1608762952
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 10212 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1608762952
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1608762952
transform 1 0 9660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 7820 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1608762952
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608762952
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1608762952
transform 1 0 5428 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608762952
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_45
timestamp 1608762952
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_56
timestamp 1608762952
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1608762952
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608762952
transform 1 0 4416 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 1608762952
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 2760 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 1932 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608762952
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1608762952
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1608762952
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1608762952
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_15
timestamp 1608762952
transform 1 0 2484 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608762952
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608762952
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1608762952
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1608762952
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1608762952
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_207
timestamp 1608762952
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_203
timestamp 1608762952
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1608762952
transform 1 0 19412 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_195
timestamp 1608762952
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_191
timestamp 1608762952
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1608762952
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 16744 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1608762952
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_173
timestamp 1608762952
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_177
timestamp 1608762952
transform 1 0 17388 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1608762952
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608762952
transform 1 0 16284 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1608762952
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608762952
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1608762952
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1608762952
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1608762952
transform 1 0 13156 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1608762952
transform 1 0 14168 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1608762952
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_140
timestamp 1608762952
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608762952
transform 1 0 11960 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_105
timestamp 1608762952
transform 1 0 10764 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_111
timestamp 1608762952
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_115
timestamp 1608762952
transform 1 0 11684 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608762952
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1608762952
transform 1 0 10396 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1608762952
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608762952
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1608762952
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608762952
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_86
timestamp 1608762952
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 7544 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1608762952
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1608762952
transform 1 0 5244 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608762952
transform 1 0 6532 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 5704 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp 1608762952
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1608762952
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_53
timestamp 1608762952
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_57
timestamp 1608762952
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608762952
transform 1 0 4232 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608762952
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1608762952
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1608762952
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1608762952
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608762952
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 1748 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608762952
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1608762952
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1608762952
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_13
timestamp 1608762952
transform 1 0 2300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1608762952
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608762952
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_212
timestamp 1608762952
transform 1 0 20608 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1608762952
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_204
timestamp 1608762952
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_208
timestamp 1608762952
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608762952
transform 1 0 17388 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608762952
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1608762952
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1608762952
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 15732 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1608762952
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 14076 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_139
timestamp 1608762952
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608762952
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1608762952
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608762952
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_114
timestamp 1608762952
transform 1 0 11592 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1608762952
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1608762952
transform 1 0 9476 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1608762952
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1608762952
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_104
timestamp 1608762952
transform 1 0 10672 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608762952
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1608762952
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608762952
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_54
timestamp 1608762952
transform 1 0 6072 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1608762952
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_42
timestamp 1608762952
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_46
timestamp 1608762952
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_50
timestamp 1608762952
transform 1 0 5704 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608762952
transform 1 0 3404 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1608762952
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_24
timestamp 1608762952
transform 1 0 3312 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1608762952
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_38
timestamp 1608762952
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608762952
transform 1 0 2116 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608762952
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1608762952
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_20
timestamp 1608762952
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608762952
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608762952
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608762952
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1608762952
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1608762952
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1608762952
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1608762952
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_198
timestamp 1608762952
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_202
timestamp 1608762952
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1608762952
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1608762952
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_192
timestamp 1608762952
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1608762952
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1608762952
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608762952
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_177
timestamp 1608762952
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1608762952
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1608762952
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_182
timestamp 1608762952
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_186
timestamp 1608762952
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1608762952
transform 1 0 16560 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 16376 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1608762952
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_164
timestamp 1608762952
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_164
timestamp 1608762952
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1608762952
transform 1 0 15364 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608762952
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_155
timestamp 1608762952
transform 1 0 15364 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1608762952
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1608762952
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1608762952
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1608762952
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608762952
transform 1 0 14352 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 13340 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1608762952
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_132
timestamp 1608762952
transform 1 0 13248 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1608762952
transform 1 0 13708 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_143
timestamp 1608762952
transform 1 0 14260 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_131
timestamp 1608762952
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 11684 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1608762952
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608762952
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_117
timestamp 1608762952
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1608762952
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1608762952
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1608762952
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_113
timestamp 1608762952
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 10028 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1608762952
transform 1 0 10304 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_98
timestamp 1608762952
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608762952
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1608762952
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1608762952
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1608762952
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 8648 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608762952
transform 1 0 8096 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1608762952
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1608762952
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_75
timestamp 1608762952
transform 1 0 8004 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_79
timestamp 1608762952
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk
timestamp 1608762952
transform 1 0 7728 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1608762952
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1608762952
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_66
timestamp 1608762952
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_70
timestamp 1608762952
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762952
transform 1 0 5704 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1608762952
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1608762952
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608762952
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1608762952
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1608762952
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608762952
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_48
timestamp 1608762952
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608762952
transform 1 0 3496 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608762952
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608762952
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_24
timestamp 1608762952
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1608762952
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1608762952
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762952
transform 1 0 1840 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608762952
transform 1 0 2852 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_17
timestamp 1608762952
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608762952
transform 1 0 1840 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608762952
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608762952
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1608762952
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608762952
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1608762952
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1608762952
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608762952
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608762952
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1608762952
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1608762952
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1608762952
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_198
timestamp 1608762952
transform 1 0 19320 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_168
timestamp 1608762952
transform 1 0 16560 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_174
timestamp 1608762952
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_178
timestamp 1608762952
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1608762952
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_186
timestamp 1608762952
transform 1 0 18216 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 16008 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_164
timestamp 1608762952
transform 1 0 16192 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 15640 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_160
timestamp 1608762952
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608762952
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1608762952
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_146
timestamp 1608762952
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1608762952
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_129
timestamp 1608762952
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1608762952
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_137
timestamp 1608762952
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1608762952
transform 1 0 14076 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 11776 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_106
timestamp 1608762952
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1608762952
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_114
timestamp 1608762952
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_118
timestamp 1608762952
transform 1 0 11960 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_124
timestamp 1608762952
transform 1 0 12512 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608762952
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1608762952
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1608762952
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1608762952
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1608762952
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_101
timestamp 1608762952
transform 1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1608762952
transform 1 0 8464 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1608762952
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1608762952
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_72
timestamp 1608762952
transform 1 0 7728 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_76
timestamp 1608762952
transform 1 0 8096 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_79
timestamp 1608762952
transform 1 0 8372 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1608762952
transform 1 0 6808 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608762952
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_55
timestamp 1608762952
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1608762952
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_47
timestamp 1608762952
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_51
timestamp 1608762952
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_43
timestamp 1608762952
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1608762952
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_36
timestamp 1608762952
transform 1 0 4416 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1608762952
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608762952
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1608762952
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1608762952
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_21
timestamp 1608762952
transform 1 0 3036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1608762952
transform 1 0 2760 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608762952
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608762952
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1608762952
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1608762952
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1608762952
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_15
timestamp 1608762952
transform 1 0 2484 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608762952
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1608762952
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1608762952
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608762952
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_168
timestamp 1608762952
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1608762952
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_176
timestamp 1608762952
transform 1 0 17296 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1608762952
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1608762952
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_164
timestamp 1608762952
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1608762952
transform 1 0 15640 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1608762952
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1608762952
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1608762952
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_146
timestamp 1608762952
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1608762952
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1608762952
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1608762952
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_129
timestamp 1608762952
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp 1608762952
transform 1 0 13340 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_138
timestamp 1608762952
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_142
timestamp 1608762952
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608762952
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 1608762952
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_110
timestamp 1608762952
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_116
timestamp 1608762952
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1608762952
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1608762952
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_90
timestamp 1608762952
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_94
timestamp 1608762952
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_98
timestamp 1608762952
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_102
timestamp 1608762952
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 7912 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608762952
transform 1 0 6900 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_72
timestamp 1608762952
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608762952
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1608762952
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1608762952
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_52
timestamp 1608762952
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_56
timestamp 1608762952
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1608762952
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1608762952
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1608762952
transform 1 0 4232 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608762952
transform 1 0 4692 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1608762952
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_32
timestamp 1608762952
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_37
timestamp 1608762952
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 2208 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608762952
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1608762952
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_8
timestamp 1608762952
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608762952
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608762952
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1608762952
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1608762952
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1608762952
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_198
timestamp 1608762952
transform 1 0 19320 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_174
timestamp 1608762952
transform 1 0 17112 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_186
timestamp 1608762952
transform 1 0 18216 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608762952
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1608762952
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1608762952
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_158
timestamp 1608762952
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_162
timestamp 1608762952
transform 1 0 16008 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1608762952
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1608762952
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1608762952
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_137
timestamp 1608762952
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1608762952
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 1608762952
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1608762952
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1608762952
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1608762952
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1608762952
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_117
timestamp 1608762952
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1608762952
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1608762952
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608762952
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_105
timestamp 1608762952
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1608762952
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_97
timestamp 1608762952
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608762952
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1608762952
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608762952
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1608762952
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1608762952
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_86
timestamp 1608762952
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762952
transform 1 0 7084 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1608762952
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762952
transform 1 0 5060 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_59
timestamp 1608762952
transform 1 0 6532 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608762952
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608762952
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1608762952
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1608762952
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608762952
transform 1 0 1472 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608762952
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 2024 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608762952
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1608762952
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1608762952
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_8
timestamp 1608762952
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_16
timestamp 1608762952
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608762952
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_209
timestamp 1608762952
transform 1 0 20332 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_217
timestamp 1608762952
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608762952
transform 1 0 18492 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1608762952
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_188
timestamp 1608762952
transform 1 0 18400 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1608762952
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_197
timestamp 1608762952
transform 1 0 19228 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608762952
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_172
timestamp 1608762952
transform 1 0 16928 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1608762952
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1608762952
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_148
timestamp 1608762952
transform 1 0 14720 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_160
timestamp 1608762952
transform 1 0 15824 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_144
timestamp 1608762952
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_140
timestamp 1608762952
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1608762952
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1608762952
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1608762952
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_128
timestamp 1608762952
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608762952
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1608762952
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_108
timestamp 1608762952
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_112
timestamp 1608762952
transform 1 0 11408 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1608762952
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_123
timestamp 1608762952
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608762952
transform 1 0 9476 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_89
timestamp 1608762952
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_100
timestamp 1608762952
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_104
timestamp 1608762952
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608762952
transform 1 0 8464 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1608762952
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608762952
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608762952
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_55
timestamp 1608762952
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608762952
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762952
transform 1 0 3036 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762952
transform 1 0 4692 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1608762952
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762952
transform 1 0 1840 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608762952
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1608762952
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1608762952
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1608762952
transform 1 0 2392 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_18
timestamp 1608762952
transform 1 0 2760 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608762952
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608762952
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1608762952
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1608762952
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1608762952
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608762952
transform 1 0 19044 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608762952
transform 1 0 19596 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_190
timestamp 1608762952
transform 1 0 18584 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_194
timestamp 1608762952
transform 1 0 18952 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_199
timestamp 1608762952
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_205
timestamp 1608762952
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1608762952
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608762952
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1608762952
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1608762952
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1608762952
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1608762952
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_132
timestamp 1608762952
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_136
timestamp 1608762952
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_140
timestamp 1608762952
transform 1 0 13984 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1608762952
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_121
timestamp 1608762952
transform 1 0 12236 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_117
timestamp 1608762952
transform 1 0 11868 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 11316 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_113
timestamp 1608762952
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1608762952
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1608762952
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_101
timestamp 1608762952
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1608762952
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608762952
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1608762952
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1608762952
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1608762952
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_87
timestamp 1608762952
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608762952
transform 1 0 8280 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608762952
transform 1 0 7268 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1608762952
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_76
timestamp 1608762952
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608762952
transform 1 0 6808 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608762952
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1608762952
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608762952
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608762952
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_44
timestamp 1608762952
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_48
timestamp 1608762952
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_52
timestamp 1608762952
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_56
timestamp 1608762952
transform 1 0 6256 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608762952
transform 1 0 4324 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608762952
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1608762952
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608762952
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_21
timestamp 1608762952
transform 1 0 3036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1608762952
transform 1 0 3496 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1608762952
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp 1608762952
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608762952
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1608762952
transform 1 0 2484 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1608762952
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1608762952
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1608762952
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1608762952
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_11
timestamp 1608762952
transform 1 0 2116 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_17
timestamp 1608762952
transform 1 0 2668 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608762952
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608762952
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608762952
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1608762952
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1608762952
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1608762952
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1608762952
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_212
timestamp 1608762952
transform 1 0 20608 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1608762952
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608762952
transform 1 0 19872 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608762952
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1608762952
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_202
timestamp 1608762952
transform 1 0 19688 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_203
timestamp 1608762952
transform 1 0 19780 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1608762952
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1608762952
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_192
timestamp 1608762952
transform 1 0 18768 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_197
timestamp 1608762952
transform 1 0 19228 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608762952
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1608762952
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_175
timestamp 1608762952
transform 1 0 17204 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_184
timestamp 1608762952
transform 1 0 18032 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608762952
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp 1608762952
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1608762952
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1608762952
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1608762952
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_163
timestamp 1608762952
transform 1 0 16100 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_126
timestamp 1608762952
transform 1 0 12696 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_138
timestamp 1608762952
transform 1 0 13800 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1608762952
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1608762952
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_114
timestamp 1608762952
transform 1 0 11592 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608762952
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608762952
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_117
timestamp 1608762952
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1608762952
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1608762952
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608762952
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1608762952
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1608762952
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_108
timestamp 1608762952
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_112
timestamp 1608762952
transform 1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608762952
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1608762952
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_101
timestamp 1608762952
transform 1 0 10396 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_100
timestamp 1608762952
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1608762952
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1608762952
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608762952
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1608762952
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1608762952
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1608762952
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_88
timestamp 1608762952
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1608762952
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_84
timestamp 1608762952
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1608762952
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1608762952
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1608762952
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_73
timestamp 1608762952
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_77
timestamp 1608762952
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_81
timestamp 1608762952
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_76
timestamp 1608762952
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_80
timestamp 1608762952
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608762952
transform 1 0 7268 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1608762952
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1608762952
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1608762952
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1608762952
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1608762952
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1608762952
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608762952
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1608762952
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1608762952
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_60
timestamp 1608762952
transform 1 0 6624 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1608762952
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_56
timestamp 1608762952
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_53
timestamp 1608762952
transform 1 0 5980 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_56
timestamp 1608762952
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1608762952
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_50
timestamp 1608762952
transform 1 0 5704 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_49
timestamp 1608762952
transform 1 0 5612 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1608762952
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_42
timestamp 1608762952
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1608762952
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_45
timestamp 1608762952
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_41
timestamp 1608762952
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608762952
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1608762952
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1608762952
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_36
timestamp 1608762952
transform 1 0 4416 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_35
timestamp 1608762952
transform 1 0 4324 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608762952
transform 1 0 3496 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1608762952
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1608762952
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1608762952
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1608762952
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1608762952
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1608762952
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1608762952
transform 1 0 2484 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_19
timestamp 1608762952
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_17
timestamp 1608762952
transform 1 0 2668 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1608762952
transform 1 0 2300 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1608762952
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_13
timestamp 1608762952
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1608762952
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1608762952
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_7
timestamp 1608762952
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_7
timestamp 1608762952
transform 1 0 1748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608762952
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608762952
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1608762952
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1608762952
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608762952
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608762952
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1608762952
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_210
timestamp 1608762952
transform 1 0 20424 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_215
timestamp 1608762952
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1608762952
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1608762952
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1608762952
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608762952
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1608762952
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1608762952
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1608762952
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1608762952
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1608762952
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608762952
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1608762952
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1608762952
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1608762952
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_87
timestamp 1608762952
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_91
timestamp 1608762952
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_103
timestamp 1608762952
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_83
timestamp 1608762952
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_79
timestamp 1608762952
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_75
timestamp 1608762952
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_70
timestamp 1608762952
transform 1 0 7544 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1608762952
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1608762952
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608762952
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1608762952
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_58
timestamp 1608762952
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1608762952
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_mem_left_track_1.prog_clk_A
timestamp 1608762952
transform 1 0 5888 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_50
timestamp 1608762952
transform 1 0 5704 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_46
timestamp 1608762952
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_42
timestamp 1608762952
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_38
timestamp 1608762952
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1608762952
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_34
timestamp 1608762952
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_29
timestamp 1608762952
transform 1 0 3772 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608762952
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_25
timestamp 1608762952
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1608762952
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_21
timestamp 1608762952
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608762952
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1608762952
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1608762952
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1608762952
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1608762952
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_13
timestamp 1608762952
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1608762952
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608762952
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608762952
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1608762952
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1608762952
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1608762952
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1608762952
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1608762952
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608762952
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1608762952
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1608762952
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1608762952
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1608762952
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1608762952
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1608762952
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608762952
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1608762952
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1608762952
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608762952
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1608762952
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1608762952
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_72
timestamp 1608762952
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_76
timestamp 1608762952
transform 1 0 8096 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_60
timestamp 1608762952
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_55
timestamp 1608762952
transform 1 0 6164 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608762952
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_51
timestamp 1608762952
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_47
timestamp 1608762952
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608762952
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_43
timestamp 1608762952
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1608762952
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_39
timestamp 1608762952
transform 1 0 4692 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608762952
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1608762952
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1608762952
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1608762952
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_25
timestamp 1608762952
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608762952
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1608762952
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 2484 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 2852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1608762952
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1608762952
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1608762952
transform 1 0 2300 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_17
timestamp 1608762952
transform 1 0 2668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608762952
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1608762952
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1608762952
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608762952
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1608762952
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1608762952
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1608762952
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1608762952
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1608762952
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608762952
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1608762952
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1608762952
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1608762952
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1608762952
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_66
timestamp 1608762952
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1608762952
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1608762952
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608762952
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1608762952
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1608762952
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608762952
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608762952
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1608762952
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1608762952
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp 1608762952
transform 1 0 3588 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_32
timestamp 1608762952
transform 1 0 4048 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_40
timestamp 1608762952
transform 1 0 4784 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608762952
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608762952
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1608762952
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1608762952
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1608762952
transform 1 0 2116 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_14
timestamp 1608762952
transform 1 0 2392 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_19
timestamp 1608762952
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608762952
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608762952
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1608762952
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1608762952
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1608762952
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1608762952
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1608762952
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608762952
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1608762952
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1608762952
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1608762952
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1608762952
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1608762952
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1608762952
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608762952
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1608762952
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1608762952
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_69
timestamp 1608762952
transform 1 0 7452 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_81
timestamp 1608762952
transform 1 0 8556 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608762952
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_45
timestamp 1608762952
transform 1 0 5244 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_57
timestamp 1608762952
transform 1 0 6348 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608762952
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_21
timestamp 1608762952
transform 1 0 3036 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1608762952
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_32
timestamp 1608762952
transform 1 0 4048 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_40
timestamp 1608762952
transform 1 0 4784 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608762952
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608762952
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608762952
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1608762952
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608762952
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608762952
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608762952
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1608762952
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1608762952
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1608762952
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1608762952
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1608762952
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608762952
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608762952
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1608762952
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1608762952
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1608762952
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1608762952
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1608762952
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608762952
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608762952
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1608762952
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1608762952
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1608762952
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1608762952
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1608762952
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608762952
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608762952
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608762952
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608762952
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608762952
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1608762952
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1608762952
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608762952
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608762952
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608762952
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1608762952
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1608762952
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608762952
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608762952
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1608762952
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608762952
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608762952
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608762952
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608762952
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51
timestamp 1608762952
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1608762952
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608762952
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608762952
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608762952
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608762952
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608762952
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608762952
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608762952
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608762952
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608762952
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608762952
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608762952
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1608762952
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
<< labels >>
rlabel metal3 s 22000 11432 22800 11552 4 ccff_head
port 1 nsew
rlabel metal2 s 11426 0 11482 800 4 ccff_tail
port 2 nsew
rlabel metal3 s 0 4224 800 4344 4 chanx_left_in[0]
port 3 nsew
rlabel metal3 s 0 8984 800 9104 4 chanx_left_in[10]
port 4 nsew
rlabel metal3 s 0 9392 800 9512 4 chanx_left_in[11]
port 5 nsew
rlabel metal3 s 0 9936 800 10056 4 chanx_left_in[12]
port 6 nsew
rlabel metal3 s 0 10344 800 10464 4 chanx_left_in[13]
port 7 nsew
rlabel metal3 s 0 10752 800 10872 4 chanx_left_in[14]
port 8 nsew
rlabel metal3 s 0 11296 800 11416 4 chanx_left_in[15]
port 9 nsew
rlabel metal3 s 0 11704 800 11824 4 chanx_left_in[16]
port 10 nsew
rlabel metal3 s 0 12248 800 12368 4 chanx_left_in[17]
port 11 nsew
rlabel metal3 s 0 12656 800 12776 4 chanx_left_in[18]
port 12 nsew
rlabel metal3 s 0 13200 800 13320 4 chanx_left_in[19]
port 13 nsew
rlabel metal3 s 0 4768 800 4888 4 chanx_left_in[1]
port 14 nsew
rlabel metal3 s 0 5176 800 5296 4 chanx_left_in[2]
port 15 nsew
rlabel metal3 s 0 5720 800 5840 4 chanx_left_in[3]
port 16 nsew
rlabel metal3 s 0 6128 800 6248 4 chanx_left_in[4]
port 17 nsew
rlabel metal3 s 0 6672 800 6792 4 chanx_left_in[5]
port 18 nsew
rlabel metal3 s 0 7080 800 7200 4 chanx_left_in[6]
port 19 nsew
rlabel metal3 s 0 7488 800 7608 4 chanx_left_in[7]
port 20 nsew
rlabel metal3 s 0 8032 800 8152 4 chanx_left_in[8]
port 21 nsew
rlabel metal3 s 0 8440 800 8560 4 chanx_left_in[9]
port 22 nsew
rlabel metal3 s 0 13608 800 13728 4 chanx_left_out[0]
port 23 nsew
rlabel metal3 s 0 18232 800 18352 4 chanx_left_out[10]
port 24 nsew
rlabel metal3 s 0 18776 800 18896 4 chanx_left_out[11]
port 25 nsew
rlabel metal3 s 0 19184 800 19304 4 chanx_left_out[12]
port 26 nsew
rlabel metal3 s 0 19728 800 19848 4 chanx_left_out[13]
port 27 nsew
rlabel metal3 s 0 20136 800 20256 4 chanx_left_out[14]
port 28 nsew
rlabel metal3 s 0 20544 800 20664 4 chanx_left_out[15]
port 29 nsew
rlabel metal3 s 0 21088 800 21208 4 chanx_left_out[16]
port 30 nsew
rlabel metal3 s 0 21496 800 21616 4 chanx_left_out[17]
port 31 nsew
rlabel metal3 s 0 22040 800 22160 4 chanx_left_out[18]
port 32 nsew
rlabel metal3 s 0 22448 800 22568 4 chanx_left_out[19]
port 33 nsew
rlabel metal3 s 0 14016 800 14136 4 chanx_left_out[1]
port 34 nsew
rlabel metal3 s 0 14560 800 14680 4 chanx_left_out[2]
port 35 nsew
rlabel metal3 s 0 14968 800 15088 4 chanx_left_out[3]
port 36 nsew
rlabel metal3 s 0 15512 800 15632 4 chanx_left_out[4]
port 37 nsew
rlabel metal3 s 0 15920 800 16040 4 chanx_left_out[5]
port 38 nsew
rlabel metal3 s 0 16464 800 16584 4 chanx_left_out[6]
port 39 nsew
rlabel metal3 s 0 16872 800 16992 4 chanx_left_out[7]
port 40 nsew
rlabel metal3 s 0 17280 800 17400 4 chanx_left_out[8]
port 41 nsew
rlabel metal3 s 0 17824 800 17944 4 chanx_left_out[9]
port 42 nsew
rlabel metal2 s 3790 22000 3846 22800 4 chany_top_in[0]
port 43 nsew
rlabel metal2 s 8390 22000 8446 22800 4 chany_top_in[10]
port 44 nsew
rlabel metal2 s 8850 22000 8906 22800 4 chany_top_in[11]
port 45 nsew
rlabel metal2 s 9310 22000 9366 22800 4 chany_top_in[12]
port 46 nsew
rlabel metal2 s 9770 22000 9826 22800 4 chany_top_in[13]
port 47 nsew
rlabel metal2 s 10230 22000 10286 22800 4 chany_top_in[14]
port 48 nsew
rlabel metal2 s 10690 22000 10746 22800 4 chany_top_in[15]
port 49 nsew
rlabel metal2 s 11150 22000 11206 22800 4 chany_top_in[16]
port 50 nsew
rlabel metal2 s 11610 22000 11666 22800 4 chany_top_in[17]
port 51 nsew
rlabel metal2 s 11978 22000 12034 22800 4 chany_top_in[18]
port 52 nsew
rlabel metal2 s 12438 22000 12494 22800 4 chany_top_in[19]
port 53 nsew
rlabel metal2 s 4250 22000 4306 22800 4 chany_top_in[1]
port 54 nsew
rlabel metal2 s 4710 22000 4766 22800 4 chany_top_in[2]
port 55 nsew
rlabel metal2 s 5170 22000 5226 22800 4 chany_top_in[3]
port 56 nsew
rlabel metal2 s 5630 22000 5686 22800 4 chany_top_in[4]
port 57 nsew
rlabel metal2 s 6090 22000 6146 22800 4 chany_top_in[5]
port 58 nsew
rlabel metal2 s 6550 22000 6606 22800 4 chany_top_in[6]
port 59 nsew
rlabel metal2 s 7010 22000 7066 22800 4 chany_top_in[7]
port 60 nsew
rlabel metal2 s 7470 22000 7526 22800 4 chany_top_in[8]
port 61 nsew
rlabel metal2 s 7930 22000 7986 22800 4 chany_top_in[9]
port 62 nsew
rlabel metal2 s 12898 22000 12954 22800 4 chany_top_out[0]
port 63 nsew
rlabel metal2 s 17498 22000 17554 22800 4 chany_top_out[10]
port 64 nsew
rlabel metal2 s 17958 22000 18014 22800 4 chany_top_out[11]
port 65 nsew
rlabel metal2 s 18418 22000 18474 22800 4 chany_top_out[12]
port 66 nsew
rlabel metal2 s 18878 22000 18934 22800 4 chany_top_out[13]
port 67 nsew
rlabel metal2 s 19338 22000 19394 22800 4 chany_top_out[14]
port 68 nsew
rlabel metal2 s 19798 22000 19854 22800 4 chany_top_out[15]
port 69 nsew
rlabel metal2 s 20258 22000 20314 22800 4 chany_top_out[16]
port 70 nsew
rlabel metal2 s 20718 22000 20774 22800 4 chany_top_out[17]
port 71 nsew
rlabel metal2 s 21178 22000 21234 22800 4 chany_top_out[18]
port 72 nsew
rlabel metal2 s 21638 22000 21694 22800 4 chany_top_out[19]
port 73 nsew
rlabel metal2 s 13358 22000 13414 22800 4 chany_top_out[1]
port 74 nsew
rlabel metal2 s 13818 22000 13874 22800 4 chany_top_out[2]
port 75 nsew
rlabel metal2 s 14278 22000 14334 22800 4 chany_top_out[3]
port 76 nsew
rlabel metal2 s 14738 22000 14794 22800 4 chany_top_out[4]
port 77 nsew
rlabel metal2 s 15198 22000 15254 22800 4 chany_top_out[5]
port 78 nsew
rlabel metal2 s 15658 22000 15714 22800 4 chany_top_out[6]
port 79 nsew
rlabel metal2 s 16118 22000 16174 22800 4 chany_top_out[7]
port 80 nsew
rlabel metal2 s 16578 22000 16634 22800 4 chany_top_out[8]
port 81 nsew
rlabel metal2 s 17038 22000 17094 22800 4 chany_top_out[9]
port 82 nsew
rlabel metal3 s 0 2456 800 2576 4 left_bottom_grid_pin_11_
port 83 nsew
rlabel metal3 s 0 2864 800 2984 4 left_bottom_grid_pin_13_
port 84 nsew
rlabel metal3 s 0 3408 800 3528 4 left_bottom_grid_pin_15_
port 85 nsew
rlabel metal3 s 0 3816 800 3936 4 left_bottom_grid_pin_17_
port 86 nsew
rlabel metal3 s 0 144 800 264 4 left_bottom_grid_pin_1_
port 87 nsew
rlabel metal3 s 0 552 800 672 4 left_bottom_grid_pin_3_
port 88 nsew
rlabel metal3 s 0 960 800 1080 4 left_bottom_grid_pin_5_
port 89 nsew
rlabel metal3 s 0 1504 800 1624 4 left_bottom_grid_pin_7_
port 90 nsew
rlabel metal3 s 0 1912 800 2032 4 left_bottom_grid_pin_9_
port 91 nsew
rlabel metal2 s 22098 22000 22154 22800 4 prog_clk_0_N_in
port 92 nsew
rlabel metal2 s 202 22000 258 22800 4 top_left_grid_pin_42_
port 93 nsew
rlabel metal2 s 570 22000 626 22800 4 top_left_grid_pin_43_
port 94 nsew
rlabel metal2 s 1030 22000 1086 22800 4 top_left_grid_pin_44_
port 95 nsew
rlabel metal2 s 1490 22000 1546 22800 4 top_left_grid_pin_45_
port 96 nsew
rlabel metal2 s 1950 22000 2006 22800 4 top_left_grid_pin_46_
port 97 nsew
rlabel metal2 s 2410 22000 2466 22800 4 top_left_grid_pin_47_
port 98 nsew
rlabel metal2 s 2870 22000 2926 22800 4 top_left_grid_pin_48_
port 99 nsew
rlabel metal2 s 3330 22000 3386 22800 4 top_left_grid_pin_49_
port 100 nsew
rlabel metal2 s 22558 22000 22614 22800 4 top_right_grid_pin_1_
port 101 nsew
rlabel metal4 s 4376 2128 4696 20176 4 VPWR
port 102 nsew
rlabel metal4 s 7808 2128 8128 20176 4 VGND
port 103 nsew
<< properties >>
string FIXED_BBOX 0 0 22800 22800
string GDS_FILE /ef/openfpga/openlane/runs/sb_2__0_/results/magic/sb_2__0_.gds
string GDS_END 1340612
string GDS_START 81916
<< end >>
