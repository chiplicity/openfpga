VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__2_
  CLASS BLOCK ;
  FOREIGN cbx_1__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 85.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 82.600 5.890 85.000 ;
    END
  END IO_ISOL_N
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 2.400 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 82.600 16.930 85.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 2.400 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 82.600 27.970 85.000 ;
    END
  END SC_OUT_TOP
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.400 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.400 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 2.400 ;
    END
  END bottom_grid_pin_11_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 2.400 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 2.400 ;
    END
  END bottom_grid_pin_13_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 2.400 ;
    END
  END bottom_grid_pin_15_
  PIN bottom_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 2.400 ;
    END
  END bottom_grid_pin_1_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 2.400 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.400 ;
    END
  END bottom_grid_pin_3_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 2.400 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END bottom_grid_pin_5_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 2.400 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 2.400 ;
    END
  END bottom_grid_pin_7_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 2.400 ;
    END
  END bottom_grid_pin_8_
  PIN bottom_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END bottom_grid_pin_9_
  PIN bottom_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END bottom_width_0_height_0__pin_0_
  PIN bottom_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 2.400 ;
    END
  END bottom_width_0_height_0__pin_1_lower
  PIN bottom_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 2.400 ;
    END
  END bottom_width_0_height_0__pin_1_upper
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 82.600 39.010 85.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 82.600 50.050 85.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 2.400 44.840 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 2.400 65.240 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 2.400 67.280 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 2.400 69.320 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.400 71.360 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 2.400 75.440 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.400 81.560 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 2.400 46.880 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.400 50.960 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 2.400 53.000 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 2.400 55.040 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 2.400 61.160 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 2.400 23.760 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 2.400 27.840 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 2.400 36.000 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 2.400 38.040 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 2.400 40.080 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 2.400 42.120 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 2.400 5.400 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.400 11.520 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 2.400 19.680 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 42.880 100.000 43.480 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 63.960 100.000 64.560 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 66.000 100.000 66.600 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 68.720 100.000 69.320 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 70.760 100.000 71.360 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 72.800 100.000 73.400 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 74.840 100.000 75.440 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 76.880 100.000 77.480 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 78.920 100.000 79.520 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 80.960 100.000 81.560 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 83.000 100.000 83.600 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 44.920 100.000 45.520 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 46.960 100.000 47.560 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 49.000 100.000 49.600 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 51.720 100.000 52.320 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 53.760 100.000 54.360 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 55.800 100.000 56.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 57.840 100.000 58.440 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 59.880 100.000 60.480 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 61.920 100.000 62.520 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 0.720 100.000 1.320 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 21.800 100.000 22.400 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 23.840 100.000 24.440 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 25.880 100.000 26.480 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 27.920 100.000 28.520 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 29.960 100.000 30.560 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 32.000 100.000 32.600 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 34.720 100.000 35.320 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 36.760 100.000 37.360 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 38.800 100.000 39.400 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 40.840 100.000 41.440 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 2.760 100.000 3.360 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 4.800 100.000 5.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 6.840 100.000 7.440 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 8.880 100.000 9.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 10.920 100.000 11.520 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 12.960 100.000 13.560 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 15.000 100.000 15.600 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 17.720 100.000 18.320 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 19.760 100.000 20.360 ;
    END
  END chanx_right_out[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.850 82.600 72.130 85.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 82.600 83.170 85.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 82.600 94.210 85.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END prog_clk_0_S_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END prog_clk_0_W_out
  PIN top_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 82.600 61.090 85.000 ;
    END
  END top_grid_pin_0_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.545 10.640 21.145 73.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.375 10.640 35.975 73.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 73.525 ;
      LAYER met1 ;
        RECT 1.910 4.800 97.450 76.120 ;
      LAYER met2 ;
        RECT 1.940 82.320 5.330 83.485 ;
        RECT 6.170 82.320 16.370 83.485 ;
        RECT 17.210 82.320 27.410 83.485 ;
        RECT 28.250 82.320 38.450 83.485 ;
        RECT 39.290 82.320 49.490 83.485 ;
        RECT 50.330 82.320 60.530 83.485 ;
        RECT 61.370 82.320 71.570 83.485 ;
        RECT 72.410 82.320 82.610 83.485 ;
        RECT 83.450 82.320 93.650 83.485 ;
        RECT 94.490 82.320 97.420 83.485 ;
        RECT 1.940 2.680 97.420 82.320 ;
        RECT 2.490 0.835 5.790 2.680 ;
        RECT 6.630 0.835 10.390 2.680 ;
        RECT 11.230 0.835 14.990 2.680 ;
        RECT 15.830 0.835 19.590 2.680 ;
        RECT 20.430 0.835 24.190 2.680 ;
        RECT 25.030 0.835 28.790 2.680 ;
        RECT 29.630 0.835 33.390 2.680 ;
        RECT 34.230 0.835 37.530 2.680 ;
        RECT 38.370 0.835 42.130 2.680 ;
        RECT 42.970 0.835 46.730 2.680 ;
        RECT 47.570 0.835 51.330 2.680 ;
        RECT 52.170 0.835 55.930 2.680 ;
        RECT 56.770 0.835 60.530 2.680 ;
        RECT 61.370 0.835 65.130 2.680 ;
        RECT 65.970 0.835 69.270 2.680 ;
        RECT 70.110 0.835 73.870 2.680 ;
        RECT 74.710 0.835 78.470 2.680 ;
        RECT 79.310 0.835 83.070 2.680 ;
        RECT 83.910 0.835 87.670 2.680 ;
        RECT 88.510 0.835 92.270 2.680 ;
        RECT 93.110 0.835 96.870 2.680 ;
      LAYER met3 ;
        RECT 2.800 82.600 97.200 83.465 ;
        RECT 2.400 81.960 97.600 82.600 ;
        RECT 2.800 80.560 97.200 81.960 ;
        RECT 2.400 79.920 97.600 80.560 ;
        RECT 2.800 78.520 97.200 79.920 ;
        RECT 2.400 77.880 97.600 78.520 ;
        RECT 2.800 76.480 97.200 77.880 ;
        RECT 2.400 75.840 97.600 76.480 ;
        RECT 2.800 74.440 97.200 75.840 ;
        RECT 2.400 73.800 97.600 74.440 ;
        RECT 2.800 72.400 97.200 73.800 ;
        RECT 2.400 71.760 97.600 72.400 ;
        RECT 2.800 70.360 97.200 71.760 ;
        RECT 2.400 69.720 97.600 70.360 ;
        RECT 2.800 68.320 97.200 69.720 ;
        RECT 2.400 67.680 97.600 68.320 ;
        RECT 2.800 67.000 97.600 67.680 ;
        RECT 2.800 66.280 97.200 67.000 ;
        RECT 2.400 65.640 97.200 66.280 ;
        RECT 2.800 65.600 97.200 65.640 ;
        RECT 2.800 64.960 97.600 65.600 ;
        RECT 2.800 64.240 97.200 64.960 ;
        RECT 2.400 63.600 97.200 64.240 ;
        RECT 2.800 63.560 97.200 63.600 ;
        RECT 2.800 62.920 97.600 63.560 ;
        RECT 2.800 62.200 97.200 62.920 ;
        RECT 2.400 61.560 97.200 62.200 ;
        RECT 2.800 61.520 97.200 61.560 ;
        RECT 2.800 60.880 97.600 61.520 ;
        RECT 2.800 60.160 97.200 60.880 ;
        RECT 2.400 59.520 97.200 60.160 ;
        RECT 2.800 59.480 97.200 59.520 ;
        RECT 2.800 58.840 97.600 59.480 ;
        RECT 2.800 58.120 97.200 58.840 ;
        RECT 2.400 57.480 97.200 58.120 ;
        RECT 2.800 57.440 97.200 57.480 ;
        RECT 2.800 56.800 97.600 57.440 ;
        RECT 2.800 56.080 97.200 56.800 ;
        RECT 2.400 55.440 97.200 56.080 ;
        RECT 2.800 55.400 97.200 55.440 ;
        RECT 2.800 54.760 97.600 55.400 ;
        RECT 2.800 54.040 97.200 54.760 ;
        RECT 2.400 53.400 97.200 54.040 ;
        RECT 2.800 53.360 97.200 53.400 ;
        RECT 2.800 52.720 97.600 53.360 ;
        RECT 2.800 52.000 97.200 52.720 ;
        RECT 2.400 51.360 97.200 52.000 ;
        RECT 2.800 51.320 97.200 51.360 ;
        RECT 2.800 50.000 97.600 51.320 ;
        RECT 2.800 49.960 97.200 50.000 ;
        RECT 2.400 49.320 97.200 49.960 ;
        RECT 2.800 48.600 97.200 49.320 ;
        RECT 2.800 47.960 97.600 48.600 ;
        RECT 2.800 47.920 97.200 47.960 ;
        RECT 2.400 47.280 97.200 47.920 ;
        RECT 2.800 46.560 97.200 47.280 ;
        RECT 2.800 45.920 97.600 46.560 ;
        RECT 2.800 45.880 97.200 45.920 ;
        RECT 2.400 45.240 97.200 45.880 ;
        RECT 2.800 44.520 97.200 45.240 ;
        RECT 2.800 43.880 97.600 44.520 ;
        RECT 2.800 43.840 97.200 43.880 ;
        RECT 2.400 42.520 97.200 43.840 ;
        RECT 2.800 42.480 97.200 42.520 ;
        RECT 2.800 41.840 97.600 42.480 ;
        RECT 2.800 41.120 97.200 41.840 ;
        RECT 2.400 40.480 97.200 41.120 ;
        RECT 2.800 40.440 97.200 40.480 ;
        RECT 2.800 39.800 97.600 40.440 ;
        RECT 2.800 39.080 97.200 39.800 ;
        RECT 2.400 38.440 97.200 39.080 ;
        RECT 2.800 38.400 97.200 38.440 ;
        RECT 2.800 37.760 97.600 38.400 ;
        RECT 2.800 37.040 97.200 37.760 ;
        RECT 2.400 36.400 97.200 37.040 ;
        RECT 2.800 36.360 97.200 36.400 ;
        RECT 2.800 35.720 97.600 36.360 ;
        RECT 2.800 35.000 97.200 35.720 ;
        RECT 2.400 34.360 97.200 35.000 ;
        RECT 2.800 34.320 97.200 34.360 ;
        RECT 2.800 33.000 97.600 34.320 ;
        RECT 2.800 32.960 97.200 33.000 ;
        RECT 2.400 32.320 97.200 32.960 ;
        RECT 2.800 31.600 97.200 32.320 ;
        RECT 2.800 30.960 97.600 31.600 ;
        RECT 2.800 30.920 97.200 30.960 ;
        RECT 2.400 30.280 97.200 30.920 ;
        RECT 2.800 29.560 97.200 30.280 ;
        RECT 2.800 28.920 97.600 29.560 ;
        RECT 2.800 28.880 97.200 28.920 ;
        RECT 2.400 28.240 97.200 28.880 ;
        RECT 2.800 27.520 97.200 28.240 ;
        RECT 2.800 26.880 97.600 27.520 ;
        RECT 2.800 26.840 97.200 26.880 ;
        RECT 2.400 26.200 97.200 26.840 ;
        RECT 2.800 25.480 97.200 26.200 ;
        RECT 2.800 24.840 97.600 25.480 ;
        RECT 2.800 24.800 97.200 24.840 ;
        RECT 2.400 24.160 97.200 24.800 ;
        RECT 2.800 23.440 97.200 24.160 ;
        RECT 2.800 22.800 97.600 23.440 ;
        RECT 2.800 22.760 97.200 22.800 ;
        RECT 2.400 22.120 97.200 22.760 ;
        RECT 2.800 21.400 97.200 22.120 ;
        RECT 2.800 20.760 97.600 21.400 ;
        RECT 2.800 20.720 97.200 20.760 ;
        RECT 2.400 20.080 97.200 20.720 ;
        RECT 2.800 19.360 97.200 20.080 ;
        RECT 2.800 18.720 97.600 19.360 ;
        RECT 2.800 18.680 97.200 18.720 ;
        RECT 2.400 18.040 97.200 18.680 ;
        RECT 2.800 17.320 97.200 18.040 ;
        RECT 2.800 16.640 97.600 17.320 ;
        RECT 2.400 16.000 97.600 16.640 ;
        RECT 2.800 14.600 97.200 16.000 ;
        RECT 2.400 13.960 97.600 14.600 ;
        RECT 2.800 12.560 97.200 13.960 ;
        RECT 2.400 11.920 97.600 12.560 ;
        RECT 2.800 10.520 97.200 11.920 ;
        RECT 2.400 9.880 97.600 10.520 ;
        RECT 2.800 8.480 97.200 9.880 ;
        RECT 2.400 7.840 97.600 8.480 ;
        RECT 2.800 6.440 97.200 7.840 ;
        RECT 2.400 5.800 97.600 6.440 ;
        RECT 2.800 4.400 97.200 5.800 ;
        RECT 2.400 3.760 97.600 4.400 ;
        RECT 2.800 2.360 97.200 3.760 ;
        RECT 2.400 1.720 97.600 2.360 ;
        RECT 2.800 0.855 97.200 1.720 ;
      LAYER met4 ;
        RECT 21.455 74.080 80.450 81.425 ;
        RECT 21.545 10.640 33.975 74.080 ;
        RECT 36.375 10.640 80.450 74.080 ;
  END
END cbx_1__2_
END LIBRARY

