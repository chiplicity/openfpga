magic
tech sky130A
magscale 1 2
timestamp 1606475969
<< locali >>
rect 5917 8891 5951 9129
rect 14105 6171 14139 6341
rect 12081 5627 12115 5729
rect 6561 5015 6595 5253
rect 10333 5151 10367 5253
rect 9413 4675 9447 4709
rect 9413 4641 9597 4675
rect 8585 4063 8619 4165
rect 9597 3995 9631 4165
rect 10701 3383 10735 3485
rect 13369 2907 13403 3077
<< viali >>
rect 1961 20009 1995 20043
rect 1777 19873 1811 19907
rect 7021 19465 7055 19499
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 6837 19261 6871 19295
rect 1961 19125 1995 19159
rect 2513 19125 2547 19159
rect 7481 18921 7515 18955
rect 3157 18853 3191 18887
rect 2145 18785 2179 18819
rect 2881 18785 2915 18819
rect 7297 18785 7331 18819
rect 2329 18717 2363 18751
rect 2513 18377 2547 18411
rect 3065 18377 3099 18411
rect 7205 18241 7239 18275
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 2881 18173 2915 18207
rect 7021 18173 7055 18207
rect 1961 18037 1995 18071
rect 1869 17833 1903 17867
rect 3157 17833 3191 17867
rect 2513 17765 2547 17799
rect 8033 17765 8067 17799
rect 10333 17765 10367 17799
rect 1685 17697 1719 17731
rect 2237 17697 2271 17731
rect 2973 17697 3007 17731
rect 7757 17697 7791 17731
rect 10057 17697 10091 17731
rect 1777 17289 1811 17323
rect 10701 17289 10735 17323
rect 5549 17221 5583 17255
rect 9137 17221 9171 17255
rect 2329 17153 2363 17187
rect 6193 17153 6227 17187
rect 8585 17153 8619 17187
rect 9781 17153 9815 17187
rect 11345 17153 11379 17187
rect 1593 17085 1627 17119
rect 2145 17085 2179 17119
rect 2881 17085 2915 17119
rect 8401 17085 8435 17119
rect 3157 17017 3191 17051
rect 11069 17017 11103 17051
rect 11713 17017 11747 17051
rect 3985 16949 4019 16983
rect 5917 16949 5951 16983
rect 6009 16949 6043 16983
rect 9505 16949 9539 16983
rect 9597 16949 9631 16983
rect 11161 16949 11195 16983
rect 3341 16745 3375 16779
rect 5733 16745 5767 16779
rect 7389 16745 7423 16779
rect 9137 16745 9171 16779
rect 11069 16745 11103 16779
rect 12725 16745 12759 16779
rect 1961 16677 1995 16711
rect 2697 16677 2731 16711
rect 1685 16609 1719 16643
rect 2421 16609 2455 16643
rect 3157 16609 3191 16643
rect 4353 16609 4387 16643
rect 4620 16609 4654 16643
rect 6276 16609 6310 16643
rect 9689 16609 9723 16643
rect 9956 16609 9990 16643
rect 11345 16609 11379 16643
rect 11612 16609 11646 16643
rect 6009 16541 6043 16575
rect 7941 16541 7975 16575
rect 2973 16201 3007 16235
rect 4905 16201 4939 16235
rect 5181 16201 5215 16235
rect 7205 16201 7239 16235
rect 11529 16201 11563 16235
rect 2329 16065 2363 16099
rect 3525 16065 3559 16099
rect 5733 16065 5767 16099
rect 6193 16065 6227 16099
rect 7849 16065 7883 16099
rect 10149 16065 10183 16099
rect 1501 15997 1535 16031
rect 2053 15997 2087 16031
rect 2789 15997 2823 16031
rect 5549 15997 5583 16031
rect 7573 15997 7607 16031
rect 8224 15997 8258 16031
rect 10416 15997 10450 16031
rect 3792 15929 3826 15963
rect 8484 15929 8518 15963
rect 1685 15861 1719 15895
rect 5641 15861 5675 15895
rect 7665 15861 7699 15895
rect 9597 15861 9631 15895
rect 1685 15657 1719 15691
rect 2789 15657 2823 15691
rect 4261 15657 4295 15691
rect 8953 15657 8987 15691
rect 9689 15657 9723 15691
rect 10977 15657 11011 15691
rect 2329 15589 2363 15623
rect 6184 15589 6218 15623
rect 10149 15589 10183 15623
rect 10609 15589 10643 15623
rect 1501 15521 1535 15555
rect 2053 15521 2087 15555
rect 3157 15521 3191 15555
rect 3249 15521 3283 15555
rect 4629 15521 4663 15555
rect 4721 15521 4755 15555
rect 5917 15521 5951 15555
rect 7840 15521 7874 15555
rect 10057 15521 10091 15555
rect 11345 15521 11379 15555
rect 3341 15453 3375 15487
rect 4813 15453 4847 15487
rect 7573 15453 7607 15487
rect 10241 15453 10275 15487
rect 11437 15453 11471 15487
rect 11621 15453 11655 15487
rect 5181 15317 5215 15351
rect 7297 15317 7331 15351
rect 11805 15317 11839 15351
rect 4169 15113 4203 15147
rect 4629 15113 4663 15147
rect 5733 15113 5767 15147
rect 8033 15113 8067 15147
rect 10609 15113 10643 15147
rect 1685 15045 1719 15079
rect 7021 15045 7055 15079
rect 2237 14977 2271 15011
rect 2789 14977 2823 15011
rect 5181 14977 5215 15011
rect 6285 14977 6319 15011
rect 7573 14977 7607 15011
rect 8677 14977 8711 15011
rect 1501 14909 1535 14943
rect 2053 14909 2087 14943
rect 3056 14909 3090 14943
rect 4997 14909 5031 14943
rect 6193 14909 6227 14943
rect 9229 14909 9263 14943
rect 7481 14841 7515 14875
rect 7849 14841 7883 14875
rect 9474 14841 9508 14875
rect 4537 14773 4571 14807
rect 5089 14773 5123 14807
rect 6101 14773 6135 14807
rect 7389 14773 7423 14807
rect 8401 14773 8435 14807
rect 8493 14773 8527 14807
rect 8953 14773 8987 14807
rect 1685 14569 1719 14603
rect 3433 14569 3467 14603
rect 4445 14569 4479 14603
rect 2320 14501 2354 14535
rect 4813 14501 4847 14535
rect 6644 14501 6678 14535
rect 9045 14501 9079 14535
rect 1501 14433 1535 14467
rect 2053 14433 2087 14467
rect 4905 14433 4939 14467
rect 8953 14433 8987 14467
rect 9956 14433 9990 14467
rect 4997 14365 5031 14399
rect 5917 14365 5951 14399
rect 6377 14365 6411 14399
rect 9229 14365 9263 14399
rect 9689 14365 9723 14399
rect 7757 14297 7791 14331
rect 8585 14229 8619 14263
rect 11069 14229 11103 14263
rect 3433 14025 3467 14059
rect 5641 14025 5675 14059
rect 9965 14025 9999 14059
rect 2053 13889 2087 13923
rect 4261 13889 4295 13923
rect 1777 13821 1811 13855
rect 2513 13821 2547 13855
rect 2789 13821 2823 13855
rect 3249 13821 3283 13855
rect 6837 13821 6871 13855
rect 7104 13821 7138 13855
rect 8585 13821 8619 13855
rect 3801 13753 3835 13787
rect 4528 13753 4562 13787
rect 5917 13753 5951 13787
rect 8852 13753 8886 13787
rect 10241 13753 10275 13787
rect 8217 13685 8251 13719
rect 3525 13481 3559 13515
rect 5457 13481 5491 13515
rect 5733 13481 5767 13515
rect 6101 13481 6135 13515
rect 8953 13481 8987 13515
rect 9689 13481 9723 13515
rect 2145 13413 2179 13447
rect 4344 13413 4378 13447
rect 9045 13413 9079 13447
rect 10057 13413 10091 13447
rect 1869 13345 1903 13379
rect 2605 13345 2639 13379
rect 3341 13345 3375 13379
rect 4077 13345 4111 13379
rect 7297 13345 7331 13379
rect 7941 13345 7975 13379
rect 8033 13345 8067 13379
rect 10149 13345 10183 13379
rect 2789 13277 2823 13311
rect 6193 13277 6227 13311
rect 6285 13277 6319 13311
rect 8217 13277 8251 13311
rect 9137 13277 9171 13311
rect 10241 13277 10275 13311
rect 7573 13209 7607 13243
rect 8585 13209 8619 13243
rect 7113 13141 7147 13175
rect 6009 12937 6043 12971
rect 9045 12937 9079 12971
rect 10057 12937 10091 12971
rect 2053 12801 2087 12835
rect 7205 12801 7239 12835
rect 7665 12801 7699 12835
rect 1777 12733 1811 12767
rect 2881 12733 2915 12767
rect 4629 12733 4663 12767
rect 10241 12733 10275 12767
rect 3126 12665 3160 12699
rect 4896 12665 4930 12699
rect 7932 12665 7966 12699
rect 4261 12597 4295 12631
rect 6285 12597 6319 12631
rect 1685 12393 1719 12427
rect 2053 12393 2087 12427
rect 4537 12393 4571 12427
rect 4905 12393 4939 12427
rect 9689 12393 9723 12427
rect 10057 12325 10091 12359
rect 1501 12257 1535 12291
rect 2421 12257 2455 12291
rect 4445 12257 4479 12291
rect 5549 12257 5583 12291
rect 5816 12257 5850 12291
rect 7564 12257 7598 12291
rect 19533 12257 19567 12291
rect 2513 12189 2547 12223
rect 2697 12189 2731 12223
rect 3065 12189 3099 12223
rect 4997 12189 5031 12223
rect 5181 12189 5215 12223
rect 7297 12189 7331 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 4261 12121 4295 12155
rect 8677 12121 8711 12155
rect 6929 12053 6963 12087
rect 19717 12053 19751 12087
rect 3433 11849 3467 11883
rect 3709 11849 3743 11883
rect 6469 11849 6503 11883
rect 7665 11849 7699 11883
rect 10701 11849 10735 11883
rect 7021 11781 7055 11815
rect 4261 11713 4295 11747
rect 8217 11713 8251 11747
rect 9321 11713 9355 11747
rect 2053 11645 2087 11679
rect 2320 11645 2354 11679
rect 4077 11645 4111 11679
rect 5089 11645 5123 11679
rect 7205 11645 7239 11679
rect 19073 11645 19107 11679
rect 5356 11577 5390 11611
rect 8033 11577 8067 11611
rect 8677 11577 8711 11611
rect 9588 11577 9622 11611
rect 4169 11509 4203 11543
rect 8125 11509 8159 11543
rect 19257 11509 19291 11543
rect 1409 11305 1443 11339
rect 1777 11305 1811 11339
rect 2421 11305 2455 11339
rect 4445 11305 4479 11339
rect 5457 11305 5491 11339
rect 6929 11305 6963 11339
rect 8585 11305 8619 11339
rect 11069 11305 11103 11339
rect 4813 11237 4847 11271
rect 6469 11237 6503 11271
rect 2789 11169 2823 11203
rect 4905 11169 4939 11203
rect 5825 11169 5859 11203
rect 7297 11169 7331 11203
rect 7389 11169 7423 11203
rect 8953 11169 8987 11203
rect 9689 11169 9723 11203
rect 9956 11169 9990 11203
rect 18619 11169 18653 11203
rect 1869 11101 1903 11135
rect 2053 11101 2087 11135
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 5089 11101 5123 11135
rect 5917 11101 5951 11135
rect 6101 11101 6135 11135
rect 7573 11101 7607 11135
rect 9045 11101 9079 11135
rect 9229 11101 9263 11135
rect 18797 11033 18831 11067
rect 2973 10761 3007 10795
rect 3709 10761 3743 10795
rect 6469 10761 6503 10795
rect 9413 10761 9447 10795
rect 9137 10693 9171 10727
rect 1593 10625 1627 10659
rect 4353 10625 4387 10659
rect 5089 10625 5123 10659
rect 10057 10625 10091 10659
rect 1860 10557 1894 10591
rect 7389 10557 7423 10591
rect 7757 10557 7791 10591
rect 8013 10557 8047 10591
rect 11069 10557 11103 10591
rect 18245 10557 18279 10591
rect 4077 10489 4111 10523
rect 5356 10489 5390 10523
rect 9781 10489 9815 10523
rect 10425 10489 10459 10523
rect 4169 10421 4203 10455
rect 7205 10421 7239 10455
rect 9873 10421 9907 10455
rect 10885 10421 10919 10455
rect 18429 10421 18463 10455
rect 2789 10217 2823 10251
rect 5733 10217 5767 10251
rect 8217 10217 8251 10251
rect 8585 10217 8619 10251
rect 11345 10217 11379 10251
rect 3157 10149 3191 10183
rect 3249 10081 3283 10115
rect 4620 10081 4654 10115
rect 6837 10081 6871 10115
rect 7104 10081 7138 10115
rect 8953 10081 8987 10115
rect 9873 10081 9907 10115
rect 3341 10013 3375 10047
rect 4353 10013 4387 10047
rect 9045 10013 9079 10047
rect 9229 10013 9263 10047
rect 2973 9673 3007 9707
rect 4905 9673 4939 9707
rect 11069 9673 11103 9707
rect 5181 9605 5215 9639
rect 7849 9605 7883 9639
rect 8861 9605 8895 9639
rect 5733 9537 5767 9571
rect 7389 9537 7423 9571
rect 8401 9537 8435 9571
rect 9413 9537 9447 9571
rect 1593 9469 1627 9503
rect 3525 9469 3559 9503
rect 3792 9469 3826 9503
rect 5641 9469 5675 9503
rect 7205 9469 7239 9503
rect 9229 9469 9263 9503
rect 9689 9469 9723 9503
rect 9945 9469 9979 9503
rect 1860 9401 1894 9435
rect 6285 9401 6319 9435
rect 8217 9401 8251 9435
rect 9321 9401 9355 9435
rect 5549 9333 5583 9367
rect 6837 9333 6871 9367
rect 7297 9333 7331 9367
rect 8309 9333 8343 9367
rect 2789 9129 2823 9163
rect 4445 9129 4479 9163
rect 5917 9129 5951 9163
rect 6101 9129 6135 9163
rect 8493 9129 8527 9163
rect 3525 9061 3559 9095
rect 1676 8993 1710 9027
rect 4537 8993 4571 9027
rect 5457 8993 5491 9027
rect 1409 8925 1443 8959
rect 3065 8925 3099 8959
rect 4721 8925 4755 8959
rect 5549 8925 5583 8959
rect 5641 8925 5675 8959
rect 6469 9061 6503 9095
rect 7113 8993 7147 9027
rect 8585 8993 8619 9027
rect 10140 8993 10174 9027
rect 6561 8925 6595 8959
rect 6653 8925 6687 8959
rect 7297 8925 7331 8959
rect 8769 8925 8803 8959
rect 9873 8925 9907 8959
rect 5917 8857 5951 8891
rect 4077 8789 4111 8823
rect 5089 8789 5123 8823
rect 8125 8789 8159 8823
rect 11253 8789 11287 8823
rect 1777 8585 1811 8619
rect 4445 8585 4479 8619
rect 5733 8585 5767 8619
rect 9229 8585 9263 8619
rect 10977 8585 11011 8619
rect 11253 8585 11287 8619
rect 4169 8517 4203 8551
rect 2237 8449 2271 8483
rect 2421 8449 2455 8483
rect 4905 8449 4939 8483
rect 4997 8449 5031 8483
rect 6377 8449 6411 8483
rect 7297 8449 7331 8483
rect 2789 8381 2823 8415
rect 4813 8381 4847 8415
rect 5641 8381 5675 8415
rect 6193 8381 6227 8415
rect 9413 8381 9447 8415
rect 9597 8381 9631 8415
rect 11437 8381 11471 8415
rect 3056 8313 3090 8347
rect 6837 8313 6871 8347
rect 7564 8313 7598 8347
rect 9864 8313 9898 8347
rect 2145 8245 2179 8279
rect 5457 8245 5491 8279
rect 6101 8245 6135 8279
rect 8677 8245 8711 8279
rect 2237 8041 2271 8075
rect 2697 8041 2731 8075
rect 4077 8041 4111 8075
rect 7941 8041 7975 8075
rect 8309 8041 8343 8075
rect 10609 8041 10643 8075
rect 11161 8041 11195 8075
rect 16681 8041 16715 8075
rect 2605 7973 2639 8007
rect 7389 7973 7423 8007
rect 11621 7973 11655 8007
rect 15568 7973 15602 8007
rect 3893 7905 3927 7939
rect 4445 7905 4479 7939
rect 5448 7905 5482 7939
rect 7297 7905 7331 7939
rect 9689 7905 9723 7939
rect 10517 7905 10551 7939
rect 11529 7905 11563 7939
rect 2789 7837 2823 7871
rect 4537 7837 4571 7871
rect 4721 7837 4755 7871
rect 5181 7837 5215 7871
rect 7573 7837 7607 7871
rect 8401 7837 8435 7871
rect 8493 7837 8527 7871
rect 10793 7837 10827 7871
rect 11713 7837 11747 7871
rect 15301 7837 15335 7871
rect 10149 7769 10183 7803
rect 3709 7701 3743 7735
rect 6561 7701 6595 7735
rect 6929 7701 6963 7735
rect 1961 7497 1995 7531
rect 6837 7497 6871 7531
rect 8125 7497 8159 7531
rect 14289 7429 14323 7463
rect 2513 7361 2547 7395
rect 3617 7361 3651 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 8677 7361 8711 7395
rect 10333 7361 10367 7395
rect 14933 7361 14967 7395
rect 4445 7293 4479 7327
rect 4712 7293 4746 7327
rect 7205 7293 7239 7327
rect 8493 7293 8527 7327
rect 12173 7293 12207 7327
rect 16957 7293 16991 7327
rect 2329 7225 2363 7259
rect 10600 7225 10634 7259
rect 14749 7225 14783 7259
rect 17233 7225 17267 7259
rect 2421 7157 2455 7191
rect 2973 7157 3007 7191
rect 3341 7157 3375 7191
rect 3433 7157 3467 7191
rect 5825 7157 5859 7191
rect 6285 7157 6319 7191
rect 8585 7157 8619 7191
rect 11713 7157 11747 7191
rect 11989 7157 12023 7191
rect 13645 7157 13679 7191
rect 14657 7157 14691 7191
rect 15577 7157 15611 7191
rect 4077 6953 4111 6987
rect 4445 6953 4479 6987
rect 14473 6953 14507 6987
rect 10333 6885 10367 6919
rect 11244 6885 11278 6919
rect 2228 6817 2262 6851
rect 4537 6817 4571 6851
rect 5365 6817 5399 6851
rect 5724 6817 5758 6851
rect 7369 6817 7403 6851
rect 13093 6817 13127 6851
rect 13360 6817 13394 6851
rect 15568 6817 15602 6851
rect 16957 6817 16991 6851
rect 1961 6749 1995 6783
rect 4721 6749 4755 6783
rect 5457 6749 5491 6783
rect 7113 6749 7147 6783
rect 10425 6749 10459 6783
rect 10609 6749 10643 6783
rect 10977 6749 11011 6783
rect 12633 6749 12667 6783
rect 15301 6749 15335 6783
rect 17233 6749 17267 6783
rect 3341 6681 3375 6715
rect 6837 6681 6871 6715
rect 5181 6613 5215 6647
rect 8493 6613 8527 6647
rect 9965 6613 9999 6647
rect 12357 6613 12391 6647
rect 16681 6613 16715 6647
rect 2789 6409 2823 6443
rect 4997 6409 5031 6443
rect 13921 6409 13955 6443
rect 15209 6409 15243 6443
rect 14105 6341 14139 6375
rect 6285 6273 6319 6307
rect 7389 6273 7423 6307
rect 8217 6273 8251 6307
rect 10425 6273 10459 6307
rect 11621 6273 11655 6307
rect 12541 6273 12575 6307
rect 1409 6205 1443 6239
rect 3617 6205 3651 6239
rect 3884 6205 3918 6239
rect 6009 6205 6043 6239
rect 7205 6205 7239 6239
rect 8484 6205 8518 6239
rect 10241 6205 10275 6239
rect 11437 6205 11471 6239
rect 14749 6273 14783 6307
rect 15761 6273 15795 6307
rect 14565 6205 14599 6239
rect 15669 6205 15703 6239
rect 16313 6205 16347 6239
rect 1676 6137 1710 6171
rect 7297 6137 7331 6171
rect 12808 6137 12842 6171
rect 14105 6137 14139 6171
rect 14657 6137 14691 6171
rect 16580 6137 16614 6171
rect 3065 6069 3099 6103
rect 5641 6069 5675 6103
rect 6101 6069 6135 6103
rect 6837 6069 6871 6103
rect 9597 6069 9631 6103
rect 9873 6069 9907 6103
rect 10333 6069 10367 6103
rect 11069 6069 11103 6103
rect 11529 6069 11563 6103
rect 14197 6069 14231 6103
rect 15577 6069 15611 6103
rect 17693 6069 17727 6103
rect 1501 5865 1535 5899
rect 1869 5865 1903 5899
rect 4077 5865 4111 5899
rect 9045 5865 9079 5899
rect 13553 5865 13587 5899
rect 14289 5865 14323 5899
rect 17417 5865 17451 5899
rect 10762 5797 10796 5831
rect 14197 5797 14231 5831
rect 16304 5797 16338 5831
rect 2881 5729 2915 5763
rect 4445 5729 4479 5763
rect 5549 5729 5583 5763
rect 5816 5729 5850 5763
rect 7573 5729 7607 5763
rect 8953 5729 8987 5763
rect 9689 5729 9723 5763
rect 10425 5729 10459 5763
rect 10517 5729 10551 5763
rect 12081 5729 12115 5763
rect 12440 5729 12474 5763
rect 15025 5729 15059 5763
rect 15301 5729 15335 5763
rect 17693 5729 17727 5763
rect 1961 5661 1995 5695
rect 2145 5661 2179 5695
rect 2973 5661 3007 5695
rect 3065 5661 3099 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 7665 5661 7699 5695
rect 7849 5661 7883 5695
rect 9229 5661 9263 5695
rect 12173 5661 12207 5695
rect 14381 5661 14415 5695
rect 15485 5661 15519 5695
rect 16037 5661 16071 5695
rect 8585 5593 8619 5627
rect 10241 5593 10275 5627
rect 11897 5593 11931 5627
rect 12081 5593 12115 5627
rect 2513 5525 2547 5559
rect 6929 5525 6963 5559
rect 7205 5525 7239 5559
rect 13829 5525 13863 5559
rect 14841 5525 14875 5559
rect 17877 5525 17911 5559
rect 5733 5321 5767 5355
rect 8217 5321 8251 5355
rect 6561 5253 6595 5287
rect 10149 5253 10183 5287
rect 10333 5253 10367 5287
rect 10425 5253 10459 5287
rect 2421 5185 2455 5219
rect 3341 5185 3375 5219
rect 4813 5185 4847 5219
rect 6377 5185 6411 5219
rect 4629 5117 4663 5151
rect 2145 5049 2179 5083
rect 10977 5185 11011 5219
rect 13001 5185 13035 5219
rect 15669 5185 15703 5219
rect 15853 5185 15887 5219
rect 16865 5185 16899 5219
rect 6837 5117 6871 5151
rect 8769 5117 8803 5151
rect 9025 5117 9059 5151
rect 10333 5117 10367 5151
rect 12909 5117 12943 5151
rect 13645 5117 13679 5151
rect 14381 5117 14415 5151
rect 15577 5117 15611 5151
rect 17233 5117 17267 5151
rect 7104 5049 7138 5083
rect 10885 5049 10919 5083
rect 11897 5049 11931 5083
rect 12817 5049 12851 5083
rect 13921 5049 13955 5083
rect 14657 5049 14691 5083
rect 16589 5049 16623 5083
rect 1777 4981 1811 5015
rect 2237 4981 2271 5015
rect 2789 4981 2823 5015
rect 3157 4981 3191 5015
rect 3249 4981 3283 5015
rect 4261 4981 4295 5015
rect 4721 4981 4755 5015
rect 6101 4981 6135 5015
rect 6193 4981 6227 5015
rect 6561 4981 6595 5015
rect 10793 4981 10827 5015
rect 12449 4981 12483 5015
rect 15209 4981 15243 5015
rect 16221 4981 16255 5015
rect 16681 4981 16715 5015
rect 1409 4777 1443 4811
rect 4997 4777 5031 4811
rect 5549 4777 5583 4811
rect 6561 4777 6595 4811
rect 14197 4777 14231 4811
rect 8217 4709 8251 4743
rect 9413 4709 9447 4743
rect 9934 4709 9968 4743
rect 18328 4709 18362 4743
rect 2136 4641 2170 4675
rect 4905 4641 4939 4675
rect 5917 4641 5951 4675
rect 6009 4641 6043 4675
rect 6929 4641 6963 4675
rect 9597 4641 9631 4675
rect 12449 4641 12483 4675
rect 14105 4641 14139 4675
rect 15752 4641 15786 4675
rect 17141 4641 17175 4675
rect 18061 4641 18095 4675
rect 1869 4573 1903 4607
rect 5089 4573 5123 4607
rect 6101 4573 6135 4607
rect 7021 4573 7055 4607
rect 7205 4573 7239 4607
rect 8309 4573 8343 4607
rect 8401 4573 8435 4607
rect 9689 4573 9723 4607
rect 11345 4573 11379 4607
rect 12725 4573 12759 4607
rect 14381 4573 14415 4607
rect 15485 4573 15519 4607
rect 17325 4573 17359 4607
rect 13737 4505 13771 4539
rect 3249 4437 3283 4471
rect 4537 4437 4571 4471
rect 7849 4437 7883 4471
rect 11069 4437 11103 4471
rect 16865 4437 16899 4471
rect 19441 4437 19475 4471
rect 6469 4233 6503 4267
rect 14749 4233 14783 4267
rect 16405 4233 16439 4267
rect 16681 4233 16715 4267
rect 8585 4165 8619 4199
rect 2605 4097 2639 4131
rect 6837 4097 6871 4131
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 9597 4165 9631 4199
rect 9413 4097 9447 4131
rect 2329 4029 2363 4063
rect 2973 4029 3007 4063
rect 3240 4029 3274 4063
rect 5089 4029 5123 4063
rect 8585 4029 8619 4063
rect 9229 4029 9263 4063
rect 17233 4097 17267 4131
rect 9781 4029 9815 4063
rect 10048 4029 10082 4063
rect 11437 4029 11471 4063
rect 12633 4029 12667 4063
rect 13369 4029 13403 4063
rect 15025 4029 15059 4063
rect 15281 4029 15315 4063
rect 5356 3961 5390 3995
rect 9597 3961 9631 3995
rect 11713 3961 11747 3995
rect 12909 3961 12943 3995
rect 13636 3961 13670 3995
rect 17049 3961 17083 3995
rect 1961 3893 1995 3927
rect 2421 3893 2455 3927
rect 4353 3893 4387 3927
rect 7757 3893 7791 3927
rect 8125 3893 8159 3927
rect 8769 3893 8803 3927
rect 9137 3893 9171 3927
rect 11161 3893 11195 3927
rect 17141 3893 17175 3927
rect 13921 3689 13955 3723
rect 15853 3689 15887 3723
rect 18337 3689 18371 3723
rect 4077 3621 4111 3655
rect 6837 3621 6871 3655
rect 10333 3621 10367 3655
rect 11152 3621 11186 3655
rect 1593 3553 1627 3587
rect 1860 3553 1894 3587
rect 4804 3553 4838 3587
rect 6745 3553 6779 3587
rect 8024 3553 8058 3587
rect 10241 3553 10275 3587
rect 12797 3553 12831 3587
rect 14381 3553 14415 3587
rect 15945 3553 15979 3587
rect 16497 3553 16531 3587
rect 17233 3553 17267 3587
rect 17785 3553 17819 3587
rect 19993 3553 20027 3587
rect 4537 3485 4571 3519
rect 6929 3485 6963 3519
rect 7757 3485 7791 3519
rect 10425 3485 10459 3519
rect 10701 3485 10735 3519
rect 10885 3485 10919 3519
rect 12541 3485 12575 3519
rect 14657 3485 14691 3519
rect 16129 3485 16163 3519
rect 16681 3485 16715 3519
rect 6377 3417 6411 3451
rect 15485 3417 15519 3451
rect 2973 3349 3007 3383
rect 5917 3349 5951 3383
rect 9137 3349 9171 3383
rect 9873 3349 9907 3383
rect 10701 3349 10735 3383
rect 12265 3349 12299 3383
rect 17417 3349 17451 3383
rect 17969 3349 18003 3383
rect 20177 3349 20211 3383
rect 3525 3145 3559 3179
rect 5273 3145 5307 3179
rect 5733 3145 5767 3179
rect 11345 3077 11379 3111
rect 13369 3077 13403 3111
rect 13461 3077 13495 3111
rect 3893 3009 3927 3043
rect 6285 3009 6319 3043
rect 9505 3009 9539 3043
rect 10609 3009 10643 3043
rect 11989 3009 12023 3043
rect 2145 2941 2179 2975
rect 2412 2941 2446 2975
rect 4160 2941 4194 2975
rect 7297 2941 7331 2975
rect 7564 2941 7598 2975
rect 10333 2941 10367 2975
rect 11805 2941 11839 2975
rect 12449 2941 12483 2975
rect 14013 3009 14047 3043
rect 18429 3009 18463 3043
rect 14473 2941 14507 2975
rect 15025 2941 15059 2975
rect 15761 2941 15795 2975
rect 16497 2941 16531 2975
rect 17049 2941 17083 2975
rect 18245 2941 18279 2975
rect 20545 2941 20579 2975
rect 9321 2873 9355 2907
rect 12725 2873 12759 2907
rect 13369 2873 13403 2907
rect 13921 2873 13955 2907
rect 15301 2873 15335 2907
rect 16037 2873 16071 2907
rect 6101 2805 6135 2839
rect 6193 2805 6227 2839
rect 8677 2805 8711 2839
rect 8953 2805 8987 2839
rect 9413 2805 9447 2839
rect 9965 2805 9999 2839
rect 10425 2805 10459 2839
rect 11713 2805 11747 2839
rect 13829 2805 13863 2839
rect 14657 2805 14691 2839
rect 16681 2805 16715 2839
rect 17233 2805 17267 2839
rect 20729 2805 20763 2839
rect 1961 2601 1995 2635
rect 2329 2601 2363 2635
rect 2421 2601 2455 2635
rect 3433 2601 3467 2635
rect 5365 2601 5399 2635
rect 5457 2601 5491 2635
rect 6929 2601 6963 2635
rect 7389 2601 7423 2635
rect 8401 2601 8435 2635
rect 9045 2601 9079 2635
rect 9781 2601 9815 2635
rect 12081 2601 12115 2635
rect 3341 2533 3375 2567
rect 8493 2533 8527 2567
rect 10149 2533 10183 2567
rect 7297 2465 7331 2499
rect 10793 2465 10827 2499
rect 11069 2465 11103 2499
rect 11529 2465 11563 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 13737 2465 13771 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 16037 2465 16071 2499
rect 16681 2465 16715 2499
rect 2605 2397 2639 2431
rect 3617 2397 3651 2431
rect 5549 2397 5583 2431
rect 7481 2397 7515 2431
rect 8677 2397 8711 2431
rect 10241 2397 10275 2431
rect 10425 2397 10459 2431
rect 2973 2329 3007 2363
rect 4997 2329 5031 2363
rect 8033 2329 8067 2363
rect 11713 2261 11747 2295
rect 12817 2261 12851 2295
rect 13369 2261 13403 2295
rect 13921 2261 13955 2295
rect 14473 2261 14507 2295
rect 15025 2261 15059 2295
rect 15669 2261 15703 2295
rect 16221 2261 16255 2295
rect 16865 2261 16899 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 7009 19499 7067 19505
rect 7009 19496 7021 19499
rect 4120 19468 7021 19496
rect 4120 19456 4126 19468
rect 7009 19465 7021 19468
rect 7055 19465 7067 19499
rect 7009 19459 7067 19465
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 1854 19292 1860 19304
rect 1811 19264 1860 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 2314 19292 2320 19304
rect 2275 19264 2320 19292
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 7190 19292 7196 19304
rect 6871 19264 7196 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 2866 19224 2872 19236
rect 1964 19196 2872 19224
rect 1964 19165 1992 19196
rect 2866 19184 2872 19196
rect 2924 19184 2930 19236
rect 1949 19159 2007 19165
rect 1949 19125 1961 19159
rect 1995 19125 2007 19159
rect 1949 19119 2007 19125
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2774 19156 2780 19168
rect 2547 19128 2780 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 3786 18912 3792 18964
rect 3844 18952 3850 18964
rect 7469 18955 7527 18961
rect 7469 18952 7481 18955
rect 3844 18924 7481 18952
rect 3844 18912 3850 18924
rect 7469 18921 7481 18924
rect 7515 18921 7527 18955
rect 7469 18915 7527 18921
rect 2314 18844 2320 18896
rect 2372 18884 2378 18896
rect 3145 18887 3203 18893
rect 3145 18884 3157 18887
rect 2372 18856 3157 18884
rect 2372 18844 2378 18856
rect 3145 18853 3157 18856
rect 3191 18853 3203 18887
rect 3145 18847 3203 18853
rect 2133 18819 2191 18825
rect 2133 18785 2145 18819
rect 2179 18816 2191 18819
rect 2869 18819 2927 18825
rect 2179 18788 2452 18816
rect 2179 18785 2191 18788
rect 2133 18779 2191 18785
rect 1762 18708 1768 18760
rect 1820 18748 1826 18760
rect 2317 18751 2375 18757
rect 2317 18748 2329 18751
rect 1820 18720 2329 18748
rect 1820 18708 1826 18720
rect 2317 18717 2329 18720
rect 2363 18717 2375 18751
rect 2317 18711 2375 18717
rect 2424 18680 2452 18788
rect 2869 18785 2881 18819
rect 2915 18785 2927 18819
rect 7282 18816 7288 18828
rect 7243 18788 7288 18816
rect 2869 18779 2927 18785
rect 2884 18748 2912 18779
rect 7282 18776 7288 18788
rect 7340 18776 7346 18828
rect 8478 18748 8484 18760
rect 2884 18720 8484 18748
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 7742 18680 7748 18692
rect 2424 18652 7748 18680
rect 7742 18640 7748 18652
rect 7800 18640 7806 18692
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 2774 18408 2780 18420
rect 2547 18380 2780 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 3050 18408 3056 18420
rect 3011 18380 3056 18408
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 7190 18272 7196 18284
rect 7151 18244 7196 18272
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18204 1823 18207
rect 2038 18204 2044 18216
rect 1811 18176 2044 18204
rect 1811 18173 1823 18176
rect 1765 18167 1823 18173
rect 2038 18164 2044 18176
rect 2096 18164 2102 18216
rect 2314 18204 2320 18216
rect 2275 18176 2320 18204
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18173 2927 18207
rect 2869 18167 2927 18173
rect 7009 18207 7067 18213
rect 7009 18173 7021 18207
rect 7055 18204 7067 18207
rect 7098 18204 7104 18216
rect 7055 18176 7104 18204
rect 7055 18173 7067 18176
rect 7009 18167 7067 18173
rect 2884 18136 2912 18167
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 10318 18136 10324 18148
rect 2884 18108 10324 18136
rect 10318 18096 10324 18108
rect 10376 18096 10382 18148
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 1857 17867 1915 17873
rect 1857 17864 1869 17867
rect 1820 17836 1869 17864
rect 1820 17824 1826 17836
rect 1857 17833 1869 17836
rect 1903 17833 1915 17867
rect 3142 17864 3148 17876
rect 3103 17836 3148 17864
rect 1857 17827 1915 17833
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 2314 17756 2320 17808
rect 2372 17796 2378 17808
rect 2501 17799 2559 17805
rect 2501 17796 2513 17799
rect 2372 17768 2513 17796
rect 2372 17756 2378 17768
rect 2501 17765 2513 17768
rect 2547 17765 2559 17799
rect 2501 17759 2559 17765
rect 7282 17756 7288 17808
rect 7340 17796 7346 17808
rect 8021 17799 8079 17805
rect 8021 17796 8033 17799
rect 7340 17768 8033 17796
rect 7340 17756 7346 17768
rect 8021 17765 8033 17768
rect 8067 17765 8079 17799
rect 10318 17796 10324 17808
rect 10279 17768 10324 17796
rect 8021 17759 8079 17765
rect 10318 17756 10324 17768
rect 10376 17756 10382 17808
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17728 1731 17731
rect 1946 17728 1952 17740
rect 1719 17700 1952 17728
rect 1719 17697 1731 17700
rect 1673 17691 1731 17697
rect 1946 17688 1952 17700
rect 2004 17688 2010 17740
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17697 2283 17731
rect 2225 17691 2283 17697
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 7650 17728 7656 17740
rect 3007 17700 7656 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 2240 17660 2268 17691
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 7745 17731 7803 17737
rect 7745 17697 7757 17731
rect 7791 17728 7803 17731
rect 9214 17728 9220 17740
rect 7791 17700 9220 17728
rect 7791 17697 7803 17700
rect 7745 17691 7803 17697
rect 9214 17688 9220 17700
rect 9272 17688 9278 17740
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 10686 17728 10692 17740
rect 10091 17700 10692 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 7282 17660 7288 17672
rect 2240 17632 7288 17660
rect 7282 17620 7288 17632
rect 7340 17620 7346 17672
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1762 17320 1768 17332
rect 1723 17292 1768 17320
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 10686 17320 10692 17332
rect 10647 17292 10692 17320
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 2038 17212 2044 17264
rect 2096 17252 2102 17264
rect 5537 17255 5595 17261
rect 2096 17224 2360 17252
rect 2096 17212 2102 17224
rect 2332 17193 2360 17224
rect 5537 17221 5549 17255
rect 5583 17221 5595 17255
rect 5537 17215 5595 17221
rect 9125 17255 9183 17261
rect 9125 17221 9137 17255
rect 9171 17221 9183 17255
rect 9125 17215 9183 17221
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17153 2375 17187
rect 5552 17184 5580 17215
rect 6178 17184 6184 17196
rect 2317 17147 2375 17153
rect 2424 17156 5580 17184
rect 6139 17156 6184 17184
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17116 1639 17119
rect 2038 17116 2044 17128
rect 1627 17088 2044 17116
rect 1627 17085 1639 17088
rect 1581 17079 1639 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17116 2191 17119
rect 2424 17116 2452 17156
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 8573 17187 8631 17193
rect 8573 17184 8585 17187
rect 7708 17156 8585 17184
rect 7708 17144 7714 17156
rect 8573 17153 8585 17156
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 2179 17088 2452 17116
rect 2869 17119 2927 17125
rect 2179 17085 2191 17088
rect 2133 17079 2191 17085
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 8389 17119 8447 17125
rect 2915 17088 8340 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 1946 17008 1952 17060
rect 2004 17048 2010 17060
rect 3145 17051 3203 17057
rect 3145 17048 3157 17051
rect 2004 17020 3157 17048
rect 2004 17008 2010 17020
rect 3145 17017 3157 17020
rect 3191 17017 3203 17051
rect 7190 17048 7196 17060
rect 3145 17011 3203 17017
rect 3896 17020 7196 17048
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 3896 16980 3924 17020
rect 7190 17008 7196 17020
rect 7248 17008 7254 17060
rect 8312 17048 8340 17088
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 9140 17116 9168 17215
rect 9766 17184 9772 17196
rect 9727 17156 9772 17184
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 11330 17184 11336 17196
rect 11291 17156 11336 17184
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 8435 17088 9168 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 8754 17048 8760 17060
rect 8312 17020 8760 17048
rect 8754 17008 8760 17020
rect 8812 17008 8818 17060
rect 11057 17051 11115 17057
rect 11057 17017 11069 17051
rect 11103 17048 11115 17051
rect 11701 17051 11759 17057
rect 11701 17048 11713 17051
rect 11103 17020 11713 17048
rect 11103 17017 11115 17020
rect 11057 17011 11115 17017
rect 11701 17017 11713 17020
rect 11747 17017 11759 17051
rect 11701 17011 11759 17017
rect 1728 16952 3924 16980
rect 3973 16983 4031 16989
rect 1728 16940 1734 16952
rect 3973 16949 3985 16983
rect 4019 16980 4031 16983
rect 5534 16980 5540 16992
rect 4019 16952 5540 16980
rect 4019 16949 4031 16952
rect 3973 16943 4031 16949
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 5902 16980 5908 16992
rect 5863 16952 5908 16980
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 6052 16952 6097 16980
rect 6052 16940 6058 16952
rect 9122 16940 9128 16992
rect 9180 16980 9186 16992
rect 9493 16983 9551 16989
rect 9493 16980 9505 16983
rect 9180 16952 9505 16980
rect 9180 16940 9186 16952
rect 9493 16949 9505 16952
rect 9539 16949 9551 16983
rect 9493 16943 9551 16949
rect 9585 16983 9643 16989
rect 9585 16949 9597 16983
rect 9631 16980 9643 16983
rect 9674 16980 9680 16992
rect 9631 16952 9680 16980
rect 9631 16949 9643 16952
rect 9585 16943 9643 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 3326 16776 3332 16788
rect 3287 16748 3332 16776
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 5721 16779 5779 16785
rect 5721 16745 5733 16779
rect 5767 16776 5779 16779
rect 5767 16748 6132 16776
rect 5767 16745 5779 16748
rect 5721 16739 5779 16745
rect 1854 16668 1860 16720
rect 1912 16708 1918 16720
rect 1949 16711 2007 16717
rect 1949 16708 1961 16711
rect 1912 16680 1961 16708
rect 1912 16668 1918 16680
rect 1949 16677 1961 16680
rect 1995 16677 2007 16711
rect 1949 16671 2007 16677
rect 2038 16668 2044 16720
rect 2096 16708 2102 16720
rect 2685 16711 2743 16717
rect 2685 16708 2697 16711
rect 2096 16680 2697 16708
rect 2096 16668 2102 16680
rect 2685 16677 2697 16680
rect 2731 16677 2743 16711
rect 5166 16708 5172 16720
rect 2685 16671 2743 16677
rect 2976 16680 5172 16708
rect 1670 16640 1676 16652
rect 1631 16612 1676 16640
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 2409 16643 2467 16649
rect 2409 16609 2421 16643
rect 2455 16640 2467 16643
rect 2976 16640 3004 16680
rect 5166 16668 5172 16680
rect 5224 16668 5230 16720
rect 3142 16640 3148 16652
rect 2455 16612 3004 16640
rect 3103 16612 3148 16640
rect 2455 16609 2467 16612
rect 2409 16603 2467 16609
rect 3142 16600 3148 16612
rect 3200 16600 3206 16652
rect 3510 16600 3516 16652
rect 3568 16640 3574 16652
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 3568 16612 4353 16640
rect 3568 16600 3574 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 4608 16643 4666 16649
rect 4608 16609 4620 16643
rect 4654 16640 4666 16643
rect 4890 16640 4896 16652
rect 4654 16612 4896 16640
rect 4654 16609 4666 16612
rect 4608 16603 4666 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 6104 16640 6132 16748
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 7377 16779 7435 16785
rect 7377 16776 7389 16779
rect 6236 16748 7389 16776
rect 6236 16736 6242 16748
rect 7377 16745 7389 16748
rect 7423 16745 7435 16779
rect 9122 16776 9128 16788
rect 9083 16748 9128 16776
rect 7377 16739 7435 16745
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 10410 16776 10416 16788
rect 9824 16748 10416 16776
rect 9824 16736 9830 16748
rect 10410 16736 10416 16748
rect 10468 16776 10474 16788
rect 11057 16779 11115 16785
rect 11057 16776 11069 16779
rect 10468 16748 11069 16776
rect 10468 16736 10474 16748
rect 11057 16745 11069 16748
rect 11103 16745 11115 16779
rect 11057 16739 11115 16745
rect 11330 16736 11336 16788
rect 11388 16776 11394 16788
rect 12713 16779 12771 16785
rect 12713 16776 12725 16779
rect 11388 16748 12725 16776
rect 11388 16736 11394 16748
rect 12713 16745 12725 16748
rect 12759 16776 12771 16779
rect 18966 16776 18972 16788
rect 12759 16748 18972 16776
rect 12759 16745 12771 16748
rect 12713 16739 12771 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 10134 16708 10140 16720
rect 9692 16680 10140 16708
rect 6270 16649 6276 16652
rect 6264 16640 6276 16649
rect 6104 16612 6276 16640
rect 6264 16603 6276 16612
rect 6270 16600 6276 16603
rect 6328 16600 6334 16652
rect 9692 16649 9720 16680
rect 10134 16668 10140 16680
rect 10192 16708 10198 16720
rect 10192 16680 11376 16708
rect 10192 16668 10198 16680
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 9944 16643 10002 16649
rect 9944 16609 9956 16643
rect 9990 16640 10002 16643
rect 10226 16640 10232 16652
rect 9990 16612 10232 16640
rect 9990 16609 10002 16612
rect 9944 16603 10002 16609
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 11348 16649 11376 16680
rect 11606 16649 11612 16652
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 11600 16603 11612 16649
rect 11664 16640 11670 16652
rect 11664 16612 11700 16640
rect 11606 16600 11612 16603
rect 11664 16600 11670 16612
rect 5810 16532 5816 16584
rect 5868 16572 5874 16584
rect 5997 16575 6055 16581
rect 5997 16572 6009 16575
rect 5868 16544 6009 16572
rect 5868 16532 5874 16544
rect 5997 16541 6009 16544
rect 6043 16541 6055 16575
rect 7926 16572 7932 16584
rect 7887 16544 7932 16572
rect 5997 16535 6055 16541
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 2958 16232 2964 16244
rect 2919 16204 2964 16232
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 4890 16232 4896 16244
rect 4851 16204 4896 16232
rect 4890 16192 4896 16204
rect 4948 16192 4954 16244
rect 5166 16232 5172 16244
rect 5127 16204 5172 16232
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 7190 16232 7196 16244
rect 7151 16204 7196 16232
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 11517 16235 11575 16241
rect 11517 16201 11529 16235
rect 11563 16232 11575 16235
rect 11606 16232 11612 16244
rect 11563 16204 11612 16232
rect 11563 16201 11575 16204
rect 11517 16195 11575 16201
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 2317 16099 2375 16105
rect 2317 16065 2329 16099
rect 2363 16096 2375 16099
rect 3142 16096 3148 16108
rect 2363 16068 3148 16096
rect 2363 16065 2375 16068
rect 2317 16059 2375 16065
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 3510 16096 3516 16108
rect 3471 16068 3516 16096
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 4908 16096 4936 16192
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 4908 16068 5733 16096
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 5721 16059 5779 16065
rect 5902 16056 5908 16108
rect 5960 16096 5966 16108
rect 6181 16099 6239 16105
rect 6181 16096 6193 16099
rect 5960 16068 6193 16096
rect 5960 16056 5966 16068
rect 6181 16065 6193 16068
rect 6227 16065 6239 16099
rect 6181 16059 6239 16065
rect 7837 16099 7895 16105
rect 7837 16065 7849 16099
rect 7883 16096 7895 16099
rect 10134 16096 10140 16108
rect 7883 16068 8156 16096
rect 10095 16068 10140 16096
rect 7883 16065 7895 16068
rect 7837 16059 7895 16065
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 15997 1547 16031
rect 2038 16028 2044 16040
rect 1999 16000 2044 16028
rect 1489 15991 1547 15997
rect 1504 15960 1532 15991
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2682 15988 2688 16040
rect 2740 16028 2746 16040
rect 2777 16031 2835 16037
rect 2777 16028 2789 16031
rect 2740 16000 2789 16028
rect 2740 15988 2746 16000
rect 2777 15997 2789 16000
rect 2823 15997 2835 16031
rect 5534 16028 5540 16040
rect 5495 16000 5540 16028
rect 2777 15991 2835 15997
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 7561 16031 7619 16037
rect 7561 15997 7573 16031
rect 7607 16028 7619 16031
rect 7926 16028 7932 16040
rect 7607 16000 7932 16028
rect 7607 15997 7619 16000
rect 7561 15991 7619 15997
rect 7926 15988 7932 16000
rect 7984 15988 7990 16040
rect 3780 15963 3838 15969
rect 1504 15932 2820 15960
rect 2792 15904 2820 15932
rect 3780 15929 3792 15963
rect 3826 15960 3838 15963
rect 4154 15960 4160 15972
rect 3826 15932 4160 15960
rect 3826 15929 3838 15932
rect 3780 15923 3838 15929
rect 4154 15920 4160 15932
rect 4212 15960 4218 15972
rect 4798 15960 4804 15972
rect 4212 15932 4804 15960
rect 4212 15920 4218 15932
rect 4798 15920 4804 15932
rect 4856 15920 4862 15972
rect 8128 15960 8156 16068
rect 10134 16056 10140 16068
rect 10192 16056 10198 16108
rect 8202 15988 8208 16040
rect 8260 16037 8266 16040
rect 10410 16037 10416 16040
rect 8260 16028 8270 16037
rect 10404 16028 10416 16037
rect 8260 16000 8305 16028
rect 10371 16000 10416 16028
rect 8260 15991 8270 16000
rect 10404 15991 10416 16000
rect 8260 15988 8266 15991
rect 10410 15988 10416 15991
rect 10468 15988 10474 16040
rect 8472 15963 8530 15969
rect 8472 15960 8484 15963
rect 8128 15932 8484 15960
rect 8472 15929 8484 15932
rect 8518 15960 8530 15963
rect 8938 15960 8944 15972
rect 8518 15932 8944 15960
rect 8518 15929 8530 15932
rect 8472 15923 8530 15929
rect 8938 15920 8944 15932
rect 8996 15920 9002 15972
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 2774 15852 2780 15904
rect 2832 15852 2838 15904
rect 5626 15892 5632 15904
rect 5587 15864 5632 15892
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 7650 15892 7656 15904
rect 7611 15864 7656 15892
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 9585 15895 9643 15901
rect 9585 15861 9597 15895
rect 9631 15892 9643 15895
rect 10226 15892 10232 15904
rect 9631 15864 10232 15892
rect 9631 15861 9643 15864
rect 9585 15855 9643 15861
rect 10226 15852 10232 15864
rect 10284 15852 10290 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 2777 15691 2835 15697
rect 2777 15688 2789 15691
rect 2096 15660 2789 15688
rect 2096 15648 2102 15660
rect 2777 15657 2789 15660
rect 2823 15657 2835 15691
rect 2777 15651 2835 15657
rect 4249 15691 4307 15697
rect 4249 15657 4261 15691
rect 4295 15688 4307 15691
rect 5626 15688 5632 15700
rect 4295 15660 5632 15688
rect 4295 15657 4307 15660
rect 4249 15651 4307 15657
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 8938 15688 8944 15700
rect 8899 15660 8944 15688
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10965 15691 11023 15697
rect 10965 15657 10977 15691
rect 11011 15688 11023 15691
rect 11146 15688 11152 15700
rect 11011 15660 11152 15688
rect 11011 15657 11023 15660
rect 10965 15651 11023 15657
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 2317 15623 2375 15629
rect 2317 15589 2329 15623
rect 2363 15620 2375 15623
rect 2682 15620 2688 15632
rect 2363 15592 2688 15620
rect 2363 15589 2375 15592
rect 2317 15583 2375 15589
rect 2682 15580 2688 15592
rect 2740 15580 2746 15632
rect 4062 15620 4068 15632
rect 2976 15592 4068 15620
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 1946 15552 1952 15564
rect 1535 15524 1952 15552
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15552 2099 15555
rect 2976 15552 3004 15592
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 6178 15629 6184 15632
rect 6172 15620 6184 15629
rect 6139 15592 6184 15620
rect 6172 15583 6184 15592
rect 6178 15580 6184 15583
rect 6236 15580 6242 15632
rect 8202 15620 8208 15632
rect 7484 15592 8208 15620
rect 3142 15552 3148 15564
rect 2087 15524 3004 15552
rect 3103 15524 3148 15552
rect 2087 15521 2099 15524
rect 2041 15515 2099 15521
rect 3142 15512 3148 15524
rect 3200 15512 3206 15564
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15552 3295 15555
rect 4246 15552 4252 15564
rect 3283 15524 4252 15552
rect 3283 15521 3295 15524
rect 3237 15515 3295 15521
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 4709 15555 4767 15561
rect 4709 15521 4721 15555
rect 4755 15552 4767 15555
rect 4755 15524 5212 15552
rect 4755 15521 4767 15524
rect 4709 15515 4767 15521
rect 3326 15444 3332 15496
rect 3384 15484 3390 15496
rect 3384 15456 3429 15484
rect 3384 15444 3390 15456
rect 4632 15416 4660 15515
rect 4798 15484 4804 15496
rect 4759 15456 4804 15484
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 4632 15388 4844 15416
rect 4816 15360 4844 15388
rect 4798 15308 4804 15360
rect 4856 15308 4862 15360
rect 5184 15357 5212 15524
rect 5810 15512 5816 15564
rect 5868 15552 5874 15564
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 5868 15524 5917 15552
rect 5868 15512 5874 15524
rect 5905 15521 5917 15524
rect 5951 15552 5963 15555
rect 7484 15552 7512 15592
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 10137 15623 10195 15629
rect 10137 15589 10149 15623
rect 10183 15620 10195 15623
rect 10597 15623 10655 15629
rect 10597 15620 10609 15623
rect 10183 15592 10609 15620
rect 10183 15589 10195 15592
rect 10137 15583 10195 15589
rect 10597 15589 10609 15592
rect 10643 15620 10655 15623
rect 11882 15620 11888 15632
rect 10643 15592 11888 15620
rect 10643 15589 10655 15592
rect 10597 15583 10655 15589
rect 11882 15580 11888 15592
rect 11940 15580 11946 15632
rect 5951 15524 7512 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 7484 15496 7512 15524
rect 7828 15555 7886 15561
rect 7828 15521 7840 15555
rect 7874 15552 7886 15555
rect 8662 15552 8668 15564
rect 7874 15524 8668 15552
rect 7874 15521 7886 15524
rect 7828 15515 7886 15521
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 10042 15552 10048 15564
rect 10003 15524 10048 15552
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 11333 15555 11391 15561
rect 11333 15552 11345 15555
rect 11112 15524 11345 15552
rect 11112 15512 11118 15524
rect 11333 15521 11345 15524
rect 11379 15521 11391 15555
rect 11333 15515 11391 15521
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 7561 15487 7619 15493
rect 7561 15484 7573 15487
rect 7524 15456 7573 15484
rect 7524 15444 7530 15456
rect 7561 15453 7573 15456
rect 7607 15453 7619 15487
rect 7561 15447 7619 15453
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 11425 15487 11483 15493
rect 10284 15456 10329 15484
rect 10284 15444 10290 15456
rect 11425 15453 11437 15487
rect 11471 15453 11483 15487
rect 11606 15484 11612 15496
rect 11567 15456 11612 15484
rect 11425 15447 11483 15453
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 6546 15348 6552 15360
rect 5215 15320 6552 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 7285 15351 7343 15357
rect 7285 15317 7297 15351
rect 7331 15348 7343 15351
rect 7558 15348 7564 15360
rect 7331 15320 7564 15348
rect 7331 15317 7343 15320
rect 7285 15311 7343 15317
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 11440 15348 11468 15447
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 11790 15348 11796 15360
rect 11440 15320 11796 15348
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 3510 15144 3516 15156
rect 2792 15116 3516 15144
rect 1670 15076 1676 15088
rect 1631 15048 1676 15076
rect 1670 15036 1676 15048
rect 1728 15036 1734 15088
rect 1946 14968 1952 15020
rect 2004 15008 2010 15020
rect 2792 15017 2820 15116
rect 3510 15104 3516 15116
rect 3568 15104 3574 15156
rect 4154 15144 4160 15156
rect 4115 15116 4160 15144
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 4246 15104 4252 15156
rect 4304 15144 4310 15156
rect 4617 15147 4675 15153
rect 4617 15144 4629 15147
rect 4304 15116 4629 15144
rect 4304 15104 4310 15116
rect 4617 15113 4629 15116
rect 4663 15113 4675 15147
rect 4617 15107 4675 15113
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 5994 15144 6000 15156
rect 5767 15116 6000 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 5994 15104 6000 15116
rect 6052 15104 6058 15156
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 7708 15116 8033 15144
rect 7708 15104 7714 15116
rect 8021 15113 8033 15116
rect 8067 15113 8079 15147
rect 8662 15144 8668 15156
rect 8575 15116 8668 15144
rect 8021 15107 8079 15113
rect 8662 15104 8668 15116
rect 8720 15144 8726 15156
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 8720 15116 10609 15144
rect 8720 15104 8726 15116
rect 10597 15113 10609 15116
rect 10643 15113 10655 15147
rect 10597 15107 10655 15113
rect 7009 15079 7067 15085
rect 7009 15045 7021 15079
rect 7055 15076 7067 15079
rect 8570 15076 8576 15088
rect 7055 15048 8576 15076
rect 7055 15045 7067 15048
rect 7009 15039 7067 15045
rect 8570 15036 8576 15048
rect 8628 15036 8634 15088
rect 2225 15011 2283 15017
rect 2225 15008 2237 15011
rect 2004 14980 2237 15008
rect 2004 14968 2010 14980
rect 2225 14977 2237 14980
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 2777 14971 2835 14977
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14909 1547 14943
rect 1489 14903 1547 14909
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 2792 14940 2820 14971
rect 4706 14968 4712 15020
rect 4764 15008 4770 15020
rect 5169 15011 5227 15017
rect 5169 15008 5181 15011
rect 4764 14980 5181 15008
rect 4764 14968 4770 14980
rect 5169 14977 5181 14980
rect 5215 14977 5227 15011
rect 6270 15008 6276 15020
rect 6231 14980 6276 15008
rect 5169 14971 5227 14977
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 7558 15008 7564 15020
rect 7519 14980 7564 15008
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 8680 15017 8708 15104
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 2866 14940 2872 14952
rect 2087 14912 2452 14940
rect 2792 14912 2872 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 1504 14804 1532 14903
rect 2424 14872 2452 14912
rect 2866 14900 2872 14912
rect 2924 14900 2930 14952
rect 3044 14943 3102 14949
rect 3044 14909 3056 14943
rect 3090 14940 3102 14943
rect 3326 14940 3332 14952
rect 3090 14912 3332 14940
rect 3090 14909 3102 14912
rect 3044 14903 3102 14909
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 4985 14943 5043 14949
rect 4985 14909 4997 14943
rect 5031 14940 5043 14943
rect 5994 14940 6000 14952
rect 5031 14912 6000 14940
rect 5031 14909 5043 14912
rect 4985 14903 5043 14909
rect 5994 14900 6000 14912
rect 6052 14900 6058 14952
rect 6181 14943 6239 14949
rect 6181 14909 6193 14943
rect 6227 14940 6239 14943
rect 7650 14940 7656 14952
rect 6227 14912 7656 14940
rect 6227 14909 6239 14912
rect 6181 14903 6239 14909
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 8260 14912 9229 14940
rect 8260 14900 8266 14912
rect 9217 14909 9229 14912
rect 9263 14909 9275 14943
rect 11054 14940 11060 14952
rect 9217 14903 9275 14909
rect 9324 14912 11060 14940
rect 4246 14872 4252 14884
rect 2424 14844 4252 14872
rect 4246 14832 4252 14844
rect 4304 14832 4310 14884
rect 6914 14832 6920 14884
rect 6972 14872 6978 14884
rect 7469 14875 7527 14881
rect 7469 14872 7481 14875
rect 6972 14844 7481 14872
rect 6972 14832 6978 14844
rect 7469 14841 7481 14844
rect 7515 14872 7527 14875
rect 7837 14875 7895 14881
rect 7837 14872 7849 14875
rect 7515 14844 7849 14872
rect 7515 14841 7527 14844
rect 7469 14835 7527 14841
rect 7837 14841 7849 14844
rect 7883 14841 7895 14875
rect 9324 14872 9352 14912
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 7837 14835 7895 14841
rect 8220 14844 9352 14872
rect 2682 14804 2688 14816
rect 1504 14776 2688 14804
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 4525 14807 4583 14813
rect 4525 14773 4537 14807
rect 4571 14804 4583 14807
rect 5077 14807 5135 14813
rect 5077 14804 5089 14807
rect 4571 14776 5089 14804
rect 4571 14773 4583 14776
rect 4525 14767 4583 14773
rect 5077 14773 5089 14776
rect 5123 14804 5135 14807
rect 5810 14804 5816 14816
rect 5123 14776 5816 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 6086 14804 6092 14816
rect 6047 14776 6092 14804
rect 6086 14764 6092 14776
rect 6144 14764 6150 14816
rect 7190 14764 7196 14816
rect 7248 14804 7254 14816
rect 7377 14807 7435 14813
rect 7377 14804 7389 14807
rect 7248 14776 7389 14804
rect 7248 14764 7254 14776
rect 7377 14773 7389 14776
rect 7423 14804 7435 14807
rect 8220 14804 8248 14844
rect 9398 14832 9404 14884
rect 9456 14881 9462 14884
rect 9456 14875 9520 14881
rect 9456 14841 9474 14875
rect 9508 14841 9520 14875
rect 9456 14835 9520 14841
rect 9456 14832 9462 14835
rect 7423 14776 8248 14804
rect 7423 14773 7435 14776
rect 7377 14767 7435 14773
rect 8294 14764 8300 14816
rect 8352 14804 8358 14816
rect 8389 14807 8447 14813
rect 8389 14804 8401 14807
rect 8352 14776 8401 14804
rect 8352 14764 8358 14776
rect 8389 14773 8401 14776
rect 8435 14773 8447 14807
rect 8389 14767 8447 14773
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 8941 14807 8999 14813
rect 8941 14804 8953 14807
rect 8527 14776 8953 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 8941 14773 8953 14776
rect 8987 14804 8999 14807
rect 10870 14804 10876 14816
rect 8987 14776 10876 14804
rect 8987 14773 8999 14776
rect 8941 14767 8999 14773
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 3384 14572 3433 14600
rect 3384 14560 3390 14572
rect 3421 14569 3433 14572
rect 3467 14569 3479 14603
rect 3421 14563 3479 14569
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 4212 14572 4445 14600
rect 4212 14560 4218 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 4433 14563 4491 14569
rect 4890 14560 4896 14612
rect 4948 14600 4954 14612
rect 8294 14600 8300 14612
rect 4948 14572 8300 14600
rect 4948 14560 4954 14572
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 10042 14600 10048 14612
rect 8496 14572 10048 14600
rect 2308 14535 2366 14541
rect 2308 14501 2320 14535
rect 2354 14532 2366 14535
rect 4706 14532 4712 14544
rect 2354 14504 4712 14532
rect 2354 14501 2366 14504
rect 2308 14495 2366 14501
rect 4706 14492 4712 14504
rect 4764 14492 4770 14544
rect 4801 14535 4859 14541
rect 4801 14501 4813 14535
rect 4847 14532 4859 14535
rect 5902 14532 5908 14544
rect 4847 14504 5908 14532
rect 4847 14501 4859 14504
rect 4801 14495 4859 14501
rect 5902 14492 5908 14504
rect 5960 14492 5966 14544
rect 6632 14535 6690 14541
rect 6632 14501 6644 14535
rect 6678 14532 6690 14535
rect 7558 14532 7564 14544
rect 6678 14504 7564 14532
rect 6678 14501 6690 14504
rect 6632 14495 6690 14501
rect 7558 14492 7564 14504
rect 7616 14492 7622 14544
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 2041 14467 2099 14473
rect 2041 14433 2053 14467
rect 2087 14464 2099 14467
rect 2866 14464 2872 14476
rect 2087 14436 2872 14464
rect 2087 14433 2099 14436
rect 2041 14427 2099 14433
rect 2866 14424 2872 14436
rect 2924 14424 2930 14476
rect 4724 14328 4752 14492
rect 4893 14467 4951 14473
rect 4893 14433 4905 14467
rect 4939 14464 4951 14467
rect 5718 14464 5724 14476
rect 4939 14436 5724 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 6086 14424 6092 14476
rect 6144 14464 6150 14476
rect 6454 14464 6460 14476
rect 6144 14436 6460 14464
rect 6144 14424 6150 14436
rect 6454 14424 6460 14436
rect 6512 14464 6518 14476
rect 8496 14464 8524 14572
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 9033 14535 9091 14541
rect 9033 14501 9045 14535
rect 9079 14532 9091 14535
rect 9674 14532 9680 14544
rect 9079 14504 9680 14532
rect 9079 14501 9091 14504
rect 9033 14495 9091 14501
rect 9674 14492 9680 14504
rect 9732 14492 9738 14544
rect 10134 14532 10140 14544
rect 9876 14504 10140 14532
rect 6512 14436 8524 14464
rect 8941 14467 8999 14473
rect 6512 14424 6518 14436
rect 8941 14433 8953 14467
rect 8987 14464 8999 14467
rect 9306 14464 9312 14476
rect 8987 14436 9312 14464
rect 8987 14433 8999 14436
rect 8941 14427 8999 14433
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 9876 14464 9904 14504
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 9950 14473 9956 14476
rect 9692 14436 9904 14464
rect 4982 14396 4988 14408
rect 4943 14368 4988 14396
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14365 5963 14399
rect 6362 14396 6368 14408
rect 6323 14368 6368 14396
rect 5905 14359 5963 14365
rect 5626 14328 5632 14340
rect 4724 14300 5632 14328
rect 5626 14288 5632 14300
rect 5684 14288 5690 14340
rect 5920 14260 5948 14359
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14396 9275 14399
rect 9398 14396 9404 14408
rect 9263 14368 9404 14396
rect 9263 14365 9275 14368
rect 9217 14359 9275 14365
rect 9398 14356 9404 14368
rect 9456 14356 9462 14408
rect 9692 14405 9720 14436
rect 9944 14427 9956 14473
rect 10008 14464 10014 14476
rect 10008 14436 10044 14464
rect 9950 14424 9956 14427
rect 10008 14424 10014 14436
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 7745 14331 7803 14337
rect 7745 14297 7757 14331
rect 7791 14328 7803 14331
rect 8294 14328 8300 14340
rect 7791 14300 8300 14328
rect 7791 14297 7803 14300
rect 7745 14291 7803 14297
rect 8294 14288 8300 14300
rect 8352 14328 8358 14340
rect 9122 14328 9128 14340
rect 8352 14300 9128 14328
rect 8352 14288 8358 14300
rect 9122 14288 9128 14300
rect 9180 14288 9186 14340
rect 7374 14260 7380 14272
rect 5920 14232 7380 14260
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 8573 14263 8631 14269
rect 8573 14260 8585 14263
rect 8536 14232 8585 14260
rect 8536 14220 8542 14232
rect 8573 14229 8585 14232
rect 8619 14229 8631 14263
rect 9416 14260 9444 14356
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 9416 14232 11069 14260
rect 8573 14223 8631 14229
rect 11057 14229 11069 14232
rect 11103 14229 11115 14263
rect 11057 14223 11115 14229
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 3418 14056 3424 14068
rect 3379 14028 3424 14056
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 5626 14056 5632 14068
rect 5587 14028 5632 14056
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 5994 14016 6000 14068
rect 6052 14056 6058 14068
rect 8386 14056 8392 14068
rect 6052 14028 8392 14056
rect 6052 14016 6058 14028
rect 8386 14016 8392 14028
rect 8444 14056 8450 14068
rect 9582 14056 9588 14068
rect 8444 14028 9588 14056
rect 8444 14016 8450 14028
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 9950 14056 9956 14068
rect 9911 14028 9956 14056
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 3326 13920 3332 13932
rect 2087 13892 3332 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 4062 13920 4068 13932
rect 3568 13892 4068 13920
rect 3568 13880 3574 13892
rect 4062 13880 4068 13892
rect 4120 13920 4126 13932
rect 4249 13923 4307 13929
rect 4249 13920 4261 13923
rect 4120 13892 4261 13920
rect 4120 13880 4126 13892
rect 4249 13889 4261 13892
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 1765 13855 1823 13861
rect 1765 13821 1777 13855
rect 1811 13852 1823 13855
rect 1946 13852 1952 13864
rect 1811 13824 1952 13852
rect 1811 13821 1823 13824
rect 1765 13815 1823 13821
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 2547 13824 2636 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 2608 13784 2636 13824
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 2777 13855 2835 13861
rect 2777 13852 2789 13855
rect 2740 13824 2789 13852
rect 2740 13812 2746 13824
rect 2777 13821 2789 13824
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 3237 13855 3295 13861
rect 3237 13852 3249 13855
rect 2924 13824 3249 13852
rect 2924 13812 2930 13824
rect 3237 13821 3249 13824
rect 3283 13821 3295 13855
rect 3237 13815 3295 13821
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 6822 13852 6828 13864
rect 6420 13824 6828 13852
rect 6420 13812 6426 13824
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7092 13855 7150 13861
rect 7092 13821 7104 13855
rect 7138 13852 7150 13855
rect 8294 13852 8300 13864
rect 7138 13824 8300 13852
rect 7138 13821 7150 13824
rect 7092 13815 7150 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 3050 13784 3056 13796
rect 2608 13756 3056 13784
rect 3050 13744 3056 13756
rect 3108 13744 3114 13796
rect 3142 13744 3148 13796
rect 3200 13784 3206 13796
rect 3789 13787 3847 13793
rect 3789 13784 3801 13787
rect 3200 13756 3801 13784
rect 3200 13744 3206 13756
rect 3789 13753 3801 13756
rect 3835 13753 3847 13787
rect 3789 13747 3847 13753
rect 4516 13787 4574 13793
rect 4516 13753 4528 13787
rect 4562 13784 4574 13787
rect 4982 13784 4988 13796
rect 4562 13756 4988 13784
rect 4562 13753 4574 13756
rect 4516 13747 4574 13753
rect 4982 13744 4988 13756
rect 5040 13784 5046 13796
rect 5442 13784 5448 13796
rect 5040 13756 5448 13784
rect 5040 13744 5046 13756
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 5902 13784 5908 13796
rect 5863 13756 5908 13784
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 6840 13784 6868 13812
rect 7466 13784 7472 13796
rect 6840 13756 7472 13784
rect 7466 13744 7472 13756
rect 7524 13784 7530 13796
rect 8588 13784 8616 13815
rect 9306 13812 9312 13864
rect 9364 13852 9370 13864
rect 9364 13824 10272 13852
rect 9364 13812 9370 13824
rect 7524 13756 8616 13784
rect 8840 13787 8898 13793
rect 7524 13744 7530 13756
rect 8840 13753 8852 13787
rect 8886 13784 8898 13787
rect 9030 13784 9036 13796
rect 8886 13756 9036 13784
rect 8886 13753 8898 13756
rect 8840 13747 8898 13753
rect 9030 13744 9036 13756
rect 9088 13744 9094 13796
rect 10244 13793 10272 13824
rect 10229 13787 10287 13793
rect 10229 13753 10241 13787
rect 10275 13753 10287 13787
rect 10229 13747 10287 13753
rect 8202 13716 8208 13728
rect 8163 13688 8208 13716
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 3510 13512 3516 13524
rect 3471 13484 3516 13512
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 5442 13512 5448 13524
rect 5403 13484 5448 13512
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6089 13515 6147 13521
rect 6089 13481 6101 13515
rect 6135 13512 6147 13515
rect 6362 13512 6368 13524
rect 6135 13484 6368 13512
rect 6135 13481 6147 13484
rect 6089 13475 6147 13481
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 7432 13484 8953 13512
rect 7432 13472 7438 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 8941 13475 8999 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 1486 13404 1492 13456
rect 1544 13444 1550 13456
rect 2133 13447 2191 13453
rect 2133 13444 2145 13447
rect 1544 13416 2145 13444
rect 1544 13404 1550 13416
rect 2133 13413 2145 13416
rect 2179 13413 2191 13447
rect 4154 13444 4160 13456
rect 2133 13407 2191 13413
rect 2608 13416 4160 13444
rect 1854 13376 1860 13388
rect 1815 13348 1860 13376
rect 1854 13336 1860 13348
rect 1912 13336 1918 13388
rect 2608 13385 2636 13416
rect 4154 13404 4160 13416
rect 4212 13404 4218 13456
rect 4332 13447 4390 13453
rect 4332 13413 4344 13447
rect 4378 13444 4390 13447
rect 5994 13444 6000 13456
rect 4378 13416 6000 13444
rect 4378 13413 4390 13416
rect 4332 13407 4390 13413
rect 5994 13404 6000 13416
rect 6052 13444 6058 13456
rect 6052 13416 6224 13444
rect 6052 13404 6058 13416
rect 2593 13379 2651 13385
rect 2593 13345 2605 13379
rect 2639 13345 2651 13379
rect 3326 13376 3332 13388
rect 3287 13348 3332 13376
rect 2593 13339 2651 13345
rect 3326 13336 3332 13348
rect 3384 13336 3390 13388
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 6196 13376 6224 13416
rect 8570 13404 8576 13456
rect 8628 13444 8634 13456
rect 9033 13447 9091 13453
rect 9033 13444 9045 13447
rect 8628 13416 9045 13444
rect 8628 13404 8634 13416
rect 9033 13413 9045 13416
rect 9079 13413 9091 13447
rect 9033 13407 9091 13413
rect 9582 13404 9588 13456
rect 9640 13444 9646 13456
rect 10045 13447 10103 13453
rect 10045 13444 10057 13447
rect 9640 13416 10057 13444
rect 9640 13404 9646 13416
rect 10045 13413 10057 13416
rect 10091 13413 10103 13447
rect 10045 13407 10103 13413
rect 6196 13348 6316 13376
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 6178 13308 6184 13320
rect 2832 13280 2877 13308
rect 6139 13280 6184 13308
rect 2832 13268 2838 13280
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 6288 13317 6316 13348
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 7064 13348 7297 13376
rect 7064 13336 7070 13348
rect 7285 13345 7297 13348
rect 7331 13345 7343 13379
rect 7285 13339 7343 13345
rect 7929 13379 7987 13385
rect 7929 13345 7941 13379
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13376 8079 13379
rect 8754 13376 8760 13388
rect 8067 13348 8760 13376
rect 8067 13345 8079 13348
rect 8021 13339 8079 13345
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 7944 13308 7972 13339
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10318 13376 10324 13388
rect 10183 13348 10324 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 7524 13280 7972 13308
rect 8205 13311 8263 13317
rect 7524 13268 7530 13280
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 8846 13308 8852 13320
rect 8251 13280 8852 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 9122 13268 9128 13320
rect 9180 13308 9186 13320
rect 9180 13280 9225 13308
rect 9180 13268 9186 13280
rect 9950 13268 9956 13320
rect 10008 13308 10014 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 10008 13280 10241 13308
rect 10008 13268 10014 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 7561 13243 7619 13249
rect 7561 13209 7573 13243
rect 7607 13240 7619 13243
rect 7742 13240 7748 13252
rect 7607 13212 7748 13240
rect 7607 13209 7619 13212
rect 7561 13203 7619 13209
rect 7742 13200 7748 13212
rect 7800 13200 7806 13252
rect 8573 13243 8631 13249
rect 8573 13209 8585 13243
rect 8619 13240 8631 13243
rect 8662 13240 8668 13252
rect 8619 13212 8668 13240
rect 8619 13209 8631 13212
rect 8573 13203 8631 13209
rect 8662 13200 8668 13212
rect 8720 13200 8726 13252
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 7101 13175 7159 13181
rect 7101 13172 7113 13175
rect 6880 13144 7113 13172
rect 6880 13132 6886 13144
rect 7101 13141 7113 13144
rect 7147 13141 7159 13175
rect 7101 13135 7159 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 5994 12968 6000 12980
rect 5955 12940 6000 12968
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 9030 12968 9036 12980
rect 8991 12940 9036 12968
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 10045 12971 10103 12977
rect 10045 12968 10057 12971
rect 9732 12940 10057 12968
rect 9732 12928 9738 12940
rect 10045 12937 10057 12940
rect 10091 12968 10103 12971
rect 10134 12968 10140 12980
rect 10091 12940 10140 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 2866 12900 2872 12912
rect 2056 12872 2872 12900
rect 2056 12841 2084 12872
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 6822 12860 6828 12912
rect 6880 12900 6886 12912
rect 6880 12872 7696 12900
rect 6880 12860 6886 12872
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12801 2099 12835
rect 2041 12795 2099 12801
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12832 7251 12835
rect 7466 12832 7472 12844
rect 7239 12804 7472 12832
rect 7239 12801 7251 12804
rect 7193 12795 7251 12801
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7668 12841 7696 12872
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 1762 12764 1768 12776
rect 1723 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 2682 12724 2688 12776
rect 2740 12764 2746 12776
rect 2869 12767 2927 12773
rect 2869 12764 2881 12767
rect 2740 12736 2881 12764
rect 2740 12724 2746 12736
rect 2869 12733 2881 12736
rect 2915 12764 2927 12767
rect 4062 12764 4068 12776
rect 2915 12736 4068 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 4062 12724 4068 12736
rect 4120 12764 4126 12776
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4120 12736 4629 12764
rect 4120 12724 4126 12736
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 4617 12727 4675 12733
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 7742 12764 7748 12776
rect 7340 12736 7748 12764
rect 7340 12724 7346 12736
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 10229 12767 10287 12773
rect 10229 12733 10241 12767
rect 10275 12764 10287 12767
rect 10778 12764 10784 12776
rect 10275 12736 10784 12764
rect 10275 12733 10287 12736
rect 10229 12727 10287 12733
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 2774 12656 2780 12708
rect 2832 12696 2838 12708
rect 3114 12699 3172 12705
rect 3114 12696 3126 12699
rect 2832 12668 3126 12696
rect 2832 12656 2838 12668
rect 3114 12665 3126 12668
rect 3160 12665 3172 12699
rect 3114 12659 3172 12665
rect 4884 12699 4942 12705
rect 4884 12665 4896 12699
rect 4930 12696 4942 12699
rect 5166 12696 5172 12708
rect 4930 12668 5172 12696
rect 4930 12665 4942 12668
rect 4884 12659 4942 12665
rect 5166 12656 5172 12668
rect 5224 12656 5230 12708
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 6362 12696 6368 12708
rect 5592 12668 6368 12696
rect 5592 12656 5598 12668
rect 6362 12656 6368 12668
rect 6420 12656 6426 12708
rect 7920 12699 7978 12705
rect 7920 12665 7932 12699
rect 7966 12696 7978 12699
rect 8662 12696 8668 12708
rect 7966 12668 8668 12696
rect 7966 12665 7978 12668
rect 7920 12659 7978 12665
rect 8662 12656 8668 12668
rect 8720 12656 8726 12708
rect 4249 12631 4307 12637
rect 4249 12597 4261 12631
rect 4295 12628 4307 12631
rect 4706 12628 4712 12640
rect 4295 12600 4712 12628
rect 4295 12597 4307 12600
rect 4249 12591 4307 12597
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 6270 12628 6276 12640
rect 6231 12600 6276 12628
rect 6270 12588 6276 12600
rect 6328 12588 6334 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1670 12424 1676 12436
rect 1631 12396 1676 12424
rect 1670 12384 1676 12396
rect 1728 12384 1734 12436
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 2041 12427 2099 12433
rect 2041 12424 2053 12427
rect 1912 12396 2053 12424
rect 1912 12384 1918 12396
rect 2041 12393 2053 12396
rect 2087 12393 2099 12427
rect 2041 12387 2099 12393
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4525 12427 4583 12433
rect 4525 12424 4537 12427
rect 4212 12396 4537 12424
rect 4212 12384 4218 12396
rect 4525 12393 4537 12396
rect 4571 12393 4583 12427
rect 4525 12387 4583 12393
rect 4893 12427 4951 12433
rect 4893 12393 4905 12427
rect 4939 12424 4951 12427
rect 6270 12424 6276 12436
rect 4939 12396 6276 12424
rect 4939 12393 4951 12396
rect 4893 12387 4951 12393
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 6362 12384 6368 12436
rect 6420 12384 6426 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7558 12424 7564 12436
rect 6972 12396 7564 12424
rect 6972 12384 6978 12396
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 9677 12427 9735 12433
rect 9677 12424 9689 12427
rect 8812 12396 9689 12424
rect 8812 12384 8818 12396
rect 9677 12393 9689 12396
rect 9723 12393 9735 12427
rect 9677 12387 9735 12393
rect 1504 12328 4384 12356
rect 1504 12297 1532 12328
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12257 1547 12291
rect 1489 12251 1547 12257
rect 2409 12291 2467 12297
rect 2409 12257 2421 12291
rect 2455 12288 2467 12291
rect 3694 12288 3700 12300
rect 2455 12260 3700 12288
rect 2455 12257 2467 12260
rect 2409 12251 2467 12257
rect 3694 12248 3700 12260
rect 3752 12248 3758 12300
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 2501 12223 2559 12229
rect 2501 12220 2513 12223
rect 1452 12192 2513 12220
rect 1452 12180 1458 12192
rect 2501 12189 2513 12192
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 2774 12220 2780 12232
rect 2731 12192 2780 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 2774 12180 2780 12192
rect 2832 12220 2838 12232
rect 2958 12220 2964 12232
rect 2832 12192 2964 12220
rect 2832 12180 2838 12192
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 4062 12220 4068 12232
rect 3099 12192 4068 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4249 12155 4307 12161
rect 4249 12152 4261 12155
rect 4212 12124 4261 12152
rect 4212 12112 4218 12124
rect 4249 12121 4261 12124
rect 4295 12121 4307 12155
rect 4356 12152 4384 12328
rect 5074 12316 5080 12368
rect 5132 12356 5138 12368
rect 6380 12356 6408 12384
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 5132 12328 5580 12356
rect 6380 12328 10057 12356
rect 5132 12316 5138 12328
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 5442 12288 5448 12300
rect 4479 12260 5448 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 5552 12297 5580 12328
rect 10045 12325 10057 12328
rect 10091 12325 10103 12359
rect 10045 12319 10103 12325
rect 5537 12291 5595 12297
rect 5537 12257 5549 12291
rect 5583 12257 5595 12291
rect 5537 12251 5595 12257
rect 5804 12291 5862 12297
rect 5804 12257 5816 12291
rect 5850 12288 5862 12291
rect 6362 12288 6368 12300
rect 5850 12260 6368 12288
rect 5850 12257 5862 12260
rect 5804 12251 5862 12257
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 7552 12291 7610 12297
rect 7552 12257 7564 12291
rect 7598 12288 7610 12291
rect 7834 12288 7840 12300
rect 7598 12260 7840 12288
rect 7598 12257 7610 12260
rect 7552 12251 7610 12257
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 8294 12248 8300 12300
rect 8352 12288 8358 12300
rect 19521 12291 19579 12297
rect 19521 12288 19533 12291
rect 8352 12260 19533 12288
rect 8352 12248 8358 12260
rect 19521 12257 19533 12260
rect 19567 12257 19579 12291
rect 19521 12251 19579 12257
rect 4982 12220 4988 12232
rect 4943 12192 4988 12220
rect 4982 12180 4988 12192
rect 5040 12180 5046 12232
rect 5166 12220 5172 12232
rect 5079 12192 5172 12220
rect 5166 12180 5172 12192
rect 5224 12220 5230 12232
rect 5224 12192 5488 12220
rect 5224 12180 5230 12192
rect 5258 12152 5264 12164
rect 4356 12124 5264 12152
rect 4249 12115 4307 12121
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 5460 12084 5488 12192
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6972 12192 7297 12220
rect 6972 12180 6978 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10008 12192 10149 12220
rect 10008 12180 10014 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 8662 12152 8668 12164
rect 8575 12124 8668 12152
rect 8662 12112 8668 12124
rect 8720 12152 8726 12164
rect 10244 12152 10272 12183
rect 8720 12124 10272 12152
rect 8720 12112 8726 12124
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 5460 12056 6929 12084
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 6917 12047 6975 12053
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12084 19763 12087
rect 20346 12084 20352 12096
rect 19751 12056 20352 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3421 11883 3479 11889
rect 3421 11880 3433 11883
rect 3016 11852 3433 11880
rect 3016 11840 3022 11852
rect 3421 11849 3433 11852
rect 3467 11849 3479 11883
rect 3694 11880 3700 11892
rect 3655 11852 3700 11880
rect 3421 11843 3479 11849
rect 3694 11840 3700 11852
rect 3752 11840 3758 11892
rect 3786 11840 3792 11892
rect 3844 11880 3850 11892
rect 5350 11880 5356 11892
rect 3844 11852 5356 11880
rect 3844 11840 3850 11852
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5500 11852 6224 11880
rect 5500 11840 5506 11852
rect 6196 11812 6224 11852
rect 6362 11840 6368 11892
rect 6420 11880 6426 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 6420 11852 6469 11880
rect 6420 11840 6426 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 7098 11840 7104 11892
rect 7156 11880 7162 11892
rect 7653 11883 7711 11889
rect 7653 11880 7665 11883
rect 7156 11852 7665 11880
rect 7156 11840 7162 11852
rect 7653 11849 7665 11852
rect 7699 11849 7711 11883
rect 7653 11843 7711 11849
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 7892 11852 10701 11880
rect 7892 11840 7898 11852
rect 7006 11812 7012 11824
rect 6196 11784 7012 11812
rect 7006 11772 7012 11784
rect 7064 11772 7070 11824
rect 8220 11753 8248 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 10689 11843 10747 11849
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 3160 11716 4261 11744
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 2041 11679 2099 11685
rect 2041 11676 2053 11679
rect 1636 11648 2053 11676
rect 1636 11636 1642 11648
rect 2041 11645 2053 11648
rect 2087 11645 2099 11679
rect 2041 11639 2099 11645
rect 2308 11679 2366 11685
rect 2308 11645 2320 11679
rect 2354 11676 2366 11679
rect 2866 11676 2872 11688
rect 2354 11648 2872 11676
rect 2354 11645 2366 11648
rect 2308 11639 2366 11645
rect 2056 11608 2084 11639
rect 2866 11636 2872 11648
rect 2924 11676 2930 11688
rect 3160 11676 3188 11716
rect 4249 11713 4261 11716
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11713 8263 11747
rect 9306 11744 9312 11756
rect 9267 11716 9312 11744
rect 8205 11707 8263 11713
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 4062 11676 4068 11688
rect 2924 11648 3188 11676
rect 4023 11648 4068 11676
rect 2924 11636 2930 11648
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4154 11636 4160 11688
rect 4212 11676 4218 11688
rect 5074 11676 5080 11688
rect 4212 11648 5080 11676
rect 4212 11636 4218 11648
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 7190 11676 7196 11688
rect 7151 11648 7196 11676
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 19061 11679 19119 11685
rect 19061 11645 19073 11679
rect 19107 11645 19119 11679
rect 19061 11639 19119 11645
rect 2682 11608 2688 11620
rect 2056 11580 2688 11608
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 5344 11611 5402 11617
rect 5344 11577 5356 11611
rect 5390 11608 5402 11611
rect 5718 11608 5724 11620
rect 5390 11580 5724 11608
rect 5390 11577 5402 11580
rect 5344 11571 5402 11577
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 8021 11611 8079 11617
rect 8021 11577 8033 11611
rect 8067 11608 8079 11611
rect 8665 11611 8723 11617
rect 8665 11608 8677 11611
rect 8067 11580 8677 11608
rect 8067 11577 8079 11580
rect 8021 11571 8079 11577
rect 8665 11577 8677 11580
rect 8711 11577 8723 11611
rect 8665 11571 8723 11577
rect 9306 11568 9312 11620
rect 9364 11608 9370 11620
rect 9576 11611 9634 11617
rect 9576 11608 9588 11611
rect 9364 11580 9588 11608
rect 9364 11568 9370 11580
rect 9576 11577 9588 11580
rect 9622 11608 9634 11611
rect 11054 11608 11060 11620
rect 9622 11580 11060 11608
rect 9622 11577 9634 11580
rect 9576 11571 9634 11577
rect 11054 11568 11060 11580
rect 11112 11568 11118 11620
rect 3694 11500 3700 11552
rect 3752 11540 3758 11552
rect 4062 11540 4068 11552
rect 3752 11512 4068 11540
rect 3752 11500 3758 11512
rect 4062 11500 4068 11512
rect 4120 11540 4126 11552
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 4120 11512 4169 11540
rect 4120 11500 4126 11512
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 8113 11543 8171 11549
rect 8113 11509 8125 11543
rect 8159 11540 8171 11543
rect 8570 11540 8576 11552
rect 8159 11512 8576 11540
rect 8159 11509 8171 11512
rect 8113 11503 8171 11509
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 19076 11540 19104 11639
rect 9180 11512 19104 11540
rect 19245 11543 19303 11549
rect 9180 11500 9186 11512
rect 19245 11509 19257 11543
rect 19291 11540 19303 11543
rect 19886 11540 19892 11552
rect 19291 11512 19892 11540
rect 19291 11509 19303 11512
rect 19245 11503 19303 11509
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1394 11336 1400 11348
rect 1355 11308 1400 11336
rect 1394 11296 1400 11308
rect 1452 11296 1458 11348
rect 1765 11339 1823 11345
rect 1765 11305 1777 11339
rect 1811 11336 1823 11339
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 1811 11308 2421 11336
rect 1811 11305 1823 11308
rect 1765 11299 1823 11305
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 2409 11299 2467 11305
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 4433 11339 4491 11345
rect 4433 11336 4445 11339
rect 4304 11308 4445 11336
rect 4304 11296 4310 11308
rect 4433 11305 4445 11308
rect 4479 11305 4491 11339
rect 4433 11299 4491 11305
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 5040 11308 5457 11336
rect 5040 11296 5046 11308
rect 5445 11305 5457 11308
rect 5491 11305 5503 11339
rect 5445 11299 5503 11305
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 7742 11336 7748 11348
rect 6963 11308 7748 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 9674 11336 9680 11348
rect 8720 11308 9680 11336
rect 8720 11296 8726 11308
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 11054 11336 11060 11348
rect 11015 11308 11060 11336
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 2866 11268 2872 11280
rect 2056 11240 2872 11268
rect 2056 11141 2084 11240
rect 2866 11228 2872 11240
rect 2924 11228 2930 11280
rect 2958 11228 2964 11280
rect 3016 11268 3022 11280
rect 3786 11268 3792 11280
rect 3016 11240 3792 11268
rect 3016 11228 3022 11240
rect 3786 11228 3792 11240
rect 3844 11228 3850 11280
rect 4801 11271 4859 11277
rect 4801 11237 4813 11271
rect 4847 11268 4859 11271
rect 6457 11271 6515 11277
rect 6457 11268 6469 11271
rect 4847 11240 6469 11268
rect 4847 11237 4859 11240
rect 4801 11231 4859 11237
rect 6457 11237 6469 11240
rect 6503 11237 6515 11271
rect 6457 11231 6515 11237
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 4246 11200 4252 11212
rect 2823 11172 4252 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 4246 11160 4252 11172
rect 4304 11200 4310 11212
rect 4893 11203 4951 11209
rect 4304 11172 4844 11200
rect 4304 11160 4310 11172
rect 4816 11144 4844 11172
rect 4893 11169 4905 11203
rect 4939 11200 4951 11203
rect 5166 11200 5172 11212
rect 4939 11172 5172 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5813 11203 5871 11209
rect 5813 11200 5825 11203
rect 5592 11172 5825 11200
rect 5592 11160 5598 11172
rect 5813 11169 5825 11172
rect 5859 11200 5871 11203
rect 6730 11200 6736 11212
rect 5859 11172 6736 11200
rect 5859 11169 5871 11172
rect 5813 11163 5871 11169
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 7282 11200 7288 11212
rect 7243 11172 7288 11200
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 8846 11200 8852 11212
rect 7423 11172 8852 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 8846 11160 8852 11172
rect 8904 11160 8910 11212
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 9766 11200 9772 11212
rect 9723 11172 9772 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11101 1915 11135
rect 1857 11095 1915 11101
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11101 2099 11135
rect 2041 11095 2099 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 2958 11132 2964 11144
rect 2915 11104 2964 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 1872 11064 1900 11095
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 2774 11064 2780 11076
rect 1872 11036 2780 11064
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 3068 10996 3096 11095
rect 4798 11092 4804 11144
rect 4856 11092 4862 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5718 11132 5724 11144
rect 5123 11104 5724 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5718 11092 5724 11104
rect 5776 11092 5782 11144
rect 5902 11132 5908 11144
rect 5863 11104 5908 11132
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6362 11132 6368 11144
rect 6135 11104 6368 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 7834 11132 7840 11144
rect 7607 11104 7840 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 6730 11024 6736 11076
rect 6788 11064 6794 11076
rect 8956 11064 8984 11163
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 9944 11203 10002 11209
rect 9944 11169 9956 11203
rect 9990 11200 10002 11203
rect 11146 11200 11152 11212
rect 9990 11172 11152 11200
rect 9990 11169 10002 11172
rect 9944 11163 10002 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 18598 11160 18604 11212
rect 18656 11209 18662 11212
rect 18656 11200 18665 11209
rect 18656 11172 18701 11200
rect 18656 11163 18665 11172
rect 18656 11160 18662 11163
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11132 9275 11135
rect 9306 11132 9312 11144
rect 9263 11104 9312 11132
rect 9263 11101 9275 11104
rect 9217 11095 9275 11101
rect 6788 11036 8984 11064
rect 9048 11064 9076 11095
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9398 11064 9404 11076
rect 9048 11036 9404 11064
rect 6788 11024 6794 11036
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 18785 11067 18843 11073
rect 18785 11033 18797 11067
rect 18831 11064 18843 11067
rect 19426 11064 19432 11076
rect 18831 11036 19432 11064
rect 18831 11033 18843 11036
rect 18785 11027 18843 11033
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 3326 10996 3332 11008
rect 3068 10968 3332 10996
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 4062 10956 4068 11008
rect 4120 10996 4126 11008
rect 11606 10996 11612 11008
rect 4120 10968 11612 10996
rect 4120 10956 4126 10968
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 2866 10752 2872 10804
rect 2924 10792 2930 10804
rect 2961 10795 3019 10801
rect 2961 10792 2973 10795
rect 2924 10764 2973 10792
rect 2924 10752 2930 10764
rect 2961 10761 2973 10764
rect 3007 10761 3019 10795
rect 2961 10755 3019 10761
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3108 10764 3709 10792
rect 3108 10752 3114 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 3697 10755 3755 10761
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 6457 10795 6515 10801
rect 6457 10792 6469 10795
rect 5776 10764 6469 10792
rect 5776 10752 5782 10764
rect 6457 10761 6469 10764
rect 6503 10761 6515 10795
rect 6457 10755 6515 10761
rect 9214 10752 9220 10804
rect 9272 10792 9278 10804
rect 9401 10795 9459 10801
rect 9401 10792 9413 10795
rect 9272 10764 9413 10792
rect 9272 10752 9278 10764
rect 9401 10761 9413 10764
rect 9447 10761 9459 10795
rect 9401 10755 9459 10761
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 9766 10724 9772 10736
rect 9171 10696 9772 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4890 10656 4896 10668
rect 4387 10628 4896 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5074 10656 5080 10668
rect 5035 10628 5080 10656
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 11146 10656 11152 10668
rect 10091 10628 11152 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 11664 10628 18276 10656
rect 11664 10616 11670 10628
rect 1848 10591 1906 10597
rect 1848 10557 1860 10591
rect 1894 10588 1906 10591
rect 3326 10588 3332 10600
rect 1894 10560 3332 10588
rect 1894 10557 1906 10560
rect 1848 10551 1906 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 6086 10588 6092 10600
rect 5276 10560 6092 10588
rect 4065 10523 4123 10529
rect 4065 10489 4077 10523
rect 4111 10520 4123 10523
rect 5276 10520 5304 10560
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 4111 10492 5304 10520
rect 5344 10523 5402 10529
rect 4111 10489 4123 10492
rect 4065 10483 4123 10489
rect 5344 10489 5356 10523
rect 5390 10520 5402 10523
rect 5442 10520 5448 10532
rect 5390 10492 5448 10520
rect 5390 10489 5402 10492
rect 5344 10483 5402 10489
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 6822 10452 6828 10464
rect 4203 10424 6828 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7190 10452 7196 10464
rect 7151 10424 7196 10452
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7392 10452 7420 10551
rect 7558 10548 7564 10600
rect 7616 10588 7622 10600
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7616 10560 7757 10588
rect 7616 10548 7622 10560
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 8001 10591 8059 10597
rect 8001 10588 8013 10591
rect 7892 10560 8013 10588
rect 7892 10548 7898 10560
rect 8001 10557 8013 10560
rect 8047 10588 8059 10591
rect 11054 10588 11060 10600
rect 8047 10560 8248 10588
rect 8047 10557 8059 10560
rect 8001 10551 8059 10557
rect 8220 10532 8248 10560
rect 9692 10560 10916 10588
rect 11015 10560 11060 10588
rect 8202 10480 8208 10532
rect 8260 10480 8266 10532
rect 9692 10452 9720 10560
rect 9769 10523 9827 10529
rect 9769 10489 9781 10523
rect 9815 10520 9827 10523
rect 10413 10523 10471 10529
rect 10413 10520 10425 10523
rect 9815 10492 10425 10520
rect 9815 10489 9827 10492
rect 9769 10483 9827 10489
rect 10413 10489 10425 10492
rect 10459 10489 10471 10523
rect 10888 10520 10916 10560
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 18248 10597 18276 10628
rect 18233 10591 18291 10597
rect 18233 10557 18245 10591
rect 18279 10557 18291 10591
rect 18233 10551 18291 10557
rect 11330 10520 11336 10532
rect 10888 10492 11336 10520
rect 10413 10483 10471 10489
rect 11330 10480 11336 10492
rect 11388 10480 11394 10532
rect 9858 10452 9864 10464
rect 7392 10424 9720 10452
rect 9819 10424 9864 10452
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 10873 10455 10931 10461
rect 10873 10452 10885 10455
rect 10836 10424 10885 10452
rect 10836 10412 10842 10424
rect 10873 10421 10885 10424
rect 10919 10421 10931 10455
rect 10873 10415 10931 10421
rect 18417 10455 18475 10461
rect 18417 10421 18429 10455
rect 18463 10452 18475 10455
rect 18690 10452 18696 10464
rect 18463 10424 18696 10452
rect 18463 10421 18475 10424
rect 18417 10415 18475 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2832 10220 2877 10248
rect 2832 10208 2838 10220
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5718 10248 5724 10260
rect 5500 10220 5724 10248
rect 5500 10208 5506 10220
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 8202 10248 8208 10260
rect 5828 10220 8064 10248
rect 8163 10220 8208 10248
rect 5828 10192 5856 10220
rect 3145 10183 3203 10189
rect 3145 10149 3157 10183
rect 3191 10180 3203 10183
rect 5810 10180 5816 10192
rect 3191 10152 5816 10180
rect 3191 10149 3203 10152
rect 3145 10143 3203 10149
rect 5810 10140 5816 10152
rect 5868 10140 5874 10192
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 4154 10112 4160 10124
rect 3283 10084 4160 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 4608 10115 4666 10121
rect 4608 10081 4620 10115
rect 4654 10112 4666 10115
rect 4890 10112 4896 10124
rect 4654 10084 4896 10112
rect 4654 10081 4666 10084
rect 4608 10075 4666 10081
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 6914 10112 6920 10124
rect 6871 10084 6920 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7092 10115 7150 10121
rect 7092 10081 7104 10115
rect 7138 10112 7150 10115
rect 7138 10084 7972 10112
rect 7138 10081 7150 10084
rect 7092 10075 7150 10081
rect 3326 10044 3332 10056
rect 3287 10016 3332 10044
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 3510 10004 3516 10056
rect 3568 10044 3574 10056
rect 4341 10047 4399 10053
rect 4341 10044 4353 10047
rect 3568 10016 4353 10044
rect 3568 10004 3574 10016
rect 4341 10013 4353 10016
rect 4387 10013 4399 10047
rect 4341 10007 4399 10013
rect 7944 9976 7972 10084
rect 8036 10044 8064 10220
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 9858 10248 9864 10260
rect 8619 10220 9864 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 11330 10248 11336 10260
rect 11291 10220 11336 10248
rect 11330 10208 11336 10220
rect 11388 10248 11394 10260
rect 11606 10248 11612 10260
rect 11388 10220 11612 10248
rect 11388 10208 11394 10220
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 8941 10115 8999 10121
rect 8941 10112 8953 10115
rect 8312 10084 8953 10112
rect 8312 10044 8340 10084
rect 8941 10081 8953 10084
rect 8987 10081 8999 10115
rect 8941 10075 8999 10081
rect 9861 10115 9919 10121
rect 9861 10081 9873 10115
rect 9907 10112 9919 10115
rect 10318 10112 10324 10124
rect 9907 10084 10324 10112
rect 9907 10081 9919 10084
rect 9861 10075 9919 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 9030 10044 9036 10056
rect 8036 10016 8340 10044
rect 8991 10016 9036 10044
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10044 9275 10047
rect 9766 10044 9772 10056
rect 9263 10016 9772 10044
rect 9263 10013 9275 10016
rect 9217 10007 9275 10013
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 8202 9976 8208 9988
rect 7944 9948 8208 9976
rect 8202 9936 8208 9948
rect 8260 9936 8266 9988
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 14366 9908 14372 9920
rect 4120 9880 14372 9908
rect 4120 9868 4126 9880
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 2961 9707 3019 9713
rect 2961 9673 2973 9707
rect 3007 9704 3019 9707
rect 3326 9704 3332 9716
rect 3007 9676 3332 9704
rect 3007 9673 3019 9676
rect 2961 9667 3019 9673
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 4890 9704 4896 9716
rect 3936 9676 4752 9704
rect 4851 9676 4896 9704
rect 3936 9664 3942 9676
rect 4724 9636 4752 9676
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 11057 9707 11115 9713
rect 5000 9676 11008 9704
rect 5000 9636 5028 9676
rect 5166 9636 5172 9648
rect 4724 9608 5028 9636
rect 5127 9608 5172 9636
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 6362 9636 6368 9648
rect 5368 9608 6368 9636
rect 4614 9528 4620 9580
rect 4672 9568 4678 9580
rect 5368 9568 5396 9608
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 6638 9596 6644 9648
rect 6696 9636 6702 9648
rect 6914 9636 6920 9648
rect 6696 9608 6920 9636
rect 6696 9596 6702 9608
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 7837 9639 7895 9645
rect 7837 9636 7849 9639
rect 7340 9608 7849 9636
rect 7340 9596 7346 9608
rect 7837 9605 7849 9608
rect 7883 9605 7895 9639
rect 8846 9636 8852 9648
rect 8807 9608 8852 9636
rect 7837 9599 7895 9605
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 10980 9636 11008 9676
rect 11057 9673 11069 9707
rect 11103 9704 11115 9707
rect 11146 9704 11152 9716
rect 11103 9676 11152 9704
rect 11103 9673 11115 9676
rect 11057 9667 11115 9673
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 10980 9608 11192 9636
rect 11164 9580 11192 9608
rect 5718 9568 5724 9580
rect 4672 9540 5396 9568
rect 5679 9540 5724 9568
rect 4672 9528 4678 9540
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7064 9540 7389 9568
rect 7064 9528 7070 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 8260 9540 8401 9568
rect 8260 9528 8266 9540
rect 8389 9537 8401 9540
rect 8435 9568 8447 9571
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 8435 9540 9413 9568
rect 8435 9537 8447 9540
rect 8389 9531 8447 9537
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 11146 9528 11152 9580
rect 11204 9528 11210 9580
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 1670 9500 1676 9512
rect 1627 9472 1676 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 1670 9460 1676 9472
rect 1728 9500 1734 9512
rect 3510 9500 3516 9512
rect 1728 9472 3516 9500
rect 1728 9460 1734 9472
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 3780 9503 3838 9509
rect 3780 9469 3792 9503
rect 3826 9500 3838 9503
rect 4706 9500 4712 9512
rect 3826 9472 4712 9500
rect 3826 9469 3838 9472
rect 3780 9463 3838 9469
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 5592 9472 5641 9500
rect 5592 9460 5598 9472
rect 5629 9469 5641 9472
rect 5675 9469 5687 9503
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 5629 9463 5687 9469
rect 6196 9472 7205 9500
rect 1848 9435 1906 9441
rect 1848 9401 1860 9435
rect 1894 9432 1906 9435
rect 2774 9432 2780 9444
rect 1894 9404 2780 9432
rect 1894 9401 1906 9404
rect 1848 9395 1906 9401
rect 2774 9392 2780 9404
rect 2832 9392 2838 9444
rect 5442 9392 5448 9444
rect 5500 9432 5506 9444
rect 6196 9432 6224 9472
rect 7193 9469 7205 9472
rect 7239 9500 7251 9503
rect 8478 9500 8484 9512
rect 7239 9472 8484 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 8478 9460 8484 9472
rect 8536 9500 8542 9512
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 8536 9472 9229 9500
rect 8536 9460 8542 9472
rect 9217 9469 9229 9472
rect 9263 9469 9275 9503
rect 9674 9500 9680 9512
rect 9635 9472 9680 9500
rect 9217 9463 9275 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 9933 9503 9991 9509
rect 9933 9500 9945 9503
rect 9824 9472 9945 9500
rect 9824 9460 9830 9472
rect 9933 9469 9945 9472
rect 9979 9469 9991 9503
rect 9933 9463 9991 9469
rect 5500 9404 6224 9432
rect 6273 9435 6331 9441
rect 5500 9392 5506 9404
rect 6273 9401 6285 9435
rect 6319 9432 6331 9435
rect 8205 9435 8263 9441
rect 8205 9432 8217 9435
rect 6319 9404 8217 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 8205 9401 8217 9404
rect 8251 9401 8263 9435
rect 8205 9395 8263 9401
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 9309 9435 9367 9441
rect 9309 9432 9321 9435
rect 8628 9404 9321 9432
rect 8628 9392 8634 9404
rect 9309 9401 9321 9404
rect 9355 9401 9367 9435
rect 9309 9395 9367 9401
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5810 9364 5816 9376
rect 5583 9336 5816 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6822 9364 6828 9376
rect 6783 9336 6828 9364
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 7374 9364 7380 9376
rect 7331 9336 7380 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 8297 9367 8355 9373
rect 8297 9364 8309 9367
rect 7800 9336 8309 9364
rect 7800 9324 7806 9336
rect 8297 9333 8309 9336
rect 8343 9333 8355 9367
rect 8297 9327 8355 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 4433 9163 4491 9169
rect 2832 9132 2877 9160
rect 2832 9120 2838 9132
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 4614 9160 4620 9172
rect 4479 9132 4620 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 5905 9163 5963 9169
rect 5905 9160 5917 9163
rect 4764 9132 5917 9160
rect 4764 9120 4770 9132
rect 5905 9129 5917 9132
rect 5951 9129 5963 9163
rect 6086 9160 6092 9172
rect 6047 9132 6092 9160
rect 5905 9123 5963 9129
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 6362 9120 6368 9172
rect 6420 9160 6426 9172
rect 8386 9160 8392 9172
rect 6420 9132 8392 9160
rect 6420 9120 6426 9132
rect 8386 9120 8392 9132
rect 8444 9160 8450 9172
rect 8481 9163 8539 9169
rect 8481 9160 8493 9163
rect 8444 9132 8493 9160
rect 8444 9120 8450 9132
rect 8481 9129 8493 9132
rect 8527 9129 8539 9163
rect 8481 9123 8539 9129
rect 1302 9052 1308 9104
rect 1360 9092 1366 9104
rect 3513 9095 3571 9101
rect 1360 9064 3464 9092
rect 1360 9052 1366 9064
rect 1664 9027 1722 9033
rect 1664 8993 1676 9027
rect 1710 9024 1722 9027
rect 2682 9024 2688 9036
rect 1710 8996 2688 9024
rect 1710 8993 1722 8996
rect 1664 8987 1722 8993
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 3436 9024 3464 9064
rect 3513 9061 3525 9095
rect 3559 9092 3571 9095
rect 6457 9095 6515 9101
rect 6457 9092 6469 9095
rect 3559 9064 6469 9092
rect 3559 9061 3571 9064
rect 3513 9055 3571 9061
rect 6457 9061 6469 9064
rect 6503 9061 6515 9095
rect 6457 9055 6515 9061
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 6788 9064 7696 9092
rect 6788 9052 6794 9064
rect 4522 9024 4528 9036
rect 3436 8996 4528 9024
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 5442 9024 5448 9036
rect 4632 8996 5448 9024
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8925 1455 8959
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 1397 8919 1455 8925
rect 1412 8820 1440 8919
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 4632 8956 4660 8996
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 5776 8996 7113 9024
rect 5776 8984 5782 8996
rect 7101 8993 7113 8996
rect 7147 8993 7159 9027
rect 7668 9024 7696 9064
rect 7834 9052 7840 9104
rect 7892 9092 7898 9104
rect 12066 9092 12072 9104
rect 7892 9064 12072 9092
rect 7892 9052 7898 9064
rect 12066 9052 12072 9064
rect 12124 9052 12130 9104
rect 8573 9027 8631 9033
rect 8573 9024 8585 9027
rect 7668 8996 8585 9024
rect 7101 8987 7159 8993
rect 8573 8993 8585 8996
rect 8619 8993 8631 9027
rect 8573 8987 8631 8993
rect 10128 9027 10186 9033
rect 10128 8993 10140 9027
rect 10174 9024 10186 9027
rect 10962 9024 10968 9036
rect 10174 8996 10968 9024
rect 10174 8993 10186 8996
rect 10128 8987 10186 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 3660 8928 4660 8956
rect 4709 8959 4767 8965
rect 3660 8916 3666 8928
rect 4709 8925 4721 8959
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 3234 8848 3240 8900
rect 3292 8888 3298 8900
rect 4724 8888 4752 8919
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 5040 8928 5549 8956
rect 5040 8916 5046 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 5644 8888 5672 8919
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 6420 8928 6561 8956
rect 6420 8916 6426 8928
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 7006 8956 7012 8968
rect 6687 8928 7012 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 3292 8860 5672 8888
rect 5905 8891 5963 8897
rect 3292 8848 3298 8860
rect 5905 8857 5917 8891
rect 5951 8888 5963 8891
rect 6656 8888 6684 8919
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 8803 8928 8892 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 5951 8860 6684 8888
rect 5951 8857 5963 8860
rect 5905 8851 5963 8857
rect 1670 8820 1676 8832
rect 1412 8792 1676 8820
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 4065 8823 4123 8829
rect 4065 8789 4077 8823
rect 4111 8820 4123 8823
rect 4798 8820 4804 8832
rect 4111 8792 4804 8820
rect 4111 8789 4123 8792
rect 4065 8783 4123 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 5077 8823 5135 8829
rect 5077 8820 5089 8823
rect 4948 8792 5089 8820
rect 4948 8780 4954 8792
rect 5077 8789 5089 8792
rect 5123 8789 5135 8823
rect 5077 8783 5135 8789
rect 5258 8780 5264 8832
rect 5316 8820 5322 8832
rect 7300 8820 7328 8919
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 8864 8888 8892 8928
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9732 8928 9873 8956
rect 9732 8916 9738 8928
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 8260 8860 8892 8888
rect 8260 8848 8266 8860
rect 5316 8792 7328 8820
rect 8113 8823 8171 8829
rect 5316 8780 5322 8792
rect 8113 8789 8125 8823
rect 8159 8820 8171 8823
rect 8294 8820 8300 8832
rect 8159 8792 8300 8820
rect 8159 8789 8171 8792
rect 8113 8783 8171 8789
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8864 8820 8892 8860
rect 11241 8823 11299 8829
rect 11241 8820 11253 8823
rect 8864 8792 11253 8820
rect 11241 8789 11253 8792
rect 11287 8789 11299 8823
rect 11241 8783 11299 8789
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 1762 8616 1768 8628
rect 1723 8588 1768 8616
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 2240 8588 4445 8616
rect 2240 8489 2268 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 5718 8616 5724 8628
rect 5679 8588 5724 8616
rect 4433 8579 4491 8585
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 7558 8616 7564 8628
rect 7300 8588 7564 8616
rect 2774 8548 2780 8560
rect 2424 8520 2780 8548
rect 2424 8489 2452 8520
rect 2774 8508 2780 8520
rect 2832 8508 2838 8560
rect 4157 8551 4215 8557
rect 4157 8517 4169 8551
rect 4203 8548 4215 8551
rect 7190 8548 7196 8560
rect 4203 8520 5028 8548
rect 4203 8517 4215 8520
rect 4157 8511 4215 8517
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8449 2283 8483
rect 2225 8443 2283 8449
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 2774 8412 2780 8424
rect 1728 8384 2780 8412
rect 1728 8372 1734 8384
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 4172 8412 4200 8511
rect 4890 8480 4896 8492
rect 4851 8452 4896 8480
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5000 8489 5028 8520
rect 5644 8520 7196 8548
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 4798 8412 4804 8424
rect 2976 8384 4200 8412
rect 4759 8384 4804 8412
rect 2682 8304 2688 8356
rect 2740 8344 2746 8356
rect 2976 8344 3004 8384
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 5644 8421 5672 8520
rect 7190 8508 7196 8520
rect 7248 8508 7254 8560
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 6546 8480 6552 8492
rect 6411 8452 6552 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 7300 8489 7328 8588
rect 7558 8576 7564 8588
rect 7616 8616 7622 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 7616 8588 9229 8616
rect 7616 8576 7622 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 10778 8616 10784 8628
rect 9217 8579 9275 8585
rect 9416 8588 10784 8616
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 6181 8415 6239 8421
rect 6181 8381 6193 8415
rect 6227 8412 6239 8415
rect 7098 8412 7104 8424
rect 6227 8384 7104 8412
rect 6227 8381 6239 8384
rect 6181 8375 6239 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 9122 8412 9128 8424
rect 7300 8384 9128 8412
rect 2740 8316 3004 8344
rect 3044 8347 3102 8353
rect 2740 8304 2746 8316
rect 3044 8313 3056 8347
rect 3090 8344 3102 8347
rect 3234 8344 3240 8356
rect 3090 8316 3240 8344
rect 3090 8313 3102 8316
rect 3044 8307 3102 8313
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 4062 8304 4068 8356
rect 4120 8344 4126 8356
rect 6825 8347 6883 8353
rect 4120 8316 6776 8344
rect 4120 8304 4126 8316
rect 2130 8276 2136 8288
rect 2091 8248 2136 8276
rect 2130 8236 2136 8248
rect 2188 8236 2194 8288
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5408 8248 5457 8276
rect 5408 8236 5414 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 6086 8276 6092 8288
rect 6047 8248 6092 8276
rect 5445 8239 5503 8245
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 6748 8276 6776 8316
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 7190 8344 7196 8356
rect 6871 8316 7196 8344
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 7300 8276 7328 8384
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 7552 8347 7610 8353
rect 7552 8313 7564 8347
rect 7598 8344 7610 8347
rect 8202 8344 8208 8356
rect 7598 8316 8208 8344
rect 7598 8313 7610 8316
rect 7552 8307 7610 8313
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 9232 8344 9260 8579
rect 9416 8421 9444 8588
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 10962 8616 10968 8628
rect 10923 8588 10968 8616
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 11112 8588 11253 8616
rect 11112 8576 11118 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 11241 8579 11299 8585
rect 9401 8415 9459 8421
rect 9401 8381 9413 8415
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 9674 8412 9680 8424
rect 9631 8384 9680 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 9600 8344 9628 8375
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 11425 8415 11483 8421
rect 11425 8381 11437 8415
rect 11471 8412 11483 8415
rect 11606 8412 11612 8424
rect 11471 8384 11612 8412
rect 11471 8381 11483 8384
rect 11425 8375 11483 8381
rect 11606 8372 11612 8384
rect 11664 8372 11670 8424
rect 9232 8316 9628 8344
rect 9852 8347 9910 8353
rect 9852 8313 9864 8347
rect 9898 8344 9910 8347
rect 11698 8344 11704 8356
rect 9898 8316 11704 8344
rect 9898 8313 9910 8316
rect 9852 8307 9910 8313
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 8662 8276 8668 8288
rect 6748 8248 7328 8276
rect 8623 8248 8668 8276
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2188 8044 2237 8072
rect 2188 8032 2194 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 2731 8044 4077 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4522 8032 4528 8084
rect 4580 8072 4586 8084
rect 4580 8044 5479 8072
rect 4580 8032 4586 8044
rect 2593 8007 2651 8013
rect 2593 7973 2605 8007
rect 2639 8004 2651 8007
rect 3050 8004 3056 8016
rect 2639 7976 3056 8004
rect 2639 7973 2651 7976
rect 2593 7967 2651 7973
rect 3050 7964 3056 7976
rect 3108 7964 3114 8016
rect 5350 8004 5356 8016
rect 3896 7976 5356 8004
rect 3896 7945 3924 7976
rect 5350 7964 5356 7976
rect 5408 7964 5414 8016
rect 5451 8004 5479 8044
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7929 8075 7987 8081
rect 7929 8072 7941 8075
rect 7156 8044 7941 8072
rect 7156 8032 7162 8044
rect 7929 8041 7941 8044
rect 7975 8041 7987 8075
rect 8294 8072 8300 8084
rect 8255 8044 8300 8072
rect 7929 8035 7987 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8072 10655 8075
rect 11149 8075 11207 8081
rect 11149 8072 11161 8075
rect 10643 8044 11161 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 11149 8041 11161 8044
rect 11195 8041 11207 8075
rect 11149 8035 11207 8041
rect 11698 8032 11704 8084
rect 11756 8072 11762 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 11756 8044 16681 8072
rect 11756 8032 11762 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 6454 8004 6460 8016
rect 5451 7976 6460 8004
rect 6454 7964 6460 7976
rect 6512 8004 6518 8016
rect 7377 8007 7435 8013
rect 7377 8004 7389 8007
rect 6512 7976 7389 8004
rect 6512 7964 6518 7976
rect 7377 7973 7389 7976
rect 7423 7973 7435 8007
rect 7742 8004 7748 8016
rect 7377 7967 7435 7973
rect 7484 7976 7748 8004
rect 3881 7939 3939 7945
rect 3881 7905 3893 7939
rect 3927 7905 3939 7939
rect 3881 7899 3939 7905
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 4890 7936 4896 7948
rect 4479 7908 4896 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 2682 7828 2688 7880
rect 2740 7868 2746 7880
rect 2777 7871 2835 7877
rect 2777 7868 2789 7871
rect 2740 7840 2789 7868
rect 2740 7828 2746 7840
rect 2777 7837 2789 7840
rect 2823 7837 2835 7871
rect 4448 7868 4476 7899
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 5436 7939 5494 7945
rect 5436 7905 5448 7939
rect 5482 7936 5494 7939
rect 7098 7936 7104 7948
rect 5482 7908 7104 7936
rect 5482 7905 5494 7908
rect 5436 7899 5494 7905
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7484 7936 7512 7976
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 10134 7964 10140 8016
rect 10192 8004 10198 8016
rect 11609 8007 11667 8013
rect 11609 8004 11621 8007
rect 10192 7976 11621 8004
rect 10192 7964 10198 7976
rect 11609 7973 11621 7976
rect 11655 7973 11667 8007
rect 11609 7967 11667 7973
rect 15556 8007 15614 8013
rect 15556 7973 15568 8007
rect 15602 8004 15614 8007
rect 15746 8004 15752 8016
rect 15602 7976 15752 8004
rect 15602 7973 15614 7976
rect 15556 7967 15614 7973
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 8202 7936 8208 7948
rect 7331 7908 7512 7936
rect 7576 7908 8208 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 2777 7831 2835 7837
rect 3160 7840 4476 7868
rect 2130 7760 2136 7812
rect 2188 7800 2194 7812
rect 3160 7800 3188 7840
rect 4522 7828 4528 7880
rect 4580 7868 4586 7880
rect 4709 7871 4767 7877
rect 4580 7840 4625 7868
rect 4580 7828 4586 7840
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 6362 7868 6368 7880
rect 6275 7840 6368 7868
rect 5169 7831 5227 7837
rect 2188 7772 3188 7800
rect 2188 7760 2194 7772
rect 3234 7760 3240 7812
rect 3292 7800 3298 7812
rect 4724 7800 4752 7831
rect 5184 7800 5212 7831
rect 6362 7828 6368 7840
rect 6420 7868 6426 7880
rect 7300 7868 7328 7899
rect 7576 7877 7604 7908
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 9723 7908 10517 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 11204 7908 11529 7936
rect 11204 7896 11210 7908
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 6420 7840 7328 7868
rect 7561 7871 7619 7877
rect 6420 7828 6426 7840
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8168 7840 8401 7868
rect 8168 7828 8174 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7868 8539 7871
rect 8662 7868 8668 7880
rect 8527 7840 8668 7868
rect 8527 7837 8539 7840
rect 8481 7831 8539 7837
rect 3292 7772 4752 7800
rect 4816 7772 5212 7800
rect 3292 7760 3298 7772
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 3697 7735 3755 7741
rect 3697 7732 3709 7735
rect 2832 7704 3709 7732
rect 2832 7692 2838 7704
rect 3697 7701 3709 7704
rect 3743 7732 3755 7735
rect 4816 7732 4844 7772
rect 3743 7704 4844 7732
rect 3743 7701 3755 7704
rect 3697 7695 3755 7701
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 6380 7732 6408 7828
rect 7098 7760 7104 7812
rect 7156 7800 7162 7812
rect 8496 7800 8524 7831
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 10962 7868 10968 7880
rect 10827 7840 10968 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11698 7828 11704 7880
rect 11756 7868 11762 7880
rect 11756 7840 11801 7868
rect 11756 7828 11762 7840
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15068 7840 15301 7868
rect 15068 7828 15074 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 7156 7772 8524 7800
rect 10137 7803 10195 7809
rect 7156 7760 7162 7772
rect 10137 7769 10149 7803
rect 10183 7800 10195 7803
rect 14642 7800 14648 7812
rect 10183 7772 14648 7800
rect 10183 7769 10195 7772
rect 10137 7763 10195 7769
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 6546 7732 6552 7744
rect 4948 7704 6408 7732
rect 6507 7704 6552 7732
rect 4948 7692 4954 7704
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7282 7732 7288 7744
rect 6963 7704 7288 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 1946 7528 1952 7540
rect 1907 7500 1952 7528
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 5626 7528 5632 7540
rect 3384 7500 5632 7528
rect 3384 7488 3390 7500
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 6086 7488 6092 7540
rect 6144 7528 6150 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6144 7500 6837 7528
rect 6144 7488 6150 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 8110 7528 8116 7540
rect 8071 7500 8116 7528
rect 6825 7491 6883 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 17862 7528 17868 7540
rect 10376 7500 17868 7528
rect 10376 7488 10382 7500
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 7098 7420 7104 7472
rect 7156 7460 7162 7472
rect 14277 7463 14335 7469
rect 7156 7432 7420 7460
rect 7156 7420 7162 7432
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 3602 7392 3608 7404
rect 3563 7364 3608 7392
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 7282 7392 7288 7404
rect 7243 7364 7288 7392
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7392 7401 7420 7432
rect 14277 7429 14289 7463
rect 14323 7460 14335 7463
rect 15654 7460 15660 7472
rect 14323 7432 15660 7460
rect 14323 7429 14335 7432
rect 14277 7423 14335 7429
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 8202 7352 8208 7404
rect 8260 7392 8266 7404
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8260 7364 8677 7392
rect 8260 7352 8266 7364
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 9732 7364 10333 7392
rect 9732 7352 9738 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7392 14979 7395
rect 15194 7392 15200 7404
rect 14967 7364 15200 7392
rect 14967 7361 14979 7364
rect 14921 7355 14979 7361
rect 4433 7327 4491 7333
rect 4433 7293 4445 7327
rect 4479 7324 4491 7327
rect 4522 7324 4528 7336
rect 4479 7296 4528 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 4700 7327 4758 7333
rect 4700 7293 4712 7327
rect 4746 7324 4758 7327
rect 6546 7324 6552 7336
rect 4746 7296 6552 7324
rect 4746 7293 4758 7296
rect 4700 7287 4758 7293
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 7190 7324 7196 7336
rect 7151 7296 7196 7324
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 10336 7324 10364 7355
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 10962 7324 10968 7336
rect 10336 7296 10968 7324
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 11112 7296 12173 7324
rect 11112 7284 11118 7296
rect 12161 7293 12173 7296
rect 12207 7293 12219 7327
rect 12161 7287 12219 7293
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 16945 7327 17003 7333
rect 16945 7324 16957 7327
rect 14700 7296 16957 7324
rect 14700 7284 14706 7296
rect 16945 7293 16957 7296
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 1486 7216 1492 7268
rect 1544 7256 1550 7268
rect 2317 7259 2375 7265
rect 2317 7256 2329 7259
rect 1544 7228 2329 7256
rect 1544 7216 1550 7228
rect 2317 7225 2329 7228
rect 2363 7225 2375 7259
rect 2317 7219 2375 7225
rect 4062 7216 4068 7268
rect 4120 7256 4126 7268
rect 9306 7256 9312 7268
rect 4120 7228 9312 7256
rect 4120 7216 4126 7228
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 10588 7259 10646 7265
rect 10588 7225 10600 7259
rect 10634 7256 10646 7259
rect 10778 7256 10784 7268
rect 10634 7228 10784 7256
rect 10634 7225 10646 7228
rect 10588 7219 10646 7225
rect 10778 7216 10784 7228
rect 10836 7216 10842 7268
rect 14458 7216 14464 7268
rect 14516 7256 14522 7268
rect 14737 7259 14795 7265
rect 14737 7256 14749 7259
rect 14516 7228 14749 7256
rect 14516 7216 14522 7228
rect 14737 7225 14749 7228
rect 14783 7225 14795 7259
rect 14737 7219 14795 7225
rect 17221 7259 17279 7265
rect 17221 7225 17233 7259
rect 17267 7256 17279 7259
rect 17770 7256 17776 7268
rect 17267 7228 17776 7256
rect 17267 7225 17279 7228
rect 17221 7219 17279 7225
rect 17770 7216 17776 7228
rect 17828 7216 17834 7268
rect 2409 7191 2467 7197
rect 2409 7157 2421 7191
rect 2455 7188 2467 7191
rect 2961 7191 3019 7197
rect 2961 7188 2973 7191
rect 2455 7160 2973 7188
rect 2455 7157 2467 7160
rect 2409 7151 2467 7157
rect 2961 7157 2973 7160
rect 3007 7157 3019 7191
rect 3326 7188 3332 7200
rect 3287 7160 3332 7188
rect 2961 7151 3019 7157
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 3418 7148 3424 7200
rect 3476 7188 3482 7200
rect 3476 7160 3521 7188
rect 3476 7148 3482 7160
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 4764 7160 5825 7188
rect 4764 7148 4770 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 5813 7151 5871 7157
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 7190 7188 7196 7200
rect 6319 7160 7196 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 8573 7191 8631 7197
rect 8573 7157 8585 7191
rect 8619 7188 8631 7191
rect 10502 7188 10508 7200
rect 8619 7160 10508 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 11698 7188 11704 7200
rect 11659 7160 11704 7188
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 11977 7191 12035 7197
rect 11977 7157 11989 7191
rect 12023 7188 12035 7191
rect 13170 7188 13176 7200
rect 12023 7160 13176 7188
rect 12023 7157 12035 7160
rect 11977 7151 12035 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 14182 7188 14188 7200
rect 13679 7160 14188 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 14645 7191 14703 7197
rect 14645 7188 14657 7191
rect 14424 7160 14657 7188
rect 14424 7148 14430 7160
rect 14645 7157 14657 7160
rect 14691 7157 14703 7191
rect 15562 7188 15568 7200
rect 15523 7160 15568 7188
rect 14645 7151 14703 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 4065 6987 4123 6993
rect 4065 6984 4077 6987
rect 3384 6956 4077 6984
rect 3384 6944 3390 6956
rect 4065 6953 4077 6956
rect 4111 6953 4123 6987
rect 4065 6947 4123 6953
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4433 6987 4491 6993
rect 4433 6984 4445 6987
rect 4304 6956 4445 6984
rect 4304 6944 4310 6956
rect 4433 6953 4445 6956
rect 4479 6953 4491 6987
rect 10778 6984 10784 6996
rect 10691 6956 10784 6984
rect 4433 6947 4491 6953
rect 10778 6944 10784 6956
rect 10836 6984 10842 6996
rect 14461 6987 14519 6993
rect 14461 6984 14473 6987
rect 10836 6956 14473 6984
rect 10836 6944 10842 6956
rect 14461 6953 14473 6956
rect 14507 6953 14519 6987
rect 14461 6947 14519 6953
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 10321 6919 10379 6925
rect 10321 6916 10333 6919
rect 4028 6888 10333 6916
rect 4028 6876 4034 6888
rect 10321 6885 10333 6888
rect 10367 6885 10379 6919
rect 10321 6879 10379 6885
rect 2216 6851 2274 6857
rect 2216 6817 2228 6851
rect 2262 6848 2274 6851
rect 2498 6848 2504 6860
rect 2262 6820 2504 6848
rect 2262 6817 2274 6820
rect 2216 6811 2274 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 4525 6851 4583 6857
rect 4525 6848 4537 6851
rect 3896 6820 4537 6848
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 1949 6783 2007 6789
rect 1949 6780 1961 6783
rect 1728 6752 1961 6780
rect 1728 6740 1734 6752
rect 1949 6749 1961 6752
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 3896 6780 3924 6820
rect 4525 6817 4537 6820
rect 4571 6817 4583 6851
rect 4525 6811 4583 6817
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 5350 6848 5356 6860
rect 4672 6820 5120 6848
rect 5311 6820 5356 6848
rect 4672 6808 4678 6820
rect 5092 6792 5120 6820
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5718 6857 5724 6860
rect 5712 6848 5724 6857
rect 5679 6820 5724 6848
rect 5712 6811 5724 6820
rect 5718 6808 5724 6811
rect 5776 6808 5782 6860
rect 7374 6857 7380 6860
rect 7357 6851 7380 6857
rect 7357 6848 7369 6851
rect 6840 6820 7369 6848
rect 3016 6752 3924 6780
rect 3016 6740 3022 6752
rect 3528 6724 3556 6752
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4246 6780 4252 6792
rect 4028 6752 4252 6780
rect 4028 6740 4034 6752
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5132 6752 5457 6780
rect 5132 6740 5138 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 3234 6672 3240 6724
rect 3292 6712 3298 6724
rect 3329 6715 3387 6721
rect 3329 6712 3341 6715
rect 3292 6684 3341 6712
rect 3292 6672 3298 6684
rect 3329 6681 3341 6684
rect 3375 6681 3387 6715
rect 3329 6675 3387 6681
rect 3510 6672 3516 6724
rect 3568 6672 3574 6724
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 6840 6721 6868 6820
rect 7357 6817 7369 6820
rect 7432 6848 7438 6860
rect 7432 6820 7505 6848
rect 7357 6811 7380 6817
rect 7374 6808 7380 6811
rect 7432 6808 7438 6820
rect 7098 6780 7104 6792
rect 7059 6752 7104 6780
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10192 6752 10425 6780
rect 10192 6740 10198 6752
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6780 10655 6783
rect 10796 6780 10824 6944
rect 11232 6919 11290 6925
rect 11232 6885 11244 6919
rect 11278 6916 11290 6919
rect 11698 6916 11704 6928
rect 11278 6888 11704 6916
rect 11278 6885 11290 6888
rect 11232 6879 11290 6885
rect 11698 6876 11704 6888
rect 11756 6876 11762 6928
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 13081 6851 13139 6857
rect 13081 6848 13093 6851
rect 12492 6820 13093 6848
rect 12492 6808 12498 6820
rect 13081 6817 13093 6820
rect 13127 6817 13139 6851
rect 13081 6811 13139 6817
rect 13348 6851 13406 6857
rect 13348 6817 13360 6851
rect 13394 6848 13406 6851
rect 13906 6848 13912 6860
rect 13394 6820 13912 6848
rect 13394 6817 13406 6820
rect 13348 6811 13406 6817
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15556 6851 15614 6857
rect 15556 6848 15568 6851
rect 15252 6820 15568 6848
rect 15252 6808 15258 6820
rect 15556 6817 15568 6820
rect 15602 6848 15614 6851
rect 16022 6848 16028 6860
rect 15602 6820 16028 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 16942 6848 16948 6860
rect 16903 6820 16948 6848
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 10962 6780 10968 6792
rect 10643 6752 10824 6780
rect 10923 6752 10968 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 12618 6780 12624 6792
rect 12579 6752 12624 6780
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 15068 6752 15301 6780
rect 15068 6740 15074 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17678 6780 17684 6792
rect 17267 6752 17684 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 6825 6715 6883 6721
rect 4120 6684 5304 6712
rect 4120 6672 4126 6684
rect 1578 6604 1584 6656
rect 1636 6644 1642 6656
rect 3694 6644 3700 6656
rect 1636 6616 3700 6644
rect 1636 6604 1642 6616
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 5169 6647 5227 6653
rect 5169 6644 5181 6647
rect 5132 6616 5181 6644
rect 5132 6604 5138 6616
rect 5169 6613 5181 6616
rect 5215 6613 5227 6647
rect 5276 6644 5304 6684
rect 6825 6681 6837 6715
rect 6871 6681 6883 6715
rect 9214 6712 9220 6724
rect 6825 6675 6883 6681
rect 8036 6684 9220 6712
rect 8036 6644 8064 6684
rect 9214 6672 9220 6684
rect 9272 6672 9278 6724
rect 9324 6684 11008 6712
rect 8478 6644 8484 6656
rect 5276 6616 8064 6644
rect 8439 6616 8484 6644
rect 5169 6607 5227 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 9324 6644 9352 6684
rect 8720 6616 9352 6644
rect 9953 6647 10011 6653
rect 8720 6604 8726 6616
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10778 6644 10784 6656
rect 9999 6616 10784 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 10980 6644 11008 6684
rect 11974 6644 11980 6656
rect 10980 6616 11980 6644
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12342 6644 12348 6656
rect 12303 6616 12348 6644
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16669 6647 16727 6653
rect 16669 6644 16681 6647
rect 15988 6616 16681 6644
rect 15988 6604 15994 6616
rect 16669 6613 16681 6616
rect 16715 6613 16727 6647
rect 16669 6607 16727 6613
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 2556 6412 2789 6440
rect 2556 6400 2562 6412
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 2777 6403 2835 6409
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 3602 6440 3608 6452
rect 3016 6412 3608 6440
rect 3016 6400 3022 6412
rect 3602 6400 3608 6412
rect 3660 6440 3666 6452
rect 4985 6443 5043 6449
rect 4985 6440 4997 6443
rect 3660 6412 4997 6440
rect 3660 6400 3666 6412
rect 4985 6409 4997 6412
rect 5031 6409 5043 6443
rect 4985 6403 5043 6409
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 12342 6440 12348 6452
rect 5776 6412 12348 6440
rect 5776 6400 5782 6412
rect 4890 6264 4896 6316
rect 4948 6304 4954 6316
rect 5810 6304 5816 6316
rect 4948 6276 5816 6304
rect 4948 6264 4954 6276
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 6288 6313 6316 6412
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 13906 6440 13912 6452
rect 12544 6412 13768 6440
rect 13867 6412 13912 6440
rect 7098 6332 7104 6384
rect 7156 6372 7162 6384
rect 7156 6344 8248 6372
rect 7156 6332 7162 6344
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6273 6331 6307
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 6273 6267 6331 6273
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8220 6313 8248 6344
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 11698 6372 11704 6384
rect 9272 6344 11704 6372
rect 9272 6332 9278 6344
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 11974 6332 11980 6384
rect 12032 6372 12038 6384
rect 12544 6372 12572 6412
rect 12032 6344 12572 6372
rect 13740 6372 13768 6412
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 16942 6440 16948 6452
rect 15243 6412 16948 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 14093 6375 14151 6381
rect 14093 6372 14105 6375
rect 13740 6344 14105 6372
rect 12032 6332 12038 6344
rect 14093 6341 14105 6344
rect 14139 6341 14151 6375
rect 14093 6335 14151 6341
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 3605 6239 3663 6245
rect 3605 6236 3617 6239
rect 1443 6208 3617 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 3605 6205 3617 6208
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 3872 6239 3930 6245
rect 3872 6205 3884 6239
rect 3918 6236 3930 6239
rect 4706 6236 4712 6248
rect 3918 6208 4712 6236
rect 3918 6205 3930 6208
rect 3872 6199 3930 6205
rect 1664 6171 1722 6177
rect 1664 6137 1676 6171
rect 1710 6168 1722 6171
rect 2774 6168 2780 6180
rect 1710 6140 2780 6168
rect 1710 6137 1722 6140
rect 1664 6131 1722 6137
rect 2774 6128 2780 6140
rect 2832 6168 2838 6180
rect 2958 6168 2964 6180
rect 2832 6140 2964 6168
rect 2832 6128 2838 6140
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 3620 6168 3648 6199
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5684 6208 6009 6236
rect 5684 6196 5690 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 7190 6236 7196 6248
rect 7151 6208 7196 6236
rect 5997 6199 6055 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 5074 6168 5080 6180
rect 3620 6140 5080 6168
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 5644 6140 7297 6168
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 3053 6103 3111 6109
rect 3053 6100 3065 6103
rect 1912 6072 3065 6100
rect 1912 6060 1918 6072
rect 3053 6069 3065 6072
rect 3099 6069 3111 6103
rect 3053 6063 3111 6069
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4246 6100 4252 6112
rect 4120 6072 4252 6100
rect 4120 6060 4126 6072
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 5644 6109 5672 6140
rect 7285 6137 7297 6140
rect 7331 6137 7343 6171
rect 8220 6168 8248 6267
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 10410 6304 10416 6316
rect 9364 6276 10272 6304
rect 10371 6276 10416 6304
rect 9364 6264 9370 6276
rect 8478 6245 8484 6248
rect 8472 6236 8484 6245
rect 8391 6208 8484 6236
rect 8472 6199 8484 6208
rect 8536 6236 8542 6248
rect 10244 6245 10272 6276
rect 10410 6264 10416 6276
rect 10468 6264 10474 6316
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 11330 6304 11336 6316
rect 10836 6276 11336 6304
rect 10836 6264 10842 6276
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11606 6304 11612 6316
rect 11567 6276 11612 6304
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 12492 6276 12541 6304
rect 12492 6264 12498 6276
rect 12529 6273 12541 6276
rect 12575 6273 12587 6307
rect 12529 6267 12587 6273
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 14737 6307 14795 6313
rect 14737 6304 14749 6307
rect 13596 6276 14749 6304
rect 13596 6264 13602 6276
rect 14737 6273 14749 6276
rect 14783 6273 14795 6307
rect 15746 6304 15752 6316
rect 15707 6276 15752 6304
rect 14737 6267 14795 6273
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 10229 6239 10287 6245
rect 8536 6208 10171 6236
rect 8478 6196 8484 6199
rect 8536 6196 8542 6208
rect 8754 6168 8760 6180
rect 8220 6140 8760 6168
rect 7285 6131 7343 6137
rect 8754 6128 8760 6140
rect 8812 6168 8818 6180
rect 10042 6168 10048 6180
rect 8812 6140 10048 6168
rect 8812 6128 8818 6140
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 10143 6168 10171 6208
rect 10229 6205 10241 6239
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 11425 6239 11483 6245
rect 11425 6205 11437 6239
rect 11471 6236 11483 6239
rect 12618 6236 12624 6248
rect 11471 6208 12624 6236
rect 11471 6205 11483 6208
rect 11425 6199 11483 6205
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 14550 6236 14556 6248
rect 14511 6208 14556 6236
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 15654 6236 15660 6248
rect 15615 6208 15660 6236
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 15930 6196 15936 6248
rect 15988 6236 15994 6248
rect 16301 6239 16359 6245
rect 16301 6236 16313 6239
rect 15988 6208 16313 6236
rect 15988 6196 15994 6208
rect 16301 6205 16313 6208
rect 16347 6205 16359 6239
rect 16301 6199 16359 6205
rect 10410 6168 10416 6180
rect 10143 6140 10416 6168
rect 10410 6128 10416 6140
rect 10468 6128 10474 6180
rect 12796 6171 12854 6177
rect 11072 6140 11836 6168
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6069 5687 6103
rect 5629 6063 5687 6069
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 6089 6103 6147 6109
rect 6089 6100 6101 6103
rect 5776 6072 6101 6100
rect 5776 6060 5782 6072
rect 6089 6069 6101 6072
rect 6135 6069 6147 6103
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6089 6063 6147 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 9585 6103 9643 6109
rect 9585 6069 9597 6103
rect 9631 6100 9643 6103
rect 9674 6100 9680 6112
rect 9631 6072 9680 6100
rect 9631 6069 9643 6072
rect 9585 6063 9643 6069
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 9858 6100 9864 6112
rect 9819 6072 9864 6100
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 10321 6103 10379 6109
rect 10321 6069 10333 6103
rect 10367 6100 10379 6103
rect 10962 6100 10968 6112
rect 10367 6072 10968 6100
rect 10367 6069 10379 6072
rect 10321 6063 10379 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 11072 6109 11100 6140
rect 11057 6103 11115 6109
rect 11057 6069 11069 6103
rect 11103 6069 11115 6103
rect 11057 6063 11115 6069
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11388 6072 11529 6100
rect 11388 6060 11394 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11808 6100 11836 6140
rect 12796 6137 12808 6171
rect 12842 6168 12854 6171
rect 13538 6168 13544 6180
rect 12842 6140 13544 6168
rect 12842 6137 12854 6140
rect 12796 6131 12854 6137
rect 13538 6128 13544 6140
rect 13596 6128 13602 6180
rect 14093 6171 14151 6177
rect 14093 6137 14105 6171
rect 14139 6168 14151 6171
rect 14458 6168 14464 6180
rect 14139 6140 14464 6168
rect 14139 6137 14151 6140
rect 14093 6131 14151 6137
rect 14458 6128 14464 6140
rect 14516 6168 14522 6180
rect 14645 6171 14703 6177
rect 14645 6168 14657 6171
rect 14516 6140 14657 6168
rect 14516 6128 14522 6140
rect 14645 6137 14657 6140
rect 14691 6137 14703 6171
rect 14645 6131 14703 6137
rect 16568 6171 16626 6177
rect 16568 6137 16580 6171
rect 16614 6168 16626 6171
rect 17402 6168 17408 6180
rect 16614 6140 17408 6168
rect 16614 6137 16626 6140
rect 16568 6131 16626 6137
rect 17402 6128 17408 6140
rect 17460 6128 17466 6180
rect 13722 6100 13728 6112
rect 11808 6072 13728 6100
rect 11517 6063 11575 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 14185 6103 14243 6109
rect 14185 6069 14197 6103
rect 14231 6100 14243 6103
rect 14274 6100 14280 6112
rect 14231 6072 14280 6100
rect 14231 6069 14243 6072
rect 14185 6063 14243 6069
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 16022 6060 16028 6112
rect 16080 6100 16086 6112
rect 17681 6103 17739 6109
rect 17681 6100 17693 6103
rect 16080 6072 17693 6100
rect 16080 6060 16086 6072
rect 17681 6069 17693 6072
rect 17727 6069 17739 6103
rect 17681 6063 17739 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1486 5896 1492 5908
rect 1447 5868 1492 5896
rect 1486 5856 1492 5868
rect 1544 5856 1550 5908
rect 1854 5896 1860 5908
rect 1815 5868 1860 5896
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3476 5868 4077 5896
rect 3476 5856 3482 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4246 5856 4252 5908
rect 4304 5896 4310 5908
rect 8294 5896 8300 5908
rect 4304 5868 8300 5896
rect 4304 5856 4310 5868
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 9033 5899 9091 5905
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 9858 5896 9864 5908
rect 9079 5868 9864 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 13170 5896 13176 5908
rect 10336 5868 13176 5896
rect 5718 5828 5724 5840
rect 2884 5800 5724 5828
rect 2884 5772 2912 5800
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 6822 5788 6828 5840
rect 6880 5828 6886 5840
rect 6880 5800 9904 5828
rect 6880 5788 6886 5800
rect 9876 5772 9904 5800
rect 2866 5760 2872 5772
rect 2827 5732 2872 5760
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 3878 5720 3884 5772
rect 3936 5760 3942 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 3936 5732 4445 5760
rect 3936 5720 3942 5732
rect 4433 5729 4445 5732
rect 4479 5760 4491 5763
rect 4890 5760 4896 5772
rect 4479 5732 4896 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 5074 5720 5080 5772
rect 5132 5760 5138 5772
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 5132 5732 5549 5760
rect 5132 5720 5138 5732
rect 5537 5729 5549 5732
rect 5583 5760 5595 5763
rect 5626 5760 5632 5772
rect 5583 5732 5632 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 5810 5769 5816 5772
rect 5804 5723 5816 5769
rect 5868 5760 5874 5772
rect 7558 5760 7564 5772
rect 5868 5732 5904 5760
rect 7519 5732 7564 5760
rect 5810 5720 5816 5723
rect 5868 5720 5874 5732
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 8987 5732 9689 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 9858 5720 9864 5772
rect 9916 5720 9922 5772
rect 10336 5760 10364 5868
rect 13170 5856 13176 5868
rect 13228 5856 13234 5908
rect 13538 5896 13544 5908
rect 13499 5868 13544 5896
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14274 5896 14280 5908
rect 14235 5868 14280 5896
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 17402 5896 17408 5908
rect 17363 5868 17408 5896
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 10686 5788 10692 5840
rect 10744 5837 10750 5840
rect 10744 5831 10808 5837
rect 10744 5797 10762 5831
rect 10796 5797 10808 5831
rect 14182 5828 14188 5840
rect 14143 5800 14188 5828
rect 10744 5791 10808 5797
rect 10744 5788 10750 5791
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 16292 5831 16350 5837
rect 16292 5797 16304 5831
rect 16338 5828 16350 5831
rect 16482 5828 16488 5840
rect 16338 5800 16488 5828
rect 16338 5797 16350 5800
rect 16292 5791 16350 5797
rect 16482 5788 16488 5800
rect 16540 5788 16546 5840
rect 10413 5763 10471 5769
rect 10413 5760 10425 5763
rect 10336 5732 10425 5760
rect 10413 5729 10425 5732
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 10505 5763 10563 5769
rect 10505 5729 10517 5763
rect 10551 5760 10563 5763
rect 12069 5763 12127 5769
rect 10551 5732 11560 5760
rect 10551 5729 10563 5732
rect 10505 5723 10563 5729
rect 1578 5652 1584 5704
rect 1636 5692 1642 5704
rect 1949 5695 2007 5701
rect 1949 5692 1961 5695
rect 1636 5664 1961 5692
rect 1636 5652 1642 5664
rect 1949 5661 1961 5664
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2958 5692 2964 5704
rect 2179 5664 2636 5692
rect 2919 5664 2964 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2498 5556 2504 5568
rect 2459 5528 2504 5556
rect 2498 5516 2504 5528
rect 2556 5516 2562 5568
rect 2608 5556 2636 5664
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 3068 5624 3096 5655
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 3844 5664 4537 5692
rect 3844 5652 3850 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4525 5655 4583 5661
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7064 5664 7665 5692
rect 7064 5652 7070 5664
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 7834 5692 7840 5704
rect 7795 5664 7840 5692
rect 7653 5655 7711 5661
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8662 5692 8668 5704
rect 7935 5664 8668 5692
rect 2740 5596 3096 5624
rect 2740 5584 2746 5596
rect 6546 5584 6552 5636
rect 6604 5624 6610 5636
rect 7935 5624 7963 5664
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9766 5692 9772 5704
rect 9263 5664 9772 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 6604 5596 7963 5624
rect 8573 5627 8631 5633
rect 6604 5584 6610 5596
rect 8573 5593 8585 5627
rect 8619 5624 8631 5627
rect 9858 5624 9864 5636
rect 8619 5596 9864 5624
rect 8619 5593 8631 5596
rect 8573 5587 8631 5593
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10229 5627 10287 5633
rect 10229 5624 10241 5627
rect 10100 5596 10241 5624
rect 10100 5584 10106 5596
rect 10229 5593 10241 5596
rect 10275 5624 10287 5627
rect 10520 5624 10548 5723
rect 11532 5692 11560 5732
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 12428 5763 12486 5769
rect 12428 5760 12440 5763
rect 12115 5732 12440 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 12428 5729 12440 5732
rect 12474 5760 12486 5763
rect 12986 5760 12992 5772
rect 12474 5732 12992 5760
rect 12474 5729 12486 5732
rect 12428 5723 12486 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 15013 5763 15071 5769
rect 15013 5760 15025 5763
rect 13228 5732 15025 5760
rect 13228 5720 13234 5732
rect 15013 5729 15025 5732
rect 15059 5729 15071 5763
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 15013 5723 15071 5729
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 17678 5760 17684 5772
rect 17639 5732 17684 5760
rect 17678 5720 17684 5732
rect 17736 5720 17742 5772
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 11532 5664 12173 5692
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14369 5695 14427 5701
rect 14369 5692 14381 5695
rect 13964 5664 14381 5692
rect 13964 5652 13970 5664
rect 14369 5661 14381 5664
rect 14415 5661 14427 5695
rect 15470 5692 15476 5704
rect 15431 5664 15476 5692
rect 14369 5655 14427 5661
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 15930 5692 15936 5704
rect 15571 5664 15936 5692
rect 10275 5596 10548 5624
rect 11885 5627 11943 5633
rect 10275 5593 10287 5596
rect 10229 5587 10287 5593
rect 11885 5593 11897 5627
rect 11931 5624 11943 5627
rect 12069 5627 12127 5633
rect 12069 5624 12081 5627
rect 11931 5596 12081 5624
rect 11931 5593 11943 5596
rect 11885 5587 11943 5593
rect 12069 5593 12081 5596
rect 12115 5593 12127 5627
rect 12069 5587 12127 5593
rect 2774 5556 2780 5568
rect 2608 5528 2780 5556
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 6454 5556 6460 5568
rect 4120 5528 6460 5556
rect 4120 5516 4126 5528
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5556 6975 5559
rect 7098 5556 7104 5568
rect 6963 5528 7104 5556
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7193 5559 7251 5565
rect 7193 5525 7205 5559
rect 7239 5556 7251 5559
rect 8662 5556 8668 5568
rect 7239 5528 8668 5556
rect 7239 5525 7251 5528
rect 7193 5519 7251 5525
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 13814 5556 13820 5568
rect 13775 5528 13820 5556
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 14829 5559 14887 5565
rect 14829 5525 14841 5559
rect 14875 5556 14887 5559
rect 15010 5556 15016 5568
rect 14875 5528 15016 5556
rect 14875 5525 14887 5528
rect 14829 5519 14887 5525
rect 15010 5516 15016 5528
rect 15068 5556 15074 5568
rect 15571 5556 15599 5664
rect 15930 5652 15936 5664
rect 15988 5692 15994 5704
rect 16025 5695 16083 5701
rect 16025 5692 16037 5695
rect 15988 5664 16037 5692
rect 15988 5652 15994 5664
rect 16025 5661 16037 5664
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 15068 5528 15599 5556
rect 17865 5559 17923 5565
rect 15068 5516 15074 5528
rect 17865 5525 17877 5559
rect 17911 5556 17923 5559
rect 17954 5556 17960 5568
rect 17911 5528 17960 5556
rect 17911 5525 17923 5528
rect 17865 5519 17923 5525
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 3142 5312 3148 5364
rect 3200 5352 3206 5364
rect 5721 5355 5779 5361
rect 3200 5324 5304 5352
rect 3200 5312 3206 5324
rect 5276 5284 5304 5324
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 7006 5352 7012 5364
rect 5767 5324 7012 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 7892 5324 8217 5352
rect 7892 5312 7898 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 9784 5324 10548 5352
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 5276 5256 6561 5284
rect 6549 5253 6561 5256
rect 6595 5253 6607 5287
rect 6549 5247 6607 5253
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 2590 5216 2596 5228
rect 2455 5188 2596 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 2590 5176 2596 5188
rect 2648 5176 2654 5228
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 1854 5108 1860 5160
rect 1912 5148 1918 5160
rect 2682 5148 2688 5160
rect 1912 5120 2688 5148
rect 1912 5108 1918 5120
rect 2682 5108 2688 5120
rect 2740 5148 2746 5160
rect 3344 5148 3372 5179
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4396 5188 4813 5216
rect 4396 5176 4402 5188
rect 4801 5185 4813 5188
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5216 6423 5219
rect 8220 5216 8248 5315
rect 6411 5188 6960 5216
rect 8220 5188 8892 5216
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 2740 5120 3372 5148
rect 2740 5108 2746 5120
rect 3694 5108 3700 5160
rect 3752 5148 3758 5160
rect 4617 5151 4675 5157
rect 4617 5148 4629 5151
rect 3752 5120 4629 5148
rect 3752 5108 3758 5120
rect 4617 5117 4629 5120
rect 4663 5117 4675 5151
rect 4617 5111 4675 5117
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 6822 5148 6828 5160
rect 5684 5120 6828 5148
rect 5684 5108 5690 5120
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 1394 5040 1400 5092
rect 1452 5080 1458 5092
rect 2133 5083 2191 5089
rect 2133 5080 2145 5083
rect 1452 5052 2145 5080
rect 1452 5040 1458 5052
rect 2133 5049 2145 5052
rect 2179 5049 2191 5083
rect 2133 5043 2191 5049
rect 2406 5040 2412 5092
rect 2464 5080 2470 5092
rect 2958 5080 2964 5092
rect 2464 5052 2964 5080
rect 2464 5040 2470 5052
rect 2958 5040 2964 5052
rect 3016 5040 3022 5092
rect 6932 5080 6960 5188
rect 8754 5148 8760 5160
rect 8715 5120 8760 5148
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 8864 5148 8892 5188
rect 9013 5151 9071 5157
rect 9013 5148 9025 5151
rect 8864 5120 9025 5148
rect 9013 5117 9025 5120
rect 9059 5117 9071 5151
rect 9013 5111 9071 5117
rect 7098 5089 7104 5092
rect 7092 5080 7104 5089
rect 6932 5052 7104 5080
rect 7092 5043 7104 5052
rect 7098 5040 7104 5043
rect 7156 5040 7162 5092
rect 9784 5080 9812 5324
rect 10137 5287 10195 5293
rect 10137 5253 10149 5287
rect 10183 5253 10195 5287
rect 10137 5247 10195 5253
rect 10321 5287 10379 5293
rect 10321 5253 10333 5287
rect 10367 5284 10379 5287
rect 10413 5287 10471 5293
rect 10413 5284 10425 5287
rect 10367 5256 10425 5284
rect 10367 5253 10379 5256
rect 10321 5247 10379 5253
rect 10413 5253 10425 5256
rect 10459 5253 10471 5287
rect 10520 5284 10548 5324
rect 10520 5256 15700 5284
rect 10413 5247 10471 5253
rect 10152 5216 10180 5247
rect 10686 5216 10692 5228
rect 10152 5188 10692 5216
rect 10686 5176 10692 5188
rect 10744 5216 10750 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10744 5188 10977 5216
rect 10744 5176 10750 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 12986 5216 12992 5228
rect 12947 5188 12992 5216
rect 10965 5179 11023 5185
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 15672 5225 15700 5256
rect 15657 5219 15715 5225
rect 13780 5188 14412 5216
rect 13780 5176 13786 5188
rect 10321 5151 10379 5157
rect 10321 5117 10333 5151
rect 10367 5148 10379 5151
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 10367 5120 12909 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 13633 5151 13691 5157
rect 13633 5117 13645 5151
rect 13679 5148 13691 5151
rect 13814 5148 13820 5160
rect 13679 5120 13820 5148
rect 13679 5117 13691 5120
rect 13633 5111 13691 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14384 5157 14412 5188
rect 15657 5185 15669 5219
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5216 15899 5219
rect 16482 5216 16488 5228
rect 15887 5188 16488 5216
rect 15887 5185 15899 5188
rect 15841 5179 15899 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5216 16911 5219
rect 17402 5216 17408 5228
rect 16899 5188 17408 5216
rect 16899 5185 16911 5188
rect 16853 5179 16911 5185
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 14369 5151 14427 5157
rect 14369 5117 14381 5151
rect 14415 5117 14427 5151
rect 14369 5111 14427 5117
rect 15565 5151 15623 5157
rect 15565 5117 15577 5151
rect 15611 5148 15623 5151
rect 17221 5151 17279 5157
rect 17221 5148 17233 5151
rect 15611 5120 17233 5148
rect 15611 5117 15623 5120
rect 15565 5111 15623 5117
rect 17221 5117 17233 5120
rect 17267 5117 17279 5151
rect 17221 5111 17279 5117
rect 7208 5052 9812 5080
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 2222 5012 2228 5024
rect 2183 4984 2228 5012
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 2372 4984 2789 5012
rect 2372 4972 2378 4984
rect 2777 4981 2789 4984
rect 2823 4981 2835 5015
rect 3142 5012 3148 5024
rect 3103 4984 3148 5012
rect 2777 4975 2835 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 3237 5015 3295 5021
rect 3237 4981 3249 5015
rect 3283 5012 3295 5015
rect 3326 5012 3332 5024
rect 3283 4984 3332 5012
rect 3283 4981 3295 4984
rect 3237 4975 3295 4981
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 4246 5012 4252 5024
rect 4207 4984 4252 5012
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 6086 5012 6092 5024
rect 6047 4984 6092 5012
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6178 4972 6184 5024
rect 6236 5012 6242 5024
rect 6549 5015 6607 5021
rect 6236 4984 6281 5012
rect 6236 4972 6242 4984
rect 6549 4981 6561 5015
rect 6595 5012 6607 5015
rect 7208 5012 7236 5052
rect 10594 5040 10600 5092
rect 10652 5080 10658 5092
rect 10873 5083 10931 5089
rect 10873 5080 10885 5083
rect 10652 5052 10885 5080
rect 10652 5040 10658 5052
rect 10873 5049 10885 5052
rect 10919 5049 10931 5083
rect 10873 5043 10931 5049
rect 11885 5083 11943 5089
rect 11885 5049 11897 5083
rect 11931 5080 11943 5083
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 11931 5052 12817 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 12805 5043 12863 5049
rect 13909 5083 13967 5089
rect 13909 5049 13921 5083
rect 13955 5080 13967 5083
rect 14274 5080 14280 5092
rect 13955 5052 14280 5080
rect 13955 5049 13967 5052
rect 13909 5043 13967 5049
rect 14274 5040 14280 5052
rect 14332 5040 14338 5092
rect 14550 5040 14556 5092
rect 14608 5080 14614 5092
rect 14645 5083 14703 5089
rect 14645 5080 14657 5083
rect 14608 5052 14657 5080
rect 14608 5040 14614 5052
rect 14645 5049 14657 5052
rect 14691 5049 14703 5083
rect 16577 5083 16635 5089
rect 16577 5080 16589 5083
rect 14645 5043 14703 5049
rect 15212 5052 16589 5080
rect 6595 4984 7236 5012
rect 6595 4981 6607 4984
rect 6549 4975 6607 4981
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 10781 5015 10839 5021
rect 10781 5012 10793 5015
rect 8352 4984 10793 5012
rect 8352 4972 8358 4984
rect 10781 4981 10793 4984
rect 10827 4981 10839 5015
rect 10781 4975 10839 4981
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 12618 5012 12624 5024
rect 12483 4984 12624 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 15212 5021 15240 5052
rect 16577 5049 16589 5052
rect 16623 5049 16635 5083
rect 16577 5043 16635 5049
rect 15197 5015 15255 5021
rect 15197 4981 15209 5015
rect 15243 4981 15255 5015
rect 16206 5012 16212 5024
rect 16167 4984 16212 5012
rect 15197 4975 15255 4981
rect 16206 4972 16212 4984
rect 16264 4972 16270 5024
rect 16666 4972 16672 5024
rect 16724 5012 16730 5024
rect 16724 4984 16769 5012
rect 16724 4972 16730 4984
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1394 4808 1400 4820
rect 1355 4780 1400 4808
rect 1394 4768 1400 4780
rect 1452 4768 1458 4820
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4985 4811 5043 4817
rect 4985 4808 4997 4811
rect 4304 4780 4997 4808
rect 4304 4768 4310 4780
rect 4985 4777 4997 4780
rect 5031 4777 5043 4811
rect 4985 4771 5043 4777
rect 5537 4811 5595 4817
rect 5537 4777 5549 4811
rect 5583 4808 5595 4811
rect 6178 4808 6184 4820
rect 5583 4780 6184 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 6549 4811 6607 4817
rect 6549 4777 6561 4811
rect 6595 4808 6607 4811
rect 7558 4808 7564 4820
rect 6595 4780 7564 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 14185 4811 14243 4817
rect 14185 4808 14197 4811
rect 9640 4780 14197 4808
rect 9640 4768 9646 4780
rect 14185 4777 14197 4780
rect 14231 4777 14243 4811
rect 14185 4771 14243 4777
rect 2406 4700 2412 4752
rect 2464 4740 2470 4752
rect 2464 4712 3924 4740
rect 2464 4700 2470 4712
rect 2124 4675 2182 4681
rect 2124 4641 2136 4675
rect 2170 4672 2182 4675
rect 2590 4672 2596 4684
rect 2170 4644 2596 4672
rect 2170 4641 2182 4644
rect 2124 4635 2182 4641
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4573 1915 4607
rect 1857 4567 1915 4573
rect 1872 4468 1900 4567
rect 3896 4536 3924 4712
rect 4062 4700 4068 4752
rect 4120 4740 4126 4752
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 4120 4712 8217 4740
rect 4120 4700 4126 4712
rect 8205 4709 8217 4712
rect 8251 4709 8263 4743
rect 8205 4703 8263 4709
rect 8662 4700 8668 4752
rect 8720 4740 8726 4752
rect 9401 4743 9459 4749
rect 9401 4740 9413 4743
rect 8720 4712 9413 4740
rect 8720 4700 8726 4712
rect 9401 4709 9413 4712
rect 9447 4709 9459 4743
rect 9401 4703 9459 4709
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 9922 4743 9980 4749
rect 9922 4740 9934 4743
rect 9824 4712 9934 4740
rect 9824 4700 9830 4712
rect 9922 4709 9934 4712
rect 9968 4709 9980 4743
rect 18316 4743 18374 4749
rect 9922 4703 9980 4709
rect 15488 4712 18092 4740
rect 4890 4672 4896 4684
rect 4851 4644 4896 4672
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 5905 4675 5963 4681
rect 5905 4672 5917 4675
rect 5776 4644 5917 4672
rect 5776 4632 5782 4644
rect 5905 4641 5917 4644
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6546 4672 6552 4684
rect 6043 4644 6552 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 6012 4604 6040 4635
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 6914 4672 6920 4684
rect 6875 4644 6920 4672
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4672 9643 4675
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 9631 4644 12449 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 12437 4635 12495 4641
rect 12544 4644 14105 4672
rect 5184 4576 6040 4604
rect 6089 4607 6147 4613
rect 5184 4536 5212 4576
rect 6089 4573 6101 4607
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 3896 4508 5212 4536
rect 5810 4496 5816 4548
rect 5868 4536 5874 4548
rect 6104 4536 6132 4567
rect 6454 4564 6460 4616
rect 6512 4604 6518 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6512 4576 7021 4604
rect 6512 4564 6518 4576
rect 7009 4573 7021 4576
rect 7055 4573 7067 4607
rect 7190 4604 7196 4616
rect 7151 4576 7196 4604
rect 7009 4567 7067 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 8294 4604 8300 4616
rect 8255 4576 8300 4604
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 5868 4508 6132 4536
rect 5868 4496 5874 4508
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 8404 4536 8432 4567
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9490 4604 9496 4616
rect 8812 4576 9496 4604
rect 8812 4564 8818 4576
rect 9490 4564 9496 4576
rect 9548 4604 9554 4616
rect 9677 4607 9735 4613
rect 9677 4604 9689 4607
rect 9548 4576 9689 4604
rect 9548 4564 9554 4576
rect 9677 4573 9689 4576
rect 9723 4573 9735 4607
rect 9677 4567 9735 4573
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 10836 4576 11345 4604
rect 10836 4564 10842 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 12544 4604 12572 4644
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 11664 4576 12572 4604
rect 12713 4607 12771 4613
rect 11664 4564 11670 4576
rect 12713 4573 12725 4607
rect 12759 4604 12771 4607
rect 13630 4604 13636 4616
rect 12759 4576 13636 4604
rect 12759 4573 12771 4576
rect 12713 4567 12771 4573
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4604 14427 4607
rect 14734 4604 14740 4616
rect 14415 4576 14740 4604
rect 14415 4573 14427 4576
rect 14369 4567 14427 4573
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 15488 4613 15516 4712
rect 15740 4675 15798 4681
rect 15740 4641 15752 4675
rect 15786 4672 15798 4675
rect 16114 4672 16120 4684
rect 15786 4644 16120 4672
rect 15786 4641 15798 4644
rect 15740 4635 15798 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 16206 4632 16212 4684
rect 16264 4672 16270 4684
rect 18064 4681 18092 4712
rect 18316 4709 18328 4743
rect 18362 4740 18374 4743
rect 18598 4740 18604 4752
rect 18362 4712 18604 4740
rect 18362 4709 18374 4712
rect 18316 4703 18374 4709
rect 18598 4700 18604 4712
rect 18656 4700 18662 4752
rect 17129 4675 17187 4681
rect 17129 4672 17141 4675
rect 16264 4644 17141 4672
rect 16264 4632 16270 4644
rect 17129 4641 17141 4644
rect 17175 4641 17187 4675
rect 17129 4635 17187 4641
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4641 18107 4675
rect 18049 4635 18107 4641
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 15068 4576 15485 4604
rect 15068 4564 15074 4576
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 17276 4576 17325 4604
rect 17276 4564 17282 4576
rect 17313 4573 17325 4576
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 7800 4508 8432 4536
rect 7800 4496 7806 4508
rect 10686 4496 10692 4548
rect 10744 4536 10750 4548
rect 13725 4539 13783 4545
rect 10744 4508 11183 4536
rect 10744 4496 10750 4508
rect 2222 4468 2228 4480
rect 1872 4440 2228 4468
rect 2222 4428 2228 4440
rect 2280 4428 2286 4480
rect 3234 4468 3240 4480
rect 3195 4440 3240 4468
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 4525 4471 4583 4477
rect 4525 4437 4537 4471
rect 4571 4468 4583 4471
rect 5350 4468 5356 4480
rect 4571 4440 5356 4468
rect 4571 4437 4583 4440
rect 4525 4431 4583 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 7834 4468 7840 4480
rect 7795 4440 7840 4468
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 10042 4428 10048 4480
rect 10100 4468 10106 4480
rect 11057 4471 11115 4477
rect 11057 4468 11069 4471
rect 10100 4440 11069 4468
rect 10100 4428 10106 4440
rect 11057 4437 11069 4440
rect 11103 4437 11115 4471
rect 11155 4468 11183 4508
rect 13725 4505 13737 4539
rect 13771 4536 13783 4539
rect 15102 4536 15108 4548
rect 13771 4508 15108 4536
rect 13771 4505 13783 4508
rect 13725 4499 13783 4505
rect 15102 4496 15108 4508
rect 15160 4496 15166 4548
rect 16408 4508 16988 4536
rect 16408 4468 16436 4508
rect 11155 4440 16436 4468
rect 11057 4431 11115 4437
rect 16482 4428 16488 4480
rect 16540 4468 16546 4480
rect 16850 4468 16856 4480
rect 16540 4440 16856 4468
rect 16540 4428 16546 4440
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 16960 4468 16988 4508
rect 19429 4471 19487 4477
rect 19429 4468 19441 4471
rect 16960 4440 19441 4468
rect 19429 4437 19441 4440
rect 19475 4437 19487 4471
rect 19429 4431 19487 4437
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 5718 4264 5724 4276
rect 5092 4236 5724 4264
rect 4338 4156 4344 4208
rect 4396 4196 4402 4208
rect 4890 4196 4896 4208
rect 4396 4168 4896 4196
rect 4396 4156 4402 4168
rect 4890 4156 4896 4168
rect 4948 4156 4954 4208
rect 198 4088 204 4140
rect 256 4128 262 4140
rect 2406 4128 2412 4140
rect 256 4100 2412 4128
rect 256 4088 262 4100
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2639 4100 3096 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 1762 4020 1768 4072
rect 1820 4060 1826 4072
rect 2317 4063 2375 4069
rect 2317 4060 2329 4063
rect 1820 4032 2329 4060
rect 1820 4020 1826 4032
rect 2317 4029 2329 4032
rect 2363 4029 2375 4063
rect 2317 4023 2375 4029
rect 2774 4020 2780 4072
rect 2832 4060 2838 4072
rect 2961 4063 3019 4069
rect 2961 4060 2973 4063
rect 2832 4032 2973 4060
rect 2832 4020 2838 4032
rect 2961 4029 2973 4032
rect 3007 4029 3019 4063
rect 3068 4060 3096 4100
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4982 4128 4988 4140
rect 4120 4100 4988 4128
rect 4120 4088 4126 4100
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 3234 4069 3240 4072
rect 3228 4060 3240 4069
rect 3068 4032 3240 4060
rect 2961 4023 3019 4029
rect 3228 4023 3240 4032
rect 3234 4020 3240 4023
rect 3292 4020 3298 4072
rect 4522 4020 4528 4072
rect 4580 4060 4586 4072
rect 5092 4069 5120 4236
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 6454 4264 6460 4276
rect 5868 4236 6460 4264
rect 5868 4224 5874 4236
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 11606 4264 11612 4276
rect 8904 4236 11612 4264
rect 8904 4224 8910 4236
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 14734 4264 14740 4276
rect 14695 4236 14740 4264
rect 14734 4224 14740 4236
rect 14792 4224 14798 4276
rect 16114 4224 16120 4276
rect 16172 4264 16178 4276
rect 16393 4267 16451 4273
rect 16393 4264 16405 4267
rect 16172 4236 16405 4264
rect 16172 4224 16178 4236
rect 16393 4233 16405 4236
rect 16439 4233 16451 4267
rect 16666 4264 16672 4276
rect 16627 4236 16672 4264
rect 16393 4227 16451 4233
rect 16666 4224 16672 4236
rect 16724 4224 16730 4276
rect 8573 4199 8631 4205
rect 8573 4165 8585 4199
rect 8619 4196 8631 4199
rect 9585 4199 9643 4205
rect 9585 4196 9597 4199
rect 8619 4168 9597 4196
rect 8619 4165 8631 4168
rect 8573 4159 8631 4165
rect 9585 4165 9597 4168
rect 9631 4165 9643 4199
rect 9585 4159 9643 4165
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4128 6883 4131
rect 6914 4128 6920 4140
rect 6871 4100 6920 4128
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7650 4128 7656 4140
rect 7524 4100 7656 4128
rect 7524 4088 7530 4100
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 7892 4100 8217 4128
rect 7892 4088 7898 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 9401 4131 9459 4137
rect 8352 4100 8397 4128
rect 8352 4088 8358 4100
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 14752 4128 14780 4224
rect 16850 4156 16856 4208
rect 16908 4196 16914 4208
rect 16908 4168 17264 4196
rect 16908 4156 16914 4168
rect 17236 4137 17264 4168
rect 17221 4131 17279 4137
rect 9447 4100 9904 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 5077 4063 5135 4069
rect 5077 4060 5089 4063
rect 4580 4032 5089 4060
rect 4580 4020 4586 4032
rect 5077 4029 5089 4032
rect 5123 4029 5135 4063
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 5077 4023 5135 4029
rect 5276 4032 8585 4060
rect 5276 3992 5304 4032
rect 8573 4029 8585 4032
rect 8619 4029 8631 4063
rect 8573 4023 8631 4029
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 8720 4032 9229 4060
rect 8720 4020 8726 4032
rect 9217 4029 9229 4032
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 9548 4032 9781 4060
rect 9548 4020 9554 4032
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 9876 4060 9904 4100
rect 11532 4100 13492 4128
rect 14752 4100 15148 4128
rect 10042 4069 10048 4072
rect 10036 4060 10048 4069
rect 9876 4032 10048 4060
rect 9769 4023 9827 4029
rect 10036 4023 10048 4032
rect 10042 4020 10048 4023
rect 10100 4020 10106 4072
rect 11425 4063 11483 4069
rect 11425 4060 11437 4063
rect 10520 4032 11437 4060
rect 1964 3964 5304 3992
rect 5344 3995 5402 4001
rect 1964 3933 1992 3964
rect 5344 3961 5356 3995
rect 5390 3992 5402 3995
rect 5442 3992 5448 4004
rect 5390 3964 5448 3992
rect 5390 3961 5402 3964
rect 5344 3955 5402 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 8386 3992 8392 4004
rect 7760 3964 8392 3992
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3893 2007 3927
rect 1949 3887 2007 3893
rect 2038 3884 2044 3936
rect 2096 3924 2102 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 2096 3896 2421 3924
rect 2096 3884 2102 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2409 3887 2467 3893
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4341 3927 4399 3933
rect 4341 3924 4353 3927
rect 4304 3896 4353 3924
rect 4304 3884 4310 3896
rect 4341 3893 4353 3896
rect 4387 3893 4399 3927
rect 4341 3887 4399 3893
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 7282 3924 7288 3936
rect 5040 3896 7288 3924
rect 5040 3884 5046 3896
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 7760 3933 7788 3964
rect 8386 3952 8392 3964
rect 8444 3952 8450 4004
rect 9585 3995 9643 4001
rect 9585 3961 9597 3995
rect 9631 3992 9643 3995
rect 10520 3992 10548 4032
rect 11425 4029 11437 4032
rect 11471 4029 11483 4063
rect 11425 4023 11483 4029
rect 11532 3992 11560 4100
rect 11606 4020 11612 4072
rect 11664 4060 11670 4072
rect 12066 4060 12072 4072
rect 11664 4032 12072 4060
rect 11664 4020 11670 4032
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 12618 4060 12624 4072
rect 12579 4032 12624 4060
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 13354 4060 13360 4072
rect 13267 4032 13360 4060
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 13464 4060 13492 4100
rect 15010 4060 15016 4072
rect 13464 4032 14044 4060
rect 14971 4032 15016 4060
rect 9631 3964 10548 3992
rect 10980 3964 11560 3992
rect 11701 3995 11759 4001
rect 9631 3961 9643 3964
rect 9585 3955 9643 3961
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3893 7803 3927
rect 7745 3887 7803 3893
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8570 3924 8576 3936
rect 8159 3896 8576 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8754 3924 8760 3936
rect 8715 3896 8760 3924
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 9122 3924 9128 3936
rect 9083 3896 9128 3924
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 10980 3924 11008 3964
rect 11701 3961 11713 3995
rect 11747 3992 11759 3995
rect 12526 3992 12532 4004
rect 11747 3964 12532 3992
rect 11747 3961 11759 3964
rect 11701 3955 11759 3961
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 12894 3992 12900 4004
rect 12855 3964 12900 3992
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 11146 3924 11152 3936
rect 9272 3896 11008 3924
rect 11107 3896 11152 3924
rect 9272 3884 9278 3896
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13363 3924 13391 4020
rect 13624 3995 13682 4001
rect 13624 3961 13636 3995
rect 13670 3992 13682 3995
rect 13906 3992 13912 4004
rect 13670 3964 13912 3992
rect 13670 3961 13682 3964
rect 13624 3955 13682 3961
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 14016 3992 14044 4032
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 15120 4060 15148 4100
rect 17221 4097 17233 4131
rect 17267 4097 17279 4131
rect 17221 4091 17279 4097
rect 15269 4063 15327 4069
rect 15269 4060 15281 4063
rect 15120 4032 15281 4060
rect 15269 4029 15281 4032
rect 15315 4029 15327 4063
rect 15269 4023 15327 4029
rect 17037 3995 17095 4001
rect 17037 3992 17049 3995
rect 14016 3964 17049 3992
rect 17037 3961 17049 3964
rect 17083 3961 17095 3995
rect 17037 3955 17095 3961
rect 12492 3896 13391 3924
rect 12492 3884 12498 3896
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 17129 3927 17187 3933
rect 17129 3924 17141 3927
rect 13596 3896 17141 3924
rect 13596 3884 13602 3896
rect 17129 3893 17141 3896
rect 17175 3924 17187 3927
rect 21174 3924 21180 3936
rect 17175 3896 21180 3924
rect 17175 3893 17187 3896
rect 17129 3887 17187 3893
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2004 3692 2912 3720
rect 2004 3680 2010 3692
rect 1670 3652 1676 3664
rect 1583 3624 1676 3652
rect 1596 3593 1624 3624
rect 1670 3612 1676 3624
rect 1728 3652 1734 3664
rect 2774 3652 2780 3664
rect 1728 3624 2780 3652
rect 1728 3612 1734 3624
rect 2774 3612 2780 3624
rect 2832 3612 2838 3664
rect 1854 3593 1860 3596
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3553 1639 3587
rect 1848 3584 1860 3593
rect 1815 3556 1860 3584
rect 1581 3547 1639 3553
rect 1848 3547 1860 3556
rect 1854 3544 1860 3547
rect 1912 3544 1918 3596
rect 2884 3584 2912 3692
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 13906 3720 13912 3732
rect 3016 3692 13768 3720
rect 13867 3692 13912 3720
rect 3016 3680 3022 3692
rect 4065 3655 4123 3661
rect 4065 3621 4077 3655
rect 4111 3652 4123 3655
rect 4338 3652 4344 3664
rect 4111 3624 4344 3652
rect 4111 3621 4123 3624
rect 4065 3615 4123 3621
rect 4338 3612 4344 3624
rect 4396 3612 4402 3664
rect 6825 3655 6883 3661
rect 6825 3652 6837 3655
rect 4448 3624 6837 3652
rect 3326 3584 3332 3596
rect 2884 3556 3332 3584
rect 3326 3544 3332 3556
rect 3384 3584 3390 3596
rect 4448 3584 4476 3624
rect 6825 3621 6837 3624
rect 6871 3652 6883 3655
rect 8662 3652 8668 3664
rect 6871 3624 8668 3652
rect 6871 3621 6883 3624
rect 6825 3615 6883 3621
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 10321 3655 10379 3661
rect 10321 3652 10333 3655
rect 8812 3624 10333 3652
rect 8812 3612 8818 3624
rect 10321 3621 10333 3624
rect 10367 3621 10379 3655
rect 10321 3615 10379 3621
rect 10410 3612 10416 3664
rect 10468 3652 10474 3664
rect 11146 3661 11152 3664
rect 11140 3652 11152 3661
rect 10468 3624 11152 3652
rect 10468 3612 10474 3624
rect 11140 3615 11152 3624
rect 11146 3612 11152 3615
rect 11204 3612 11210 3664
rect 3384 3556 4476 3584
rect 4792 3587 4850 3593
rect 3384 3544 3390 3556
rect 4792 3553 4804 3587
rect 4838 3584 4850 3587
rect 5074 3584 5080 3596
rect 4838 3556 5080 3584
rect 4838 3553 4850 3556
rect 4792 3547 4850 3553
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 6730 3584 6736 3596
rect 6691 3556 6736 3584
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 6840 3556 7696 3584
rect 6840 3528 6868 3556
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 4522 3516 4528 3528
rect 3936 3488 4528 3516
rect 3936 3476 3942 3488
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3485 6975 3519
rect 7668 3516 7696 3556
rect 7834 3544 7840 3596
rect 7892 3584 7898 3596
rect 8012 3587 8070 3593
rect 8012 3584 8024 3587
rect 7892 3556 8024 3584
rect 7892 3544 7898 3556
rect 8012 3553 8024 3556
rect 8058 3584 8070 3587
rect 10134 3584 10140 3596
rect 8058 3556 10140 3584
rect 8058 3553 8070 3556
rect 8012 3547 8070 3553
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10229 3587 10287 3593
rect 10229 3553 10241 3587
rect 10275 3553 10287 3587
rect 10229 3547 10287 3553
rect 7745 3519 7803 3525
rect 7745 3516 7757 3519
rect 7668 3488 7757 3516
rect 6917 3479 6975 3485
rect 7745 3485 7757 3488
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 2866 3448 2872 3460
rect 2516 3420 2872 3448
rect 1026 3340 1032 3392
rect 1084 3380 1090 3392
rect 2516 3380 2544 3420
rect 2866 3408 2872 3420
rect 2924 3408 2930 3460
rect 5460 3420 6040 3448
rect 1084 3352 2544 3380
rect 1084 3340 1090 3352
rect 2590 3340 2596 3392
rect 2648 3380 2654 3392
rect 2961 3383 3019 3389
rect 2961 3380 2973 3383
rect 2648 3352 2973 3380
rect 2648 3340 2654 3352
rect 2961 3349 2973 3352
rect 3007 3349 3019 3383
rect 2961 3343 3019 3349
rect 3326 3340 3332 3392
rect 3384 3380 3390 3392
rect 5460 3380 5488 3420
rect 3384 3352 5488 3380
rect 3384 3340 3390 3352
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 5905 3383 5963 3389
rect 5905 3380 5917 3383
rect 5868 3352 5917 3380
rect 5868 3340 5874 3352
rect 5905 3349 5917 3352
rect 5951 3349 5963 3383
rect 6012 3380 6040 3420
rect 6086 3408 6092 3460
rect 6144 3448 6150 3460
rect 6365 3451 6423 3457
rect 6365 3448 6377 3451
rect 6144 3420 6377 3448
rect 6144 3408 6150 3420
rect 6365 3417 6377 3420
rect 6411 3417 6423 3451
rect 6365 3411 6423 3417
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 6932 3448 6960 3479
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 9548 3488 10180 3516
rect 9548 3476 9554 3488
rect 6512 3420 6960 3448
rect 6512 3408 6518 3420
rect 8018 3380 8024 3392
rect 6012 3352 8024 3380
rect 5905 3343 5963 3349
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 9125 3383 9183 3389
rect 9125 3380 9137 3383
rect 8168 3352 9137 3380
rect 8168 3340 8174 3352
rect 9125 3349 9137 3352
rect 9171 3349 9183 3383
rect 9858 3380 9864 3392
rect 9819 3352 9864 3380
rect 9125 3343 9183 3349
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 10152 3380 10180 3488
rect 10244 3448 10272 3547
rect 10594 3544 10600 3596
rect 10652 3584 10658 3596
rect 10652 3556 12204 3584
rect 10652 3544 10658 3556
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 10689 3519 10747 3525
rect 10468 3488 10513 3516
rect 10468 3476 10474 3488
rect 10689 3485 10701 3519
rect 10735 3516 10747 3519
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10735 3488 10885 3516
rect 10735 3485 10747 3488
rect 10689 3479 10747 3485
rect 10873 3485 10885 3488
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 10778 3448 10784 3460
rect 10244 3420 10784 3448
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 12176 3448 12204 3556
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12785 3587 12843 3593
rect 12785 3584 12797 3587
rect 12308 3556 12797 3584
rect 12308 3544 12314 3556
rect 12785 3553 12797 3556
rect 12831 3553 12843 3587
rect 12785 3547 12843 3553
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 12492 3488 12541 3516
rect 12492 3476 12498 3488
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 12176 3420 12388 3448
rect 10689 3383 10747 3389
rect 10689 3380 10701 3383
rect 10152 3352 10701 3380
rect 10689 3349 10701 3352
rect 10735 3349 10747 3383
rect 12250 3380 12256 3392
rect 12211 3352 12256 3380
rect 10689 3343 10747 3349
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 12360 3380 12388 3420
rect 13538 3380 13544 3392
rect 12360 3352 13544 3380
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 13740 3380 13768 3692
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 15841 3723 15899 3729
rect 15841 3689 15853 3723
rect 15887 3720 15899 3723
rect 18325 3723 18383 3729
rect 18325 3720 18337 3723
rect 15887 3692 18337 3720
rect 15887 3689 15899 3692
rect 15841 3683 15899 3689
rect 18325 3689 18337 3692
rect 18371 3689 18383 3723
rect 18325 3683 18383 3689
rect 14366 3584 14372 3596
rect 14327 3556 14372 3584
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 15933 3587 15991 3593
rect 15933 3584 15945 3587
rect 15160 3556 15945 3584
rect 15160 3544 15166 3556
rect 15933 3553 15945 3556
rect 15979 3553 15991 3587
rect 15933 3547 15991 3553
rect 16485 3587 16543 3593
rect 16485 3553 16497 3587
rect 16531 3553 16543 3587
rect 17218 3584 17224 3596
rect 17179 3556 17224 3584
rect 16485 3547 16543 3553
rect 14645 3519 14703 3525
rect 14645 3485 14657 3519
rect 14691 3516 14703 3519
rect 15838 3516 15844 3528
rect 14691 3488 15844 3516
rect 14691 3485 14703 3488
rect 14645 3479 14703 3485
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 16114 3516 16120 3528
rect 16075 3488 16120 3516
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 15473 3451 15531 3457
rect 15473 3417 15485 3451
rect 15519 3448 15531 3451
rect 16500 3448 16528 3547
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 17770 3584 17776 3596
rect 17731 3556 17776 3584
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 19981 3587 20039 3593
rect 19981 3553 19993 3587
rect 20027 3553 20039 3587
rect 19981 3547 20039 3553
rect 16666 3516 16672 3528
rect 16627 3488 16672 3516
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 19996 3448 20024 3547
rect 15519 3420 16528 3448
rect 16592 3420 20024 3448
rect 15519 3417 15531 3420
rect 15473 3411 15531 3417
rect 16592 3380 16620 3420
rect 13740 3352 16620 3380
rect 17405 3383 17463 3389
rect 17405 3349 17417 3383
rect 17451 3380 17463 3383
rect 17678 3380 17684 3392
rect 17451 3352 17684 3380
rect 17451 3349 17463 3352
rect 17405 3343 17463 3349
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 17957 3383 18015 3389
rect 17957 3349 17969 3383
rect 18003 3380 18015 3383
rect 18598 3380 18604 3392
rect 18003 3352 18604 3380
rect 18003 3349 18015 3352
rect 17957 3343 18015 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 20165 3383 20223 3389
rect 20165 3349 20177 3383
rect 20211 3380 20223 3383
rect 20806 3380 20812 3392
rect 20211 3352 20812 3380
rect 20211 3349 20223 3352
rect 20165 3343 20223 3349
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 3513 3179 3571 3185
rect 3513 3176 3525 3179
rect 1912 3148 3525 3176
rect 1912 3136 1918 3148
rect 3513 3145 3525 3148
rect 3559 3145 3571 3179
rect 3513 3139 3571 3145
rect 3712 3148 5028 3176
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2972 2191 2975
rect 2222 2972 2228 2984
rect 2179 2944 2228 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 2400 2975 2458 2981
rect 2400 2941 2412 2975
rect 2446 2972 2458 2975
rect 3712 2972 3740 3148
rect 5000 3108 5028 3148
rect 5074 3136 5080 3188
rect 5132 3176 5138 3188
rect 5258 3176 5264 3188
rect 5132 3148 5264 3176
rect 5132 3136 5138 3148
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 5718 3176 5724 3188
rect 5679 3148 5724 3176
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 6086 3136 6092 3188
rect 6144 3176 6150 3188
rect 9214 3176 9220 3188
rect 6144 3148 9220 3176
rect 6144 3136 6150 3148
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 9916 3148 15056 3176
rect 9916 3136 9922 3148
rect 5000 3080 6684 3108
rect 3878 3040 3884 3052
rect 3839 3012 3884 3040
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 5810 3040 5816 3052
rect 5500 3012 5816 3040
rect 5500 3000 5506 3012
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 6273 3043 6331 3049
rect 6273 3009 6285 3043
rect 6319 3009 6331 3043
rect 6656 3040 6684 3080
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 11333 3111 11391 3117
rect 8352 3080 9628 3108
rect 8352 3068 8358 3080
rect 9493 3043 9551 3049
rect 6656 3012 7420 3040
rect 6273 3003 6331 3009
rect 2446 2944 3740 2972
rect 4148 2975 4206 2981
rect 2446 2941 2458 2944
rect 2400 2935 2458 2941
rect 4148 2941 4160 2975
rect 4194 2972 4206 2975
rect 6288 2972 6316 3003
rect 4194 2944 6316 2972
rect 4194 2941 4206 2944
rect 4148 2935 4206 2941
rect 4264 2916 4292 2944
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 6880 2944 7297 2972
rect 6880 2932 6886 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7392 2972 7420 3012
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 7552 2975 7610 2981
rect 7392 2944 7512 2972
rect 7285 2935 7343 2941
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 624 2876 4200 2904
rect 624 2864 630 2876
rect 1486 2796 1492 2848
rect 1544 2836 1550 2848
rect 3418 2836 3424 2848
rect 1544 2808 3424 2836
rect 1544 2796 1550 2808
rect 3418 2796 3424 2808
rect 3476 2796 3482 2848
rect 4172 2836 4200 2876
rect 4246 2864 4252 2916
rect 4304 2864 4310 2916
rect 5718 2864 5724 2916
rect 5776 2904 5782 2916
rect 7374 2904 7380 2916
rect 5776 2876 7380 2904
rect 5776 2864 5782 2876
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 6086 2836 6092 2848
rect 4172 2808 6092 2836
rect 6086 2796 6092 2808
rect 6144 2796 6150 2848
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 7006 2836 7012 2848
rect 6227 2808 7012 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 7484 2836 7512 2944
rect 7552 2941 7564 2975
rect 7598 2972 7610 2975
rect 7926 2972 7932 2984
rect 7598 2944 7932 2972
rect 7598 2941 7610 2944
rect 7552 2935 7610 2941
rect 7926 2932 7932 2944
rect 7984 2972 7990 2984
rect 9508 2972 9536 3003
rect 7984 2944 9536 2972
rect 9600 2972 9628 3080
rect 11333 3077 11345 3111
rect 11379 3108 11391 3111
rect 13357 3111 13415 3117
rect 13357 3108 13369 3111
rect 11379 3080 13369 3108
rect 11379 3077 11391 3080
rect 11333 3071 11391 3077
rect 13357 3077 13369 3080
rect 13403 3077 13415 3111
rect 13357 3071 13415 3077
rect 13449 3111 13507 3117
rect 13449 3077 13461 3111
rect 13495 3108 13507 3111
rect 13495 3080 14964 3108
rect 13495 3077 13507 3080
rect 13449 3071 13507 3077
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 10410 3040 10416 3052
rect 10192 3012 10416 3040
rect 10192 3000 10198 3012
rect 10410 3000 10416 3012
rect 10468 3040 10474 3052
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 10468 3012 10609 3040
rect 10468 3000 10474 3012
rect 10597 3009 10609 3012
rect 10643 3040 10655 3043
rect 10686 3040 10692 3052
rect 10643 3012 10692 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12250 3040 12256 3052
rect 12023 3012 12256 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 13906 3000 13912 3052
rect 13964 3040 13970 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13964 3012 14013 3040
rect 13964 3000 13970 3012
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 9600 2944 10333 2972
rect 7984 2932 7990 2944
rect 10321 2941 10333 2944
rect 10367 2972 10379 2975
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 10367 2944 11805 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12492 2944 12537 2972
rect 12492 2932 12498 2944
rect 12894 2932 12900 2984
rect 12952 2972 12958 2984
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 12952 2944 14473 2972
rect 12952 2932 12958 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 9309 2907 9367 2913
rect 9309 2873 9321 2907
rect 9355 2904 9367 2907
rect 9355 2876 9996 2904
rect 9355 2873 9367 2876
rect 9309 2867 9367 2873
rect 8662 2836 8668 2848
rect 7484 2808 8668 2836
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 8938 2836 8944 2848
rect 8899 2808 8944 2836
rect 8938 2796 8944 2808
rect 8996 2796 9002 2848
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 9766 2836 9772 2848
rect 9447 2808 9772 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 9968 2845 9996 2876
rect 10502 2864 10508 2916
rect 10560 2904 10566 2916
rect 11974 2904 11980 2916
rect 10560 2876 11980 2904
rect 10560 2864 10566 2876
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 12713 2907 12771 2913
rect 12713 2873 12725 2907
rect 12759 2904 12771 2907
rect 13170 2904 13176 2916
rect 12759 2876 13176 2904
rect 12759 2873 12771 2876
rect 12713 2867 12771 2873
rect 13170 2864 13176 2876
rect 13228 2864 13234 2916
rect 13357 2907 13415 2913
rect 13357 2873 13369 2907
rect 13403 2904 13415 2907
rect 13909 2907 13967 2913
rect 13909 2904 13921 2907
rect 13403 2876 13921 2904
rect 13403 2873 13415 2876
rect 13357 2867 13415 2873
rect 13909 2873 13921 2876
rect 13955 2873 13967 2907
rect 14936 2904 14964 3080
rect 15028 2981 15056 3148
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18417 3043 18475 3049
rect 18417 3040 18429 3043
rect 17920 3012 18429 3040
rect 17920 3000 17926 3012
rect 18417 3009 18429 3012
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 15013 2975 15071 2981
rect 15013 2941 15025 2975
rect 15059 2941 15071 2975
rect 15749 2975 15807 2981
rect 15749 2972 15761 2975
rect 15013 2935 15071 2941
rect 15120 2944 15761 2972
rect 15120 2904 15148 2944
rect 15749 2941 15761 2944
rect 15795 2941 15807 2975
rect 15749 2935 15807 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 16485 2975 16543 2981
rect 16485 2972 16497 2975
rect 15896 2944 16497 2972
rect 15896 2932 15902 2944
rect 16485 2941 16497 2944
rect 16531 2941 16543 2975
rect 16485 2935 16543 2941
rect 17037 2975 17095 2981
rect 17037 2941 17049 2975
rect 17083 2941 17095 2975
rect 17037 2935 17095 2941
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 21634 2972 21640 2984
rect 20579 2944 21640 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 14936 2876 15148 2904
rect 15289 2907 15347 2913
rect 13909 2867 13967 2873
rect 15289 2873 15301 2907
rect 15335 2904 15347 2907
rect 15930 2904 15936 2916
rect 15335 2876 15936 2904
rect 15335 2873 15347 2876
rect 15289 2867 15347 2873
rect 15930 2864 15936 2876
rect 15988 2864 15994 2916
rect 16025 2907 16083 2913
rect 16025 2873 16037 2907
rect 16071 2904 16083 2907
rect 17052 2904 17080 2935
rect 16071 2876 17080 2904
rect 18248 2904 18276 2935
rect 21634 2932 21640 2944
rect 21692 2932 21698 2984
rect 22554 2904 22560 2916
rect 18248 2876 22560 2904
rect 16071 2873 16083 2876
rect 16025 2867 16083 2873
rect 22554 2864 22560 2876
rect 22612 2864 22618 2916
rect 9953 2839 10011 2845
rect 9953 2805 9965 2839
rect 9999 2805 10011 2839
rect 9953 2799 10011 2805
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10413 2839 10471 2845
rect 10413 2836 10425 2839
rect 10192 2808 10425 2836
rect 10192 2796 10198 2808
rect 10413 2805 10425 2808
rect 10459 2836 10471 2839
rect 10962 2836 10968 2848
rect 10459 2808 10968 2836
rect 10459 2805 10471 2808
rect 10413 2799 10471 2805
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11514 2796 11520 2848
rect 11572 2836 11578 2848
rect 11701 2839 11759 2845
rect 11701 2836 11713 2839
rect 11572 2808 11713 2836
rect 11572 2796 11578 2808
rect 11701 2805 11713 2808
rect 11747 2805 11759 2839
rect 11701 2799 11759 2805
rect 13538 2796 13544 2848
rect 13596 2836 13602 2848
rect 13817 2839 13875 2845
rect 13817 2836 13829 2839
rect 13596 2808 13829 2836
rect 13596 2796 13602 2808
rect 13817 2805 13829 2808
rect 13863 2805 13875 2839
rect 13817 2799 13875 2805
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 14645 2839 14703 2845
rect 14645 2836 14657 2839
rect 14240 2808 14657 2836
rect 14240 2796 14246 2808
rect 14645 2805 14657 2808
rect 14691 2805 14703 2839
rect 14645 2799 14703 2805
rect 15838 2796 15844 2848
rect 15896 2836 15902 2848
rect 16669 2839 16727 2845
rect 16669 2836 16681 2839
rect 15896 2808 16681 2836
rect 15896 2796 15902 2808
rect 16669 2805 16681 2808
rect 16715 2805 16727 2839
rect 16669 2799 16727 2805
rect 16850 2796 16856 2848
rect 16908 2836 16914 2848
rect 17221 2839 17279 2845
rect 17221 2836 17233 2839
rect 16908 2808 17233 2836
rect 16908 2796 16914 2808
rect 17221 2805 17233 2808
rect 17267 2805 17279 2839
rect 17221 2799 17279 2805
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 22094 2836 22100 2848
rect 20763 2808 22100 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2038 2632 2044 2644
rect 1995 2604 2044 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 2314 2632 2320 2644
rect 2275 2604 2320 2632
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 2498 2632 2504 2644
rect 2455 2604 2504 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 3418 2632 3424 2644
rect 3379 2604 3424 2632
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 5350 2632 5356 2644
rect 5311 2604 5356 2632
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 6917 2635 6975 2641
rect 6917 2632 6929 2635
rect 5491 2604 6929 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 6917 2601 6929 2604
rect 6963 2601 6975 2635
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 6917 2595 6975 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 9033 2635 9091 2641
rect 9033 2632 9045 2635
rect 8628 2604 9045 2632
rect 8628 2592 8634 2604
rect 9033 2601 9045 2604
rect 9079 2601 9091 2635
rect 9766 2632 9772 2644
rect 9727 2604 9772 2632
rect 9033 2595 9091 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 10870 2632 10876 2644
rect 10744 2604 10876 2632
rect 10744 2592 10750 2604
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 12069 2635 12127 2641
rect 12069 2601 12081 2635
rect 12115 2632 12127 2635
rect 13538 2632 13544 2644
rect 12115 2604 13544 2632
rect 12115 2601 12127 2604
rect 12069 2595 12127 2601
rect 13538 2592 13544 2604
rect 13596 2592 13602 2644
rect 3326 2564 3332 2576
rect 2792 2536 3332 2564
rect 2314 2456 2320 2508
rect 2372 2496 2378 2508
rect 2792 2496 2820 2536
rect 3326 2524 3332 2536
rect 3384 2524 3390 2576
rect 5258 2524 5264 2576
rect 5316 2564 5322 2576
rect 8481 2567 8539 2573
rect 5316 2536 7512 2564
rect 5316 2524 5322 2536
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 2372 2468 2820 2496
rect 2976 2468 7297 2496
rect 2372 2456 2378 2468
rect 2590 2428 2596 2440
rect 2551 2400 2596 2428
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 2976 2369 3004 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 4246 2428 4252 2440
rect 3651 2400 4252 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 7484 2437 7512 2536
rect 8481 2533 8493 2567
rect 8527 2564 8539 2567
rect 8938 2564 8944 2576
rect 8527 2536 8944 2564
rect 8527 2533 8539 2536
rect 8481 2527 8539 2533
rect 8938 2524 8944 2536
rect 8996 2524 9002 2576
rect 9214 2524 9220 2576
rect 9272 2564 9278 2576
rect 9950 2564 9956 2576
rect 9272 2536 9956 2564
rect 9272 2524 9278 2536
rect 9950 2524 9956 2536
rect 10008 2564 10014 2576
rect 10137 2567 10195 2573
rect 10137 2564 10149 2567
rect 10008 2536 10149 2564
rect 10008 2524 10014 2536
rect 10137 2533 10149 2536
rect 10183 2533 10195 2567
rect 12434 2564 12440 2576
rect 10137 2527 10195 2533
rect 10244 2536 12440 2564
rect 10244 2496 10272 2536
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 7944 2468 10272 2496
rect 10781 2499 10839 2505
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 5500 2400 5549 2428
rect 5500 2388 5506 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 2961 2363 3019 2369
rect 2961 2329 2973 2363
rect 3007 2329 3019 2363
rect 2961 2323 3019 2329
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 4706 2360 4712 2372
rect 3292 2332 4712 2360
rect 3292 2320 3298 2332
rect 4706 2320 4712 2332
rect 4764 2320 4770 2372
rect 4985 2363 5043 2369
rect 4985 2329 4997 2363
rect 5031 2360 5043 2363
rect 7944 2360 7972 2468
rect 10781 2465 10793 2499
rect 10827 2465 10839 2499
rect 10781 2459 10839 2465
rect 11057 2499 11115 2505
rect 11057 2465 11069 2499
rect 11103 2496 11115 2499
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11103 2468 11529 2496
rect 11103 2465 11115 2468
rect 11057 2459 11115 2465
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 11517 2459 11575 2465
rect 8662 2428 8668 2440
rect 8623 2400 8668 2428
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 10134 2388 10140 2440
rect 10192 2428 10198 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 10192 2400 10241 2428
rect 10192 2388 10198 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10410 2428 10416 2440
rect 10371 2400 10416 2428
rect 10229 2391 10287 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 5031 2332 7972 2360
rect 8021 2363 8079 2369
rect 5031 2329 5043 2332
rect 4985 2323 5043 2329
rect 8021 2329 8033 2363
rect 8067 2360 8079 2363
rect 10796 2360 10824 2459
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12584 2468 12633 2496
rect 12584 2456 12590 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 13170 2496 13176 2508
rect 13131 2468 13176 2496
rect 12621 2459 12679 2465
rect 13170 2456 13176 2468
rect 13228 2456 13234 2508
rect 13722 2496 13728 2508
rect 13683 2468 13728 2496
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 14274 2496 14280 2508
rect 14235 2468 14280 2496
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14608 2468 14841 2496
rect 14608 2456 14614 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 14829 2459 14887 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 15930 2456 15936 2508
rect 15988 2496 15994 2508
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15988 2468 16037 2496
rect 15988 2456 15994 2468
rect 16025 2465 16037 2468
rect 16071 2465 16083 2499
rect 16666 2496 16672 2508
rect 16627 2468 16672 2496
rect 16025 2459 16083 2465
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 8067 2332 10824 2360
rect 8067 2329 8079 2332
rect 8021 2323 8079 2329
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 10134 2292 10140 2304
rect 7064 2264 10140 2292
rect 7064 2252 7070 2264
rect 10134 2252 10140 2264
rect 10192 2292 10198 2304
rect 10594 2292 10600 2304
rect 10192 2264 10600 2292
rect 10192 2252 10198 2264
rect 10594 2252 10600 2264
rect 10652 2252 10658 2304
rect 11701 2295 11759 2301
rect 11701 2261 11713 2295
rect 11747 2292 11759 2295
rect 12434 2292 12440 2304
rect 11747 2264 12440 2292
rect 11747 2261 11759 2264
rect 11701 2255 11759 2261
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2292 12863 2295
rect 12894 2292 12900 2304
rect 12851 2264 12900 2292
rect 12851 2261 12863 2264
rect 12805 2255 12863 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 13354 2292 13360 2304
rect 13315 2264 13360 2292
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 13909 2295 13967 2301
rect 13909 2292 13921 2295
rect 13780 2264 13921 2292
rect 13780 2252 13786 2264
rect 13909 2261 13921 2264
rect 13955 2261 13967 2295
rect 13909 2255 13967 2261
rect 14461 2295 14519 2301
rect 14461 2261 14473 2295
rect 14507 2292 14519 2295
rect 14642 2292 14648 2304
rect 14507 2264 14648 2292
rect 14507 2261 14519 2264
rect 14461 2255 14519 2261
rect 14642 2252 14648 2264
rect 14700 2252 14706 2304
rect 15013 2295 15071 2301
rect 15013 2261 15025 2295
rect 15059 2292 15071 2295
rect 15102 2292 15108 2304
rect 15059 2264 15108 2292
rect 15059 2261 15071 2264
rect 15013 2255 15071 2261
rect 15102 2252 15108 2264
rect 15160 2252 15166 2304
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15528 2264 15669 2292
rect 15528 2252 15534 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 16209 2295 16267 2301
rect 16209 2261 16221 2295
rect 16255 2292 16267 2295
rect 16390 2292 16396 2304
rect 16255 2264 16396 2292
rect 16255 2261 16267 2264
rect 16209 2255 16267 2261
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 17310 2292 17316 2304
rect 16899 2264 17316 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 3602 1980 3608 2032
rect 3660 2020 3666 2032
rect 4798 2020 4804 2032
rect 3660 1992 4804 2020
rect 3660 1980 3666 1992
rect 4798 1980 4804 1992
rect 4856 1980 4862 2032
rect 5994 1368 6000 1420
rect 6052 1408 6058 1420
rect 6730 1408 6736 1420
rect 6052 1380 6736 1408
rect 6052 1368 6058 1380
rect 6730 1368 6736 1380
rect 6788 1368 6794 1420
rect 11146 1368 11152 1420
rect 11204 1408 11210 1420
rect 11882 1408 11888 1420
rect 11204 1380 11888 1408
rect 11204 1368 11210 1380
rect 11882 1368 11888 1380
rect 11940 1368 11946 1420
rect 6178 552 6184 604
rect 6236 592 6242 604
rect 6270 592 6276 604
rect 6236 564 6276 592
rect 6236 552 6242 564
rect 6270 552 6276 564
rect 6328 552 6334 604
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 4068 19456 4120 19508
rect 1860 19252 1912 19304
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 7196 19252 7248 19304
rect 2872 19184 2924 19236
rect 2780 19116 2832 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 3792 18912 3844 18964
rect 2320 18844 2372 18896
rect 1768 18708 1820 18760
rect 7288 18819 7340 18828
rect 7288 18785 7297 18819
rect 7297 18785 7331 18819
rect 7331 18785 7340 18819
rect 7288 18776 7340 18785
rect 8484 18708 8536 18760
rect 7748 18640 7800 18692
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 2780 18368 2832 18420
rect 3056 18411 3108 18420
rect 3056 18377 3065 18411
rect 3065 18377 3099 18411
rect 3099 18377 3108 18411
rect 3056 18368 3108 18377
rect 7196 18275 7248 18284
rect 7196 18241 7205 18275
rect 7205 18241 7239 18275
rect 7239 18241 7248 18275
rect 7196 18232 7248 18241
rect 2044 18164 2096 18216
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 7104 18164 7156 18216
rect 10324 18096 10376 18148
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1768 17824 1820 17876
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 2320 17756 2372 17808
rect 7288 17756 7340 17808
rect 10324 17799 10376 17808
rect 10324 17765 10333 17799
rect 10333 17765 10367 17799
rect 10367 17765 10376 17799
rect 10324 17756 10376 17765
rect 1952 17688 2004 17740
rect 7656 17688 7708 17740
rect 9220 17688 9272 17740
rect 10692 17688 10744 17740
rect 7288 17620 7340 17672
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1768 17323 1820 17332
rect 1768 17289 1777 17323
rect 1777 17289 1811 17323
rect 1811 17289 1820 17323
rect 1768 17280 1820 17289
rect 10692 17323 10744 17332
rect 10692 17289 10701 17323
rect 10701 17289 10735 17323
rect 10735 17289 10744 17323
rect 10692 17280 10744 17289
rect 2044 17212 2096 17264
rect 6184 17187 6236 17196
rect 2044 17076 2096 17128
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 7656 17144 7708 17196
rect 1952 17008 2004 17060
rect 1676 16940 1728 16992
rect 7196 17008 7248 17060
rect 9772 17187 9824 17196
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 8760 17008 8812 17060
rect 5540 16940 5592 16992
rect 5908 16983 5960 16992
rect 5908 16949 5917 16983
rect 5917 16949 5951 16983
rect 5951 16949 5960 16983
rect 5908 16940 5960 16949
rect 6000 16983 6052 16992
rect 6000 16949 6009 16983
rect 6009 16949 6043 16983
rect 6043 16949 6052 16983
rect 6000 16940 6052 16949
rect 9128 16940 9180 16992
rect 9680 16940 9732 16992
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 3332 16779 3384 16788
rect 3332 16745 3341 16779
rect 3341 16745 3375 16779
rect 3375 16745 3384 16779
rect 3332 16736 3384 16745
rect 1860 16668 1912 16720
rect 2044 16668 2096 16720
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 5172 16668 5224 16720
rect 3148 16643 3200 16652
rect 3148 16609 3157 16643
rect 3157 16609 3191 16643
rect 3191 16609 3200 16643
rect 3148 16600 3200 16609
rect 3516 16600 3568 16652
rect 4896 16600 4948 16652
rect 6184 16736 6236 16788
rect 9128 16779 9180 16788
rect 9128 16745 9137 16779
rect 9137 16745 9171 16779
rect 9171 16745 9180 16779
rect 9128 16736 9180 16745
rect 9772 16736 9824 16788
rect 10416 16736 10468 16788
rect 11336 16736 11388 16788
rect 18972 16736 19024 16788
rect 6276 16643 6328 16652
rect 6276 16609 6310 16643
rect 6310 16609 6328 16643
rect 6276 16600 6328 16609
rect 10140 16668 10192 16720
rect 10232 16600 10284 16652
rect 11612 16643 11664 16652
rect 11612 16609 11646 16643
rect 11646 16609 11664 16643
rect 11612 16600 11664 16609
rect 5816 16532 5868 16584
rect 7932 16575 7984 16584
rect 7932 16541 7941 16575
rect 7941 16541 7975 16575
rect 7975 16541 7984 16575
rect 7932 16532 7984 16541
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 2964 16235 3016 16244
rect 2964 16201 2973 16235
rect 2973 16201 3007 16235
rect 3007 16201 3016 16235
rect 2964 16192 3016 16201
rect 4896 16235 4948 16244
rect 4896 16201 4905 16235
rect 4905 16201 4939 16235
rect 4939 16201 4948 16235
rect 4896 16192 4948 16201
rect 5172 16235 5224 16244
rect 5172 16201 5181 16235
rect 5181 16201 5215 16235
rect 5215 16201 5224 16235
rect 5172 16192 5224 16201
rect 7196 16235 7248 16244
rect 7196 16201 7205 16235
rect 7205 16201 7239 16235
rect 7239 16201 7248 16235
rect 7196 16192 7248 16201
rect 11612 16192 11664 16244
rect 3148 16056 3200 16108
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 5908 16056 5960 16108
rect 10140 16099 10192 16108
rect 2044 16031 2096 16040
rect 2044 15997 2053 16031
rect 2053 15997 2087 16031
rect 2087 15997 2096 16031
rect 2044 15988 2096 15997
rect 2688 15988 2740 16040
rect 5540 16031 5592 16040
rect 5540 15997 5549 16031
rect 5549 15997 5583 16031
rect 5583 15997 5592 16031
rect 5540 15988 5592 15997
rect 7932 15988 7984 16040
rect 4160 15920 4212 15972
rect 4804 15920 4856 15972
rect 10140 16065 10149 16099
rect 10149 16065 10183 16099
rect 10183 16065 10192 16099
rect 10140 16056 10192 16065
rect 8208 16031 8260 16040
rect 8208 15997 8224 16031
rect 8224 15997 8258 16031
rect 8258 15997 8260 16031
rect 10416 16031 10468 16040
rect 8208 15988 8260 15997
rect 10416 15997 10450 16031
rect 10450 15997 10468 16031
rect 10416 15988 10468 15997
rect 8944 15920 8996 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 2780 15852 2832 15904
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 10232 15852 10284 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 2044 15648 2096 15700
rect 5632 15648 5684 15700
rect 8944 15691 8996 15700
rect 8944 15657 8953 15691
rect 8953 15657 8987 15691
rect 8987 15657 8996 15691
rect 8944 15648 8996 15657
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 11152 15648 11204 15700
rect 2688 15580 2740 15632
rect 1952 15512 2004 15564
rect 4068 15580 4120 15632
rect 6184 15623 6236 15632
rect 6184 15589 6218 15623
rect 6218 15589 6236 15623
rect 6184 15580 6236 15589
rect 3148 15555 3200 15564
rect 3148 15521 3157 15555
rect 3157 15521 3191 15555
rect 3191 15521 3200 15555
rect 3148 15512 3200 15521
rect 4252 15512 4304 15564
rect 3332 15487 3384 15496
rect 3332 15453 3341 15487
rect 3341 15453 3375 15487
rect 3375 15453 3384 15487
rect 3332 15444 3384 15453
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 4804 15308 4856 15360
rect 5816 15512 5868 15564
rect 8208 15580 8260 15632
rect 11888 15580 11940 15632
rect 8668 15512 8720 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 11060 15512 11112 15564
rect 7472 15444 7524 15496
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 11612 15487 11664 15496
rect 6552 15308 6604 15360
rect 7564 15308 7616 15360
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 11796 15351 11848 15360
rect 11796 15317 11805 15351
rect 11805 15317 11839 15351
rect 11839 15317 11848 15351
rect 11796 15308 11848 15317
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 1676 15079 1728 15088
rect 1676 15045 1685 15079
rect 1685 15045 1719 15079
rect 1719 15045 1728 15079
rect 1676 15036 1728 15045
rect 1952 14968 2004 15020
rect 3516 15104 3568 15156
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 4252 15104 4304 15156
rect 6000 15104 6052 15156
rect 7656 15104 7708 15156
rect 8668 15104 8720 15156
rect 8576 15036 8628 15088
rect 4712 14968 4764 15020
rect 6276 15011 6328 15020
rect 6276 14977 6285 15011
rect 6285 14977 6319 15011
rect 6319 14977 6328 15011
rect 6276 14968 6328 14977
rect 7564 15011 7616 15020
rect 7564 14977 7573 15011
rect 7573 14977 7607 15011
rect 7607 14977 7616 15011
rect 7564 14968 7616 14977
rect 2872 14900 2924 14952
rect 3332 14900 3384 14952
rect 6000 14900 6052 14952
rect 7656 14900 7708 14952
rect 8208 14900 8260 14952
rect 4252 14832 4304 14884
rect 6920 14832 6972 14884
rect 11060 14900 11112 14952
rect 2688 14764 2740 14816
rect 5816 14764 5868 14816
rect 6092 14807 6144 14816
rect 6092 14773 6101 14807
rect 6101 14773 6135 14807
rect 6135 14773 6144 14807
rect 6092 14764 6144 14773
rect 7196 14764 7248 14816
rect 9404 14832 9456 14884
rect 8300 14764 8352 14816
rect 10876 14764 10928 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 3332 14560 3384 14612
rect 4160 14560 4212 14612
rect 4896 14560 4948 14612
rect 8300 14560 8352 14612
rect 4712 14492 4764 14544
rect 5908 14492 5960 14544
rect 7564 14492 7616 14544
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2872 14424 2924 14476
rect 5724 14424 5776 14476
rect 6092 14424 6144 14476
rect 6460 14424 6512 14476
rect 10048 14560 10100 14612
rect 9680 14492 9732 14544
rect 9312 14424 9364 14476
rect 10140 14492 10192 14544
rect 4988 14399 5040 14408
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 6368 14399 6420 14408
rect 5632 14288 5684 14340
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 9404 14356 9456 14408
rect 9956 14467 10008 14476
rect 9956 14433 9990 14467
rect 9990 14433 10008 14467
rect 9956 14424 10008 14433
rect 8300 14288 8352 14340
rect 9128 14288 9180 14340
rect 7380 14220 7432 14272
rect 8484 14220 8536 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 5632 14059 5684 14068
rect 5632 14025 5641 14059
rect 5641 14025 5675 14059
rect 5675 14025 5684 14059
rect 5632 14016 5684 14025
rect 6000 14016 6052 14068
rect 8392 14016 8444 14068
rect 9588 14016 9640 14068
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 3332 13880 3384 13932
rect 3516 13880 3568 13932
rect 4068 13880 4120 13932
rect 1952 13812 2004 13864
rect 2688 13812 2740 13864
rect 2872 13812 2924 13864
rect 6368 13812 6420 13864
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 8300 13812 8352 13864
rect 3056 13744 3108 13796
rect 3148 13744 3200 13796
rect 4988 13744 5040 13796
rect 5448 13744 5500 13796
rect 5908 13787 5960 13796
rect 5908 13753 5917 13787
rect 5917 13753 5951 13787
rect 5951 13753 5960 13787
rect 5908 13744 5960 13753
rect 7472 13744 7524 13796
rect 9312 13812 9364 13864
rect 9036 13744 9088 13796
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 5448 13515 5500 13524
rect 5448 13481 5457 13515
rect 5457 13481 5491 13515
rect 5491 13481 5500 13515
rect 5448 13472 5500 13481
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 6368 13472 6420 13524
rect 7380 13472 7432 13524
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 1492 13404 1544 13456
rect 1860 13379 1912 13388
rect 1860 13345 1869 13379
rect 1869 13345 1903 13379
rect 1903 13345 1912 13379
rect 1860 13336 1912 13345
rect 4160 13404 4212 13456
rect 6000 13404 6052 13456
rect 3332 13379 3384 13388
rect 3332 13345 3341 13379
rect 3341 13345 3375 13379
rect 3375 13345 3384 13379
rect 3332 13336 3384 13345
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 8576 13404 8628 13456
rect 9588 13404 9640 13456
rect 2780 13311 2832 13320
rect 2780 13277 2789 13311
rect 2789 13277 2823 13311
rect 2823 13277 2832 13311
rect 6184 13311 6236 13320
rect 2780 13268 2832 13277
rect 6184 13277 6193 13311
rect 6193 13277 6227 13311
rect 6227 13277 6236 13311
rect 6184 13268 6236 13277
rect 7012 13336 7064 13388
rect 7472 13268 7524 13320
rect 8760 13336 8812 13388
rect 10324 13336 10376 13388
rect 8852 13268 8904 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9956 13268 10008 13320
rect 7748 13200 7800 13252
rect 8668 13200 8720 13252
rect 6828 13132 6880 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 6000 12971 6052 12980
rect 6000 12937 6009 12971
rect 6009 12937 6043 12971
rect 6043 12937 6052 12971
rect 6000 12928 6052 12937
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 9680 12928 9732 12980
rect 10140 12928 10192 12980
rect 2872 12860 2924 12912
rect 6828 12860 6880 12912
rect 7472 12792 7524 12844
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 2688 12724 2740 12776
rect 4068 12724 4120 12776
rect 7288 12724 7340 12776
rect 7748 12724 7800 12776
rect 10784 12724 10836 12776
rect 2780 12656 2832 12708
rect 5172 12656 5224 12708
rect 5540 12656 5592 12708
rect 6368 12656 6420 12708
rect 8668 12656 8720 12708
rect 4712 12588 4764 12640
rect 6276 12631 6328 12640
rect 6276 12597 6285 12631
rect 6285 12597 6319 12631
rect 6319 12597 6328 12631
rect 6276 12588 6328 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 1676 12427 1728 12436
rect 1676 12393 1685 12427
rect 1685 12393 1719 12427
rect 1719 12393 1728 12427
rect 1676 12384 1728 12393
rect 1860 12384 1912 12436
rect 4160 12384 4212 12436
rect 6276 12384 6328 12436
rect 6368 12384 6420 12436
rect 6920 12384 6972 12436
rect 7564 12384 7616 12436
rect 8760 12384 8812 12436
rect 3700 12248 3752 12300
rect 1400 12180 1452 12232
rect 2780 12180 2832 12232
rect 2964 12180 3016 12232
rect 4068 12180 4120 12232
rect 4160 12112 4212 12164
rect 5080 12316 5132 12368
rect 5448 12248 5500 12300
rect 6368 12248 6420 12300
rect 7840 12248 7892 12300
rect 8300 12248 8352 12300
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 5264 12112 5316 12164
rect 6920 12180 6972 12232
rect 9956 12180 10008 12232
rect 8668 12155 8720 12164
rect 8668 12121 8677 12155
rect 8677 12121 8711 12155
rect 8711 12121 8720 12155
rect 8668 12112 8720 12121
rect 20352 12044 20404 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 2964 11840 3016 11892
rect 3700 11883 3752 11892
rect 3700 11849 3709 11883
rect 3709 11849 3743 11883
rect 3743 11849 3752 11883
rect 3700 11840 3752 11849
rect 3792 11840 3844 11892
rect 5356 11840 5408 11892
rect 5448 11840 5500 11892
rect 6368 11840 6420 11892
rect 7104 11840 7156 11892
rect 7840 11840 7892 11892
rect 7012 11815 7064 11824
rect 7012 11781 7021 11815
rect 7021 11781 7055 11815
rect 7055 11781 7064 11815
rect 7012 11772 7064 11781
rect 1584 11636 1636 11688
rect 2872 11636 2924 11688
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 4160 11636 4212 11688
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 2688 11568 2740 11620
rect 5724 11568 5776 11620
rect 9312 11568 9364 11620
rect 11060 11568 11112 11620
rect 3700 11500 3752 11552
rect 4068 11500 4120 11552
rect 8576 11500 8628 11552
rect 9128 11500 9180 11552
rect 19892 11500 19944 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 4252 11296 4304 11348
rect 4988 11296 5040 11348
rect 7748 11296 7800 11348
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 8668 11296 8720 11348
rect 9680 11296 9732 11348
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 2872 11228 2924 11280
rect 2964 11228 3016 11280
rect 3792 11228 3844 11280
rect 4252 11160 4304 11212
rect 5172 11160 5224 11212
rect 5540 11160 5592 11212
rect 6736 11160 6788 11212
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 8852 11160 8904 11212
rect 2964 11092 3016 11144
rect 2780 11024 2832 11076
rect 4804 11092 4856 11144
rect 5724 11092 5776 11144
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6368 11092 6420 11144
rect 7840 11092 7892 11144
rect 6736 11024 6788 11076
rect 9772 11160 9824 11212
rect 11152 11160 11204 11212
rect 18604 11203 18656 11212
rect 18604 11169 18619 11203
rect 18619 11169 18653 11203
rect 18653 11169 18656 11203
rect 18604 11160 18656 11169
rect 9312 11092 9364 11144
rect 9404 11024 9456 11076
rect 19432 11024 19484 11076
rect 3332 10956 3384 11008
rect 4068 10956 4120 11008
rect 11612 10956 11664 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 2872 10752 2924 10804
rect 3056 10752 3108 10804
rect 5724 10752 5776 10804
rect 9220 10752 9272 10804
rect 9772 10684 9824 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 4896 10616 4948 10668
rect 5080 10659 5132 10668
rect 5080 10625 5089 10659
rect 5089 10625 5123 10659
rect 5123 10625 5132 10659
rect 5080 10616 5132 10625
rect 11152 10616 11204 10668
rect 11612 10616 11664 10668
rect 3332 10548 3384 10600
rect 6092 10548 6144 10600
rect 5448 10480 5500 10532
rect 6828 10412 6880 10464
rect 7196 10455 7248 10464
rect 7196 10421 7205 10455
rect 7205 10421 7239 10455
rect 7239 10421 7248 10455
rect 7196 10412 7248 10421
rect 7564 10548 7616 10600
rect 7840 10548 7892 10600
rect 11060 10591 11112 10600
rect 8208 10480 8260 10532
rect 11060 10557 11069 10591
rect 11069 10557 11103 10591
rect 11103 10557 11112 10591
rect 11060 10548 11112 10557
rect 11336 10480 11388 10532
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 10784 10412 10836 10464
rect 18696 10412 18748 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 5448 10208 5500 10260
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 8208 10251 8260 10260
rect 5816 10140 5868 10192
rect 4160 10072 4212 10124
rect 4896 10072 4948 10124
rect 6920 10072 6972 10124
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 3516 10004 3568 10056
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 9864 10208 9916 10260
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 11612 10208 11664 10260
rect 10324 10072 10376 10124
rect 9036 10047 9088 10056
rect 9036 10013 9045 10047
rect 9045 10013 9079 10047
rect 9079 10013 9088 10047
rect 9036 10004 9088 10013
rect 9772 10004 9824 10056
rect 8208 9936 8260 9988
rect 4068 9868 4120 9920
rect 14372 9868 14424 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 3332 9664 3384 9716
rect 3884 9664 3936 9716
rect 4896 9707 4948 9716
rect 4896 9673 4905 9707
rect 4905 9673 4939 9707
rect 4939 9673 4948 9707
rect 4896 9664 4948 9673
rect 5172 9639 5224 9648
rect 5172 9605 5181 9639
rect 5181 9605 5215 9639
rect 5215 9605 5224 9639
rect 5172 9596 5224 9605
rect 4620 9528 4672 9580
rect 6368 9596 6420 9648
rect 6644 9596 6696 9648
rect 6920 9596 6972 9648
rect 7288 9596 7340 9648
rect 8852 9639 8904 9648
rect 8852 9605 8861 9639
rect 8861 9605 8895 9639
rect 8895 9605 8904 9639
rect 8852 9596 8904 9605
rect 11152 9664 11204 9716
rect 5724 9571 5776 9580
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 7012 9528 7064 9580
rect 8208 9528 8260 9580
rect 11152 9528 11204 9580
rect 1676 9460 1728 9512
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 4712 9460 4764 9512
rect 5540 9460 5592 9512
rect 2780 9392 2832 9444
rect 5448 9392 5500 9444
rect 8484 9460 8536 9512
rect 9680 9503 9732 9512
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 9772 9460 9824 9512
rect 8576 9392 8628 9444
rect 5816 9324 5868 9376
rect 6828 9367 6880 9376
rect 6828 9333 6837 9367
rect 6837 9333 6871 9367
rect 6871 9333 6880 9367
rect 6828 9324 6880 9333
rect 7380 9324 7432 9376
rect 7748 9324 7800 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 4620 9120 4672 9172
rect 4712 9120 4764 9172
rect 6092 9163 6144 9172
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 6368 9120 6420 9172
rect 8392 9120 8444 9172
rect 1308 9052 1360 9104
rect 2688 8984 2740 9036
rect 6736 9052 6788 9104
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 4528 8984 4580 8993
rect 5448 9027 5500 9036
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3608 8916 3660 8968
rect 5448 8993 5457 9027
rect 5457 8993 5491 9027
rect 5491 8993 5500 9027
rect 5448 8984 5500 8993
rect 5724 8984 5776 9036
rect 7840 9052 7892 9104
rect 12072 9052 12124 9104
rect 10968 8984 11020 9036
rect 3240 8848 3292 8900
rect 4988 8916 5040 8968
rect 6368 8916 6420 8968
rect 7012 8916 7064 8968
rect 1676 8780 1728 8832
rect 4804 8780 4856 8832
rect 4896 8780 4948 8832
rect 5264 8780 5316 8832
rect 8208 8848 8260 8900
rect 9680 8916 9732 8968
rect 8300 8780 8352 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 2780 8508 2832 8560
rect 1676 8372 1728 8424
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 4804 8415 4856 8424
rect 2688 8304 2740 8356
rect 4804 8381 4813 8415
rect 4813 8381 4847 8415
rect 4847 8381 4856 8415
rect 4804 8372 4856 8381
rect 7196 8508 7248 8560
rect 6552 8440 6604 8492
rect 7564 8576 7616 8628
rect 7104 8372 7156 8424
rect 3240 8304 3292 8356
rect 4068 8304 4120 8356
rect 2136 8279 2188 8288
rect 2136 8245 2145 8279
rect 2145 8245 2179 8279
rect 2179 8245 2188 8279
rect 2136 8236 2188 8245
rect 5356 8236 5408 8288
rect 6092 8279 6144 8288
rect 6092 8245 6101 8279
rect 6101 8245 6135 8279
rect 6135 8245 6144 8279
rect 6092 8236 6144 8245
rect 7196 8304 7248 8356
rect 9128 8372 9180 8424
rect 8208 8304 8260 8356
rect 10784 8576 10836 8628
rect 10968 8619 11020 8628
rect 10968 8585 10977 8619
rect 10977 8585 11011 8619
rect 11011 8585 11020 8619
rect 10968 8576 11020 8585
rect 11060 8576 11112 8628
rect 9680 8372 9732 8424
rect 11612 8372 11664 8424
rect 11704 8304 11756 8356
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 2136 8032 2188 8084
rect 4528 8032 4580 8084
rect 3056 7964 3108 8016
rect 5356 7964 5408 8016
rect 7104 8032 7156 8084
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 11704 8032 11756 8084
rect 6460 7964 6512 8016
rect 2688 7828 2740 7880
rect 4896 7896 4948 7948
rect 7104 7896 7156 7948
rect 7748 7964 7800 8016
rect 10140 7964 10192 8016
rect 15752 7964 15804 8016
rect 2136 7760 2188 7812
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 3240 7760 3292 7812
rect 6368 7828 6420 7880
rect 8208 7896 8260 7948
rect 11152 7896 11204 7948
rect 8116 7828 8168 7880
rect 2780 7692 2832 7744
rect 4896 7692 4948 7744
rect 7104 7760 7156 7812
rect 8668 7828 8720 7880
rect 10968 7828 11020 7880
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 15016 7828 15068 7880
rect 14648 7760 14700 7812
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 7288 7692 7340 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 1952 7531 2004 7540
rect 1952 7497 1961 7531
rect 1961 7497 1995 7531
rect 1995 7497 2004 7531
rect 1952 7488 2004 7497
rect 3332 7488 3384 7540
rect 5632 7488 5684 7540
rect 6092 7488 6144 7540
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 10324 7488 10376 7540
rect 17868 7488 17920 7540
rect 7104 7420 7156 7472
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 15660 7420 15712 7472
rect 8208 7352 8260 7404
rect 9680 7352 9732 7404
rect 4528 7284 4580 7336
rect 6552 7284 6604 7336
rect 7196 7327 7248 7336
rect 7196 7293 7205 7327
rect 7205 7293 7239 7327
rect 7239 7293 7248 7327
rect 7196 7284 7248 7293
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 15200 7352 15252 7404
rect 10968 7284 11020 7336
rect 11060 7284 11112 7336
rect 14648 7284 14700 7336
rect 1492 7216 1544 7268
rect 4068 7216 4120 7268
rect 9312 7216 9364 7268
rect 10784 7216 10836 7268
rect 14464 7216 14516 7268
rect 17776 7216 17828 7268
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 4712 7148 4764 7200
rect 7196 7148 7248 7200
rect 10508 7148 10560 7200
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 13176 7148 13228 7200
rect 14188 7148 14240 7200
rect 14372 7148 14424 7200
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 3332 6944 3384 6996
rect 4252 6944 4304 6996
rect 10784 6944 10836 6996
rect 3976 6876 4028 6928
rect 2504 6808 2556 6860
rect 1676 6740 1728 6792
rect 2964 6740 3016 6792
rect 4620 6808 4672 6860
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5356 6808 5408 6817
rect 5724 6851 5776 6860
rect 5724 6817 5758 6851
rect 5758 6817 5776 6851
rect 5724 6808 5776 6817
rect 7380 6851 7432 6860
rect 3976 6740 4028 6792
rect 4252 6740 4304 6792
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 5080 6740 5132 6792
rect 3240 6672 3292 6724
rect 3516 6672 3568 6724
rect 4068 6672 4120 6724
rect 7380 6817 7403 6851
rect 7403 6817 7432 6851
rect 7380 6808 7432 6817
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 10140 6740 10192 6792
rect 11704 6876 11756 6928
rect 12440 6808 12492 6860
rect 13912 6808 13964 6860
rect 15200 6808 15252 6860
rect 16028 6808 16080 6860
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 10968 6783 11020 6792
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 10968 6740 11020 6749
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 15016 6740 15068 6792
rect 17684 6740 17736 6792
rect 1584 6604 1636 6656
rect 3700 6604 3752 6656
rect 5080 6604 5132 6656
rect 9220 6672 9272 6724
rect 8484 6647 8536 6656
rect 8484 6613 8493 6647
rect 8493 6613 8527 6647
rect 8527 6613 8536 6647
rect 8484 6604 8536 6613
rect 8668 6604 8720 6656
rect 10784 6604 10836 6656
rect 11980 6604 12032 6656
rect 12348 6647 12400 6656
rect 12348 6613 12357 6647
rect 12357 6613 12391 6647
rect 12391 6613 12400 6647
rect 12348 6604 12400 6613
rect 15936 6604 15988 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2504 6400 2556 6452
rect 2964 6400 3016 6452
rect 3608 6400 3660 6452
rect 5724 6400 5776 6452
rect 4896 6264 4948 6316
rect 5816 6264 5868 6316
rect 12348 6400 12400 6452
rect 13912 6443 13964 6452
rect 7104 6332 7156 6384
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 9220 6332 9272 6384
rect 11704 6332 11756 6384
rect 11980 6332 12032 6384
rect 13912 6409 13921 6443
rect 13921 6409 13955 6443
rect 13955 6409 13964 6443
rect 13912 6400 13964 6409
rect 16948 6400 17000 6452
rect 2780 6128 2832 6180
rect 2964 6128 3016 6180
rect 4712 6196 4764 6248
rect 5632 6196 5684 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 5080 6128 5132 6180
rect 1860 6060 1912 6112
rect 4068 6060 4120 6112
rect 4252 6060 4304 6112
rect 9312 6264 9364 6316
rect 10416 6307 10468 6316
rect 8484 6239 8536 6248
rect 8484 6205 8518 6239
rect 8518 6205 8536 6239
rect 10416 6273 10425 6307
rect 10425 6273 10459 6307
rect 10459 6273 10468 6307
rect 10416 6264 10468 6273
rect 10784 6264 10836 6316
rect 11336 6264 11388 6316
rect 11612 6307 11664 6316
rect 11612 6273 11621 6307
rect 11621 6273 11655 6307
rect 11655 6273 11664 6307
rect 11612 6264 11664 6273
rect 12440 6264 12492 6316
rect 13544 6264 13596 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 8484 6196 8536 6205
rect 8760 6128 8812 6180
rect 10048 6128 10100 6180
rect 12624 6196 12676 6248
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 15660 6239 15712 6248
rect 15660 6205 15669 6239
rect 15669 6205 15703 6239
rect 15703 6205 15712 6239
rect 15660 6196 15712 6205
rect 15936 6196 15988 6248
rect 10416 6128 10468 6180
rect 5724 6060 5776 6112
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 9680 6060 9732 6112
rect 9864 6103 9916 6112
rect 9864 6069 9873 6103
rect 9873 6069 9907 6103
rect 9907 6069 9916 6103
rect 9864 6060 9916 6069
rect 10968 6060 11020 6112
rect 11336 6060 11388 6112
rect 13544 6128 13596 6180
rect 14464 6128 14516 6180
rect 17408 6128 17460 6180
rect 13728 6060 13780 6112
rect 14280 6060 14332 6112
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 16028 6060 16080 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 1492 5899 1544 5908
rect 1492 5865 1501 5899
rect 1501 5865 1535 5899
rect 1535 5865 1544 5899
rect 1492 5856 1544 5865
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 3424 5856 3476 5908
rect 4252 5856 4304 5908
rect 8300 5856 8352 5908
rect 9864 5856 9916 5908
rect 5724 5788 5776 5840
rect 6828 5788 6880 5840
rect 2872 5763 2924 5772
rect 2872 5729 2881 5763
rect 2881 5729 2915 5763
rect 2915 5729 2924 5763
rect 2872 5720 2924 5729
rect 3884 5720 3936 5772
rect 4896 5720 4948 5772
rect 5080 5720 5132 5772
rect 5632 5720 5684 5772
rect 5816 5763 5868 5772
rect 5816 5729 5850 5763
rect 5850 5729 5868 5763
rect 7564 5763 7616 5772
rect 5816 5720 5868 5729
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 9864 5720 9916 5772
rect 13176 5856 13228 5908
rect 13544 5899 13596 5908
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 14280 5899 14332 5908
rect 14280 5865 14289 5899
rect 14289 5865 14323 5899
rect 14323 5865 14332 5899
rect 14280 5856 14332 5865
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 10692 5788 10744 5840
rect 14188 5831 14240 5840
rect 14188 5797 14197 5831
rect 14197 5797 14231 5831
rect 14231 5797 14240 5831
rect 14188 5788 14240 5797
rect 16488 5788 16540 5840
rect 1584 5652 1636 5704
rect 2964 5695 3016 5704
rect 2504 5559 2556 5568
rect 2504 5525 2513 5559
rect 2513 5525 2547 5559
rect 2547 5525 2556 5559
rect 2504 5516 2556 5525
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 2688 5584 2740 5636
rect 3792 5652 3844 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 7012 5652 7064 5704
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 6552 5584 6604 5636
rect 8668 5652 8720 5704
rect 9772 5652 9824 5704
rect 9864 5584 9916 5636
rect 10048 5584 10100 5636
rect 12992 5720 13044 5772
rect 13176 5720 13228 5772
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 17684 5763 17736 5772
rect 17684 5729 17693 5763
rect 17693 5729 17727 5763
rect 17727 5729 17736 5763
rect 17684 5720 17736 5729
rect 13912 5652 13964 5704
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 2780 5516 2832 5568
rect 4068 5516 4120 5568
rect 6460 5516 6512 5568
rect 7104 5516 7156 5568
rect 8668 5516 8720 5568
rect 13820 5559 13872 5568
rect 13820 5525 13829 5559
rect 13829 5525 13863 5559
rect 13863 5525 13872 5559
rect 13820 5516 13872 5525
rect 15016 5516 15068 5568
rect 15936 5652 15988 5704
rect 17960 5516 18012 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 3148 5312 3200 5364
rect 7012 5312 7064 5364
rect 7840 5312 7892 5364
rect 2596 5176 2648 5228
rect 1860 5108 1912 5160
rect 2688 5108 2740 5160
rect 4344 5176 4396 5228
rect 3700 5108 3752 5160
rect 5632 5108 5684 5160
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 1400 5040 1452 5092
rect 2412 5040 2464 5092
rect 2964 5040 3016 5092
rect 8760 5151 8812 5160
rect 8760 5117 8769 5151
rect 8769 5117 8803 5151
rect 8803 5117 8812 5151
rect 8760 5108 8812 5117
rect 7104 5083 7156 5092
rect 7104 5049 7138 5083
rect 7138 5049 7156 5083
rect 7104 5040 7156 5049
rect 10692 5176 10744 5228
rect 12992 5219 13044 5228
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 13728 5176 13780 5228
rect 13820 5108 13872 5160
rect 16488 5176 16540 5228
rect 17408 5176 17460 5228
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 2320 4972 2372 5024
rect 3148 5015 3200 5024
rect 3148 4981 3157 5015
rect 3157 4981 3191 5015
rect 3191 4981 3200 5015
rect 3148 4972 3200 4981
rect 3332 4972 3384 5024
rect 4252 5015 4304 5024
rect 4252 4981 4261 5015
rect 4261 4981 4295 5015
rect 4295 4981 4304 5015
rect 4252 4972 4304 4981
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 6092 5015 6144 5024
rect 6092 4981 6101 5015
rect 6101 4981 6135 5015
rect 6135 4981 6144 5015
rect 6092 4972 6144 4981
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 10600 5040 10652 5092
rect 14280 5040 14332 5092
rect 14556 5040 14608 5092
rect 8300 4972 8352 5024
rect 12624 4972 12676 5024
rect 16212 5015 16264 5024
rect 16212 4981 16221 5015
rect 16221 4981 16255 5015
rect 16255 4981 16264 5015
rect 16212 4972 16264 4981
rect 16672 5015 16724 5024
rect 16672 4981 16681 5015
rect 16681 4981 16715 5015
rect 16715 4981 16724 5015
rect 16672 4972 16724 4981
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 1400 4811 1452 4820
rect 1400 4777 1409 4811
rect 1409 4777 1443 4811
rect 1443 4777 1452 4811
rect 1400 4768 1452 4777
rect 4252 4768 4304 4820
rect 6184 4768 6236 4820
rect 7564 4768 7616 4820
rect 9588 4768 9640 4820
rect 2412 4700 2464 4752
rect 2596 4632 2648 4684
rect 4068 4700 4120 4752
rect 8668 4700 8720 4752
rect 9772 4700 9824 4752
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 5724 4632 5776 4684
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 6552 4632 6604 4684
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 5816 4496 5868 4548
rect 6460 4564 6512 4616
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 7748 4496 7800 4548
rect 8760 4564 8812 4616
rect 9496 4564 9548 4616
rect 10784 4564 10836 4616
rect 11612 4564 11664 4616
rect 13636 4564 13688 4616
rect 14740 4564 14792 4616
rect 15016 4564 15068 4616
rect 16120 4632 16172 4684
rect 16212 4632 16264 4684
rect 18604 4700 18656 4752
rect 17224 4564 17276 4616
rect 10692 4496 10744 4548
rect 2228 4428 2280 4480
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 5356 4428 5408 4480
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 10048 4428 10100 4480
rect 15108 4496 15160 4548
rect 16488 4428 16540 4480
rect 16856 4471 16908 4480
rect 16856 4437 16865 4471
rect 16865 4437 16899 4471
rect 16899 4437 16908 4471
rect 16856 4428 16908 4437
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 4344 4156 4396 4208
rect 4896 4156 4948 4208
rect 204 4088 256 4140
rect 2412 4088 2464 4140
rect 1768 4020 1820 4072
rect 2780 4020 2832 4072
rect 4068 4088 4120 4140
rect 4988 4088 5040 4140
rect 3240 4063 3292 4072
rect 3240 4029 3274 4063
rect 3274 4029 3292 4063
rect 3240 4020 3292 4029
rect 4528 4020 4580 4072
rect 5724 4224 5776 4276
rect 5816 4224 5868 4276
rect 6460 4267 6512 4276
rect 6460 4233 6469 4267
rect 6469 4233 6503 4267
rect 6503 4233 6512 4267
rect 6460 4224 6512 4233
rect 8852 4224 8904 4276
rect 11612 4224 11664 4276
rect 14740 4267 14792 4276
rect 14740 4233 14749 4267
rect 14749 4233 14783 4267
rect 14783 4233 14792 4267
rect 14740 4224 14792 4233
rect 16120 4224 16172 4276
rect 16672 4267 16724 4276
rect 16672 4233 16681 4267
rect 16681 4233 16715 4267
rect 16715 4233 16724 4267
rect 16672 4224 16724 4233
rect 6920 4088 6972 4140
rect 7472 4088 7524 4140
rect 7656 4088 7708 4140
rect 7840 4088 7892 4140
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 16856 4156 16908 4208
rect 8668 4020 8720 4072
rect 9496 4020 9548 4072
rect 10048 4063 10100 4072
rect 10048 4029 10082 4063
rect 10082 4029 10100 4063
rect 10048 4020 10100 4029
rect 5448 3952 5500 4004
rect 2044 3884 2096 3936
rect 4252 3884 4304 3936
rect 4988 3884 5040 3936
rect 7288 3884 7340 3936
rect 8392 3952 8444 4004
rect 11612 4020 11664 4072
rect 12072 4020 12124 4072
rect 12624 4063 12676 4072
rect 12624 4029 12633 4063
rect 12633 4029 12667 4063
rect 12667 4029 12676 4063
rect 12624 4020 12676 4029
rect 13360 4063 13412 4072
rect 13360 4029 13369 4063
rect 13369 4029 13403 4063
rect 13403 4029 13412 4063
rect 13360 4020 13412 4029
rect 15016 4063 15068 4072
rect 8576 3884 8628 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 9220 3884 9272 3936
rect 12532 3952 12584 4004
rect 12900 3995 12952 4004
rect 12900 3961 12909 3995
rect 12909 3961 12943 3995
rect 12943 3961 12952 3995
rect 12900 3952 12952 3961
rect 11152 3927 11204 3936
rect 11152 3893 11161 3927
rect 11161 3893 11195 3927
rect 11195 3893 11204 3927
rect 11152 3884 11204 3893
rect 12440 3884 12492 3936
rect 13912 3952 13964 4004
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 13544 3884 13596 3936
rect 21180 3884 21232 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 1952 3680 2004 3732
rect 1676 3612 1728 3664
rect 2780 3612 2832 3664
rect 1860 3587 1912 3596
rect 1860 3553 1894 3587
rect 1894 3553 1912 3587
rect 1860 3544 1912 3553
rect 2964 3680 3016 3732
rect 13912 3723 13964 3732
rect 4344 3612 4396 3664
rect 3332 3544 3384 3596
rect 8668 3612 8720 3664
rect 8760 3612 8812 3664
rect 10416 3612 10468 3664
rect 11152 3655 11204 3664
rect 11152 3621 11186 3655
rect 11186 3621 11204 3655
rect 11152 3612 11204 3621
rect 5080 3544 5132 3596
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 3884 3476 3936 3528
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 6828 3476 6880 3528
rect 7840 3544 7892 3596
rect 10140 3544 10192 3596
rect 1032 3340 1084 3392
rect 2872 3408 2924 3460
rect 2596 3340 2648 3392
rect 3332 3340 3384 3392
rect 5816 3340 5868 3392
rect 6092 3408 6144 3460
rect 6460 3408 6512 3460
rect 9496 3476 9548 3528
rect 8024 3340 8076 3392
rect 8116 3340 8168 3392
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 10600 3544 10652 3596
rect 10416 3519 10468 3528
rect 10416 3485 10425 3519
rect 10425 3485 10459 3519
rect 10459 3485 10468 3519
rect 10416 3476 10468 3485
rect 10784 3408 10836 3460
rect 12256 3544 12308 3596
rect 12440 3476 12492 3528
rect 12256 3383 12308 3392
rect 12256 3349 12265 3383
rect 12265 3349 12299 3383
rect 12299 3349 12308 3383
rect 12256 3340 12308 3349
rect 13544 3340 13596 3392
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 14372 3587 14424 3596
rect 14372 3553 14381 3587
rect 14381 3553 14415 3587
rect 14415 3553 14424 3587
rect 14372 3544 14424 3553
rect 15108 3544 15160 3596
rect 17224 3587 17276 3596
rect 15844 3476 15896 3528
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 17224 3553 17233 3587
rect 17233 3553 17267 3587
rect 17267 3553 17276 3587
rect 17224 3544 17276 3553
rect 17776 3587 17828 3596
rect 17776 3553 17785 3587
rect 17785 3553 17819 3587
rect 17819 3553 17828 3587
rect 17776 3544 17828 3553
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 17684 3340 17736 3392
rect 18604 3340 18656 3392
rect 20812 3340 20864 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 1860 3136 1912 3188
rect 2228 2932 2280 2984
rect 5080 3136 5132 3188
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 5724 3179 5776 3188
rect 5724 3145 5733 3179
rect 5733 3145 5767 3179
rect 5767 3145 5776 3179
rect 5724 3136 5776 3145
rect 6092 3136 6144 3188
rect 9220 3136 9272 3188
rect 9864 3136 9916 3188
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 5448 3000 5500 3052
rect 5816 3000 5868 3052
rect 8300 3068 8352 3120
rect 6828 2932 6880 2984
rect 572 2864 624 2916
rect 1492 2796 1544 2848
rect 3424 2796 3476 2848
rect 4252 2864 4304 2916
rect 5724 2864 5776 2916
rect 7380 2864 7432 2916
rect 6092 2839 6144 2848
rect 6092 2805 6101 2839
rect 6101 2805 6135 2839
rect 6135 2805 6144 2839
rect 6092 2796 6144 2805
rect 7012 2796 7064 2848
rect 7932 2932 7984 2984
rect 10140 3000 10192 3052
rect 10416 3000 10468 3052
rect 10692 3000 10744 3052
rect 12256 3000 12308 3052
rect 13912 3000 13964 3052
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 12900 2932 12952 2984
rect 8668 2839 8720 2848
rect 8668 2805 8677 2839
rect 8677 2805 8711 2839
rect 8711 2805 8720 2839
rect 8668 2796 8720 2805
rect 8944 2839 8996 2848
rect 8944 2805 8953 2839
rect 8953 2805 8987 2839
rect 8987 2805 8996 2839
rect 8944 2796 8996 2805
rect 9772 2796 9824 2848
rect 10508 2864 10560 2916
rect 11980 2864 12032 2916
rect 13176 2864 13228 2916
rect 17868 3000 17920 3052
rect 15844 2932 15896 2984
rect 15936 2864 15988 2916
rect 21640 2932 21692 2984
rect 22560 2864 22612 2916
rect 10140 2796 10192 2848
rect 10968 2796 11020 2848
rect 11520 2796 11572 2848
rect 13544 2796 13596 2848
rect 14188 2796 14240 2848
rect 15844 2796 15896 2848
rect 16856 2796 16908 2848
rect 22100 2796 22152 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2044 2592 2096 2644
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 2504 2592 2556 2644
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 8576 2592 8628 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 10692 2592 10744 2644
rect 10876 2592 10928 2644
rect 13544 2592 13596 2644
rect 3332 2567 3384 2576
rect 2320 2456 2372 2508
rect 3332 2533 3341 2567
rect 3341 2533 3375 2567
rect 3375 2533 3384 2567
rect 3332 2524 3384 2533
rect 5264 2524 5316 2576
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 4252 2388 4304 2440
rect 5448 2388 5500 2440
rect 8944 2524 8996 2576
rect 9220 2524 9272 2576
rect 9956 2524 10008 2576
rect 12440 2524 12492 2576
rect 3240 2320 3292 2372
rect 4712 2320 4764 2372
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 10140 2388 10192 2440
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 12532 2456 12584 2508
rect 13176 2499 13228 2508
rect 13176 2465 13185 2499
rect 13185 2465 13219 2499
rect 13219 2465 13228 2499
rect 13176 2456 13228 2465
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 14556 2456 14608 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 15936 2456 15988 2508
rect 16672 2499 16724 2508
rect 16672 2465 16681 2499
rect 16681 2465 16715 2499
rect 16715 2465 16724 2499
rect 16672 2456 16724 2465
rect 7012 2252 7064 2304
rect 10140 2252 10192 2304
rect 10600 2252 10652 2304
rect 12440 2252 12492 2304
rect 12900 2252 12952 2304
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 13728 2252 13780 2304
rect 14648 2252 14700 2304
rect 15108 2252 15160 2304
rect 15476 2252 15528 2304
rect 16396 2252 16448 2304
rect 17316 2252 17368 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 3608 1980 3660 2032
rect 4804 1980 4856 2032
rect 6000 1368 6052 1420
rect 6736 1368 6788 1420
rect 11152 1368 11204 1420
rect 11888 1368 11940 1420
rect 6184 552 6236 604
rect 6276 552 6328 604
<< metal2 >>
rect 3606 22536 3662 22545
rect 3606 22471 3662 22480
rect 3054 22128 3110 22137
rect 3054 22063 3110 22072
rect 2870 21176 2926 21185
rect 2870 21111 2926 21120
rect 2778 20632 2834 20641
rect 2778 20567 2834 20576
rect 1950 20224 2006 20233
rect 1950 20159 2006 20168
rect 1964 20058 1992 20159
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1780 18766 1808 19858
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1766 18320 1822 18329
rect 1766 18255 1822 18264
rect 1780 17882 1808 18255
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1766 17368 1822 17377
rect 1766 17303 1768 17312
rect 1820 17303 1822 17312
rect 1768 17274 1820 17280
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16658 1716 16934
rect 1872 16726 1900 19246
rect 2332 18902 2360 19246
rect 2792 19174 2820 20567
rect 2884 19242 2912 21111
rect 2872 19236 2924 19242
rect 2872 19178 2924 19184
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2320 18896 2372 18902
rect 2320 18838 2372 18844
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 2792 18426 2820 18799
rect 3068 18426 3096 22063
rect 3146 21584 3202 21593
rect 3146 21519 3202 21528
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1964 17921 1992 18022
rect 1950 17912 2006 17921
rect 1950 17847 2006 17856
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 1964 17066 1992 17682
rect 2056 17270 2084 18158
rect 2332 17814 2360 18158
rect 3160 17882 3188 21519
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 2044 17264 2096 17270
rect 2044 17206 2096 17212
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 2056 16726 2084 17070
rect 3330 16960 3386 16969
rect 3330 16895 3386 16904
rect 3344 16794 3372 16895
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 1860 16720 1912 16726
rect 1860 16662 1912 16668
rect 2044 16720 2096 16726
rect 2044 16662 2096 16668
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 2962 16552 3018 16561
rect 2962 16487 3018 16496
rect 2976 16250 3004 16487
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3160 16114 3188 16594
rect 3528 16114 3556 16594
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 2044 16040 2096 16046
rect 1674 16008 1730 16017
rect 2044 15982 2096 15988
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 1674 15943 1730 15952
rect 1688 15910 1716 15943
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 2056 15706 2084 15982
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 1688 15609 1716 15642
rect 2700 15638 2728 15982
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2688 15632 2740 15638
rect 1674 15600 1730 15609
rect 2688 15574 2740 15580
rect 1674 15535 1730 15544
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1676 15088 1728 15094
rect 1674 15056 1676 15065
rect 1728 15056 1730 15065
rect 1964 15026 1992 15506
rect 1674 14991 1730 15000
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 1674 14648 1730 14657
rect 1674 14583 1676 14592
rect 1728 14583 1730 14592
rect 1676 14554 1728 14560
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1504 13462 1532 14418
rect 2700 13870 2728 14758
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 1492 13456 1544 13462
rect 1492 13398 1544 13404
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 1674 13288 1730 13297
rect 1674 13223 1730 13232
rect 1688 12442 1716 13223
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11354 1440 12174
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1596 10674 1624 11630
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1308 9104 1360 9110
rect 1308 9046 1360 9052
rect 204 4140 256 4146
rect 204 4082 256 4088
rect 216 480 244 4082
rect 1032 3392 1084 3398
rect 1032 3334 1084 3340
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 584 480 612 2858
rect 1044 480 1072 3334
rect 1320 649 1348 9046
rect 1688 8838 1716 9454
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8430 1716 8774
rect 1780 8634 1808 12718
rect 1872 12442 1900 13330
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1492 7268 1544 7274
rect 1492 7210 1544 7216
rect 1504 5914 1532 7210
rect 1688 6798 1716 8366
rect 1964 7546 1992 13806
rect 2792 13326 2820 15846
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2884 14482 2912 14894
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2884 12918 2912 13806
rect 3160 13802 3188 15506
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 3344 14958 3372 15438
rect 3528 15162 3556 16050
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3344 14618 3372 14894
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3422 14104 3478 14113
rect 3422 14039 3424 14048
rect 3476 14039 3478 14048
rect 3424 14010 3476 14016
rect 3528 13938 3556 15098
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2700 11626 2728 12718
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12238 2820 12650
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2976 11898 3004 12174
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2884 11286 2912 11630
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 10266 2820 11018
rect 2884 10810 2912 11222
rect 2976 11150 3004 11222
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2792 9178 2820 9386
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2700 8362 2728 8978
rect 2792 8566 2820 9114
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2136 8288 2188 8294
rect 2136 8230 2188 8236
rect 2148 8090 2176 8230
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2700 7886 2728 8298
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1596 5710 1624 6598
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1400 5092 1452 5098
rect 1400 5034 1452 5040
rect 1412 4826 1440 5034
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1596 2961 1624 5646
rect 1688 3670 1716 6734
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 5914 1900 6054
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4078 1808 4966
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1872 3602 1900 5102
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 3194 1900 3538
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1582 2952 1638 2961
rect 1582 2887 1638 2896
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1306 640 1362 649
rect 1306 575 1362 584
rect 1504 480 1532 2790
rect 1964 480 1992 3674
rect 2056 2650 2084 3878
rect 2148 3505 2176 7754
rect 2792 7750 2820 8366
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2516 6866 2544 7346
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2516 6458 2544 6802
rect 2976 6798 3004 11086
rect 3068 10810 3096 13738
rect 3344 13394 3372 13874
rect 3514 13696 3570 13705
rect 3514 13631 3570 13640
rect 3528 13530 3556 13631
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3344 10606 3372 10950
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10062 3372 10542
rect 3332 10056 3384 10062
rect 3146 10024 3202 10033
rect 3332 9998 3384 10004
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3146 9959 3202 9968
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3068 8022 3096 8910
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 3054 7848 3110 7857
rect 3054 7783 3110 7792
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2976 6186 3004 6394
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2412 5092 2464 5098
rect 2412 5034 2464 5040
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2240 4865 2268 4966
rect 2226 4856 2282 4865
rect 2226 4791 2282 4800
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2134 3496 2190 3505
rect 2134 3431 2190 3440
rect 2240 3369 2268 4422
rect 2226 3360 2282 3369
rect 2226 3295 2282 3304
rect 2240 2990 2268 3295
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 2332 2650 2360 4966
rect 2424 4758 2452 5034
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2424 4146 2452 4694
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2516 2650 2544 5510
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2608 4690 2636 5170
rect 2700 5166 2728 5578
rect 2792 5574 2820 6122
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2608 3398 2636 4626
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2792 3670 2820 4014
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2884 3466 2912 5714
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2976 5098 3004 5646
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2962 3904 3018 3913
rect 2962 3839 3018 3848
rect 2976 3738 3004 3839
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2332 480 2360 2450
rect 2608 2446 2636 3334
rect 3068 2553 3096 7783
rect 3160 5370 3188 9959
rect 3344 9722 3372 9998
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3528 9518 3556 9998
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3620 8974 3648 22471
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 4066 19816 4122 19825
rect 4066 19751 4122 19760
rect 4080 19514 4108 19751
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 7196 19304 7248 19310
rect 3790 19272 3846 19281
rect 7196 19246 7248 19252
rect 3790 19207 3846 19216
rect 3804 18970 3832 19207
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 7208 18290 7236 19246
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4908 16250 4936 16594
rect 5184 16250 5212 16662
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5552 16046 5580 16934
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 4080 15042 4108 15574
rect 4172 15162 4200 15914
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4264 15162 4292 15506
rect 4816 15502 4844 15914
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5644 15706 5672 15846
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5828 15570 5856 16526
rect 5920 16114 5948 16934
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4080 15014 4200 15042
rect 4172 14618 4200 15014
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4252 14884 4304 14890
rect 4252 14826 4304 14832
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4080 13394 4108 13874
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 12782 4108 13330
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4080 12322 4108 12718
rect 4172 12442 4200 13398
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3700 12300 3752 12306
rect 4080 12294 4200 12322
rect 3700 12242 3752 12248
rect 3712 11898 3740 12242
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3252 8362 3280 8842
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3252 7818 3280 8298
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3252 6730 3280 7754
rect 3330 7576 3386 7585
rect 3330 7511 3332 7520
rect 3384 7511 3386 7520
rect 3332 7482 3384 7488
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3344 7002 3372 7142
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3436 5914 3464 7142
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3160 3641 3188 4966
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4078 3280 4422
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3146 3632 3202 3641
rect 3344 3602 3372 4966
rect 3146 3567 3202 3576
rect 3332 3596 3384 3602
rect 3054 2544 3110 2553
rect 3054 2479 3110 2488
rect 2596 2440 2648 2446
rect 3160 2428 3188 3567
rect 3332 3538 3384 3544
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3344 2582 3372 3334
rect 3422 2952 3478 2961
rect 3422 2887 3478 2896
rect 3436 2854 3464 2887
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3436 2650 3464 2790
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3332 2576 3384 2582
rect 3332 2518 3384 2524
rect 2596 2382 2648 2388
rect 2792 2400 3188 2428
rect 2792 480 2820 2400
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 3252 480 3280 2314
rect 3528 1057 3556 6666
rect 3620 6458 3648 7346
rect 3712 6662 3740 11494
rect 3804 11286 3832 11834
rect 4080 11694 4108 12174
rect 4172 12170 4200 12294
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4172 11694 4200 12106
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4068 11552 4120 11558
rect 4066 11520 4068 11529
rect 4120 11520 4122 11529
rect 4066 11455 4122 11464
rect 4066 11384 4122 11393
rect 4264 11354 4292 14826
rect 4724 14550 4752 14962
rect 4816 14634 4844 15302
rect 6012 15162 6040 16934
rect 6196 16794 6224 17138
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6196 15638 6224 16730
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6288 15026 6316 16594
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 4816 14618 4936 14634
rect 4816 14612 4948 14618
rect 4816 14606 4896 14612
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4066 11319 4122 11328
rect 4252 11348 4304 11354
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 4080 11014 4108 11319
rect 4252 11290 4304 11296
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3882 10840 3938 10849
rect 3882 10775 3938 10784
rect 3896 9722 3924 10775
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4080 9926 4108 10367
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 4066 8528 4122 8537
rect 4066 8463 4122 8472
rect 4080 8362 4108 8463
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 4080 7274 4108 8055
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3974 7168 4030 7177
rect 3974 7103 4030 7112
rect 3988 6934 4016 7103
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4066 6760 4122 6769
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3698 5264 3754 5273
rect 3698 5199 3754 5208
rect 3712 5166 3740 5199
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3804 4298 3832 5646
rect 3712 4270 3832 4298
rect 3608 2032 3660 2038
rect 3608 1974 3660 1980
rect 3620 1601 3648 1974
rect 3606 1592 3662 1601
rect 3606 1527 3662 1536
rect 3514 1048 3570 1057
rect 3514 983 3570 992
rect 3712 480 3740 4270
rect 3896 4162 3924 5714
rect 3804 4134 3924 4162
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1490 0 1546 480
rect 1950 0 2006 480
rect 2318 0 2374 480
rect 2778 0 2834 480
rect 3238 0 3294 480
rect 3698 0 3754 480
rect 3804 241 3832 4134
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3896 3369 3924 3470
rect 3882 3360 3938 3369
rect 3882 3295 3938 3304
rect 3896 3058 3924 3295
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3988 2009 4016 6734
rect 4066 6695 4068 6704
rect 4120 6695 4122 6704
rect 4068 6666 4120 6672
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4080 6118 4108 6151
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4080 5574 4108 5743
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4080 4321 4108 4694
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3974 2000 4030 2009
rect 3974 1935 4030 1944
rect 4080 480 4108 4082
rect 4172 1170 4200 10066
rect 4264 7002 4292 11154
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4526 9616 4582 9625
rect 4526 9551 4582 9560
rect 4620 9580 4672 9586
rect 4540 9042 4568 9551
rect 4620 9522 4672 9528
rect 4632 9178 4660 9522
rect 4724 9518 4752 12582
rect 4816 11150 4844 14606
rect 4896 14554 4948 14560
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5000 13802 5028 14350
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5644 14074 5672 14282
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13530 5488 13738
rect 5736 13530 5764 14418
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5828 12866 5856 14758
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 5920 13802 5948 14486
rect 6012 14074 6040 14894
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6104 14482 6132 14758
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6380 13870 6408 14350
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 6012 12986 6040 13398
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5828 12838 6040 12866
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 5000 11354 5028 12174
rect 5092 11694 5120 12310
rect 5184 12238 5212 12650
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 5092 10674 5120 11630
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 4908 10130 4936 10610
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4908 9722 4936 10066
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5184 9654 5212 11154
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4724 9178 4752 9454
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4632 9058 4660 9114
rect 4528 9036 4580 9042
rect 4632 9030 4752 9058
rect 4528 8978 4580 8984
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4724 8242 4752 9030
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4816 8430 4844 8774
rect 4908 8498 4936 8774
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4724 8214 4844 8242
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4540 7886 4568 8026
rect 4528 7880 4580 7886
rect 4526 7848 4528 7857
rect 4580 7848 4582 7857
rect 4526 7783 4582 7792
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4528 7336 4580 7342
rect 4580 7284 4660 7290
rect 4528 7278 4660 7284
rect 4540 7262 4660 7278
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4264 6798 4292 6938
rect 4632 6866 4660 7262
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4724 6798 4752 7142
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4724 6254 4752 6734
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4264 5914 4292 6054
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4724 5710 4752 6190
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4264 4826 4292 4966
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4356 4706 4384 5170
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4264 4678 4384 4706
rect 4264 3942 4292 4678
rect 4724 4593 4752 4966
rect 4710 4584 4766 4593
rect 4710 4519 4766 4528
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4264 2922 4292 3878
rect 4356 3670 4384 4150
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4540 3534 4568 4014
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4264 2446 4292 2858
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4724 2378 4752 4519
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4816 2038 4844 8214
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4908 7750 4936 7890
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 5778 4936 6258
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4908 4214 4936 4626
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 5000 4146 5028 8910
rect 5276 8838 5304 12106
rect 5460 11898 5488 12242
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5368 11778 5396 11834
rect 5552 11778 5580 12650
rect 5368 11750 5580 11778
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5460 10266 5488 10474
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5552 9625 5580 11154
rect 5736 11150 5764 11562
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5736 10810 5764 11086
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5538 9616 5594 9625
rect 5736 9586 5764 10202
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5538 9551 5594 9560
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5460 9042 5488 9386
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 8022 5396 8230
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5368 6866 5396 7958
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 6662 5120 6734
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6186 5120 6598
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5092 5778 5120 6122
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 4172 1142 4568 1170
rect 4540 480 4568 1142
rect 5000 480 5028 3878
rect 5092 3602 5120 4558
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5092 3194 5120 3538
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5276 2582 5304 3130
rect 5368 2650 5396 4422
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5460 3058 5488 3946
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 5460 2446 5488 2994
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5552 2292 5580 9454
rect 5828 9382 5856 10134
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5736 8634 5764 8978
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5644 6254 5672 7482
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5736 6458 5764 6802
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5828 6322 5856 9318
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5846 5764 6054
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5644 5166 5672 5714
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5644 4570 5672 5102
rect 5736 4690 5764 5782
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5644 4542 5764 4570
rect 5828 4554 5856 5714
rect 5736 4282 5764 4542
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5828 4282 5856 4490
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5736 2922 5764 3130
rect 5828 3058 5856 3334
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5460 2264 5580 2292
rect 5460 480 5488 2264
rect 5920 480 5948 11086
rect 6012 1426 6040 12838
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6104 9178 6132 10542
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6104 7546 6132 8230
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6196 5114 6224 13262
rect 6380 12714 6408 13466
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6288 12442 6316 12582
rect 6380 12442 6408 12650
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6380 11898 6408 12242
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6380 11150 6408 11834
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6380 9178 6408 9590
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6380 7886 6408 8910
rect 6472 8022 6500 14418
rect 6564 12322 6592 15302
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13190 6868 13806
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6840 12918 6868 13126
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6564 12294 6684 12322
rect 6656 9654 6684 12294
rect 6840 12220 6868 12854
rect 6932 12442 6960 14826
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6920 12232 6972 12238
rect 6840 12192 6920 12220
rect 6920 12174 6972 12180
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 11082 6776 11154
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6748 9110 6776 11018
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 9382 6868 10406
rect 6932 10130 6960 12174
rect 7024 11830 7052 13330
rect 7116 11898 7144 18158
rect 7300 17814 7328 18770
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 7288 17808 7340 17814
rect 7288 17750 7340 17756
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7208 16250 7236 17002
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7012 11824 7064 11830
rect 7208 11778 7236 14758
rect 7300 12782 7328 17614
rect 7668 17202 7696 17682
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 13530 7420 14214
rect 7484 13802 7512 15438
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 15026 7604 15302
rect 7668 15162 7696 15846
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7576 14550 7604 14962
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7472 13796 7524 13802
rect 7472 13738 7524 13744
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7484 12850 7512 13262
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7576 12186 7604 12378
rect 7012 11766 7064 11772
rect 7116 11750 7236 11778
rect 7484 12158 7604 12186
rect 7116 11529 7144 11750
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7102 11520 7158 11529
rect 7102 11455 7158 11464
rect 7208 10470 7236 11630
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6564 7750 6592 8434
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7342 6592 7686
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5846 6868 6054
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6196 5086 6316 5114
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6104 3466 6132 4966
rect 6196 4826 6224 4966
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6104 2854 6132 3130
rect 6092 2848 6144 2854
rect 6288 2836 6316 5086
rect 6472 4622 6500 5510
rect 6564 4690 6592 5578
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6734 4720 6790 4729
rect 6552 4684 6604 4690
rect 6734 4655 6790 4664
rect 6552 4626 6604 4632
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6472 3466 6500 4218
rect 6748 3641 6776 4655
rect 6734 3632 6790 3641
rect 6734 3567 6736 3576
rect 6788 3567 6790 3576
rect 6736 3538 6788 3544
rect 6840 3534 6868 5102
rect 6932 4842 6960 9590
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7024 8974 7052 9522
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7208 8566 7236 10406
rect 7300 9654 7328 11154
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7116 8090 7144 8366
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7116 7818 7144 7890
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7116 7478 7144 7754
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7208 7342 7236 8298
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7410 7328 7686
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7116 6390 7144 6734
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7208 6254 7236 7142
rect 7392 7018 7420 9318
rect 7300 6990 7420 7018
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7024 5370 7052 5646
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7116 5098 7144 5510
rect 7104 5092 7156 5098
rect 7156 5052 7236 5080
rect 7104 5034 7156 5040
rect 6932 4814 7144 4842
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 4146 6960 4626
rect 7116 4468 7144 4814
rect 7208 4622 7236 5052
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7116 4440 7236 4468
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6840 2990 6868 3470
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6092 2790 6144 2796
rect 6196 2808 6316 2836
rect 7012 2848 7064 2854
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 6196 610 6224 2808
rect 7012 2790 7064 2796
rect 7024 2310 7052 2790
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6736 1420 6788 1426
rect 6736 1362 6788 1368
rect 6184 604 6236 610
rect 6184 546 6236 552
rect 6276 604 6328 610
rect 6276 546 6328 552
rect 6288 480 6316 546
rect 6748 480 6776 1362
rect 7208 480 7236 4440
rect 7300 3942 7328 6990
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 6322 7420 6802
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7484 4146 7512 12158
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7576 8634 7604 10542
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7576 4826 7604 5714
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7668 4264 7696 14894
rect 7760 13258 7788 18634
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 7944 16046 7972 16526
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15638 8248 15982
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8220 14958 8248 15574
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8312 14618 8340 14758
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8312 13870 8340 14282
rect 8496 14278 8524 18702
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 10324 18148 10376 18154
rect 10324 18090 10376 18096
rect 10336 17814 10364 18090
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 10324 17808 10376 17814
rect 10324 17750 10376 17756
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8680 15162 8708 15506
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7760 11354 7788 12718
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7852 11898 7880 12242
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7852 10606 7880 11086
rect 8220 10690 8248 13670
rect 8298 12744 8354 12753
rect 8298 12679 8354 12688
rect 8312 12306 8340 12679
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8220 10662 8340 10690
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8220 10266 8248 10474
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8312 10146 8340 10662
rect 8220 10118 8340 10146
rect 8220 9994 8248 10118
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8220 9586 8248 9930
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 8022 7788 9318
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8404 9178 8432 14010
rect 8588 13462 8616 15030
rect 8772 13546 8800 17002
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9140 16794 9168 16934
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 8944 15972 8996 15978
rect 8944 15914 8996 15920
rect 8956 15706 8984 15914
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 8680 13518 8800 13546
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8680 13258 8708 13518
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8680 12170 8708 12650
rect 8772 12442 8800 13330
rect 8852 13320 8904 13326
rect 9048 13274 9076 13738
rect 9140 13326 9168 14282
rect 8904 13268 9076 13274
rect 8852 13262 9076 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8864 13246 9076 13262
rect 9048 12986 9076 13246
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 9126 12336 9182 12345
rect 9126 12271 9182 12280
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8666 11792 8722 11801
rect 8666 11727 8722 11736
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 11354 8616 11494
rect 8680 11354 8708 11727
rect 9140 11558 9168 12271
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8864 9654 8892 11154
rect 9232 10810 9260 17682
rect 10704 17338 10732 17682
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 18970 17232 19026 17241
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 11336 17196 11388 17202
rect 18970 17167 19026 17176
rect 11336 17138 11388 17144
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 15706 9720 16934
rect 9784 16794 9812 17138
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10152 16114 10180 16662
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9324 13870 9352 14418
rect 9416 14414 9444 14826
rect 10060 14618 10088 15506
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10152 14550 10180 16050
rect 10244 15910 10272 16594
rect 10428 16046 10456 16730
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10244 15502 10272 15846
rect 11164 15706 11192 16934
rect 11348 16794 11376 17138
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 18984 16794 19012 17167
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11624 16250 11652 16594
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 11072 14958 11100 15506
rect 11624 15502 11652 16186
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9600 13462 9628 14010
rect 9692 13530 9720 14486
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9968 13326 9996 14010
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 10152 12986 10180 14486
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 9312 11756 9364 11762
rect 9508 11750 9628 11778
rect 9508 11744 9536 11750
rect 9364 11716 9536 11744
rect 9312 11698 9364 11704
rect 9600 11676 9628 11750
rect 9692 11676 9720 12922
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9600 11648 9812 11676
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9324 11150 9352 11562
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9692 11257 9720 11290
rect 9678 11248 9734 11257
rect 9784 11218 9812 11648
rect 9678 11183 9734 11192
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8850 9480 8906 9489
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 7840 9104 7892 9110
rect 7838 9072 7840 9081
rect 7892 9072 7894 9081
rect 7838 9007 7894 9016
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8362 8248 8842
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 8220 7954 8248 8298
rect 8312 8090 8340 8774
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7546 8156 7822
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8220 7410 8248 7890
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8496 7342 8524 9454
rect 8576 9444 8628 9450
rect 8850 9415 8906 9424
rect 8576 9386 8628 9392
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6254 8524 6598
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8588 6066 8616 9386
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 7886 8708 8230
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8496 6038 8616 6066
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7852 5370 7880 5646
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 8312 5030 8340 5850
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8300 4616 8352 4622
rect 8298 4584 8300 4593
rect 8352 4584 8354 4593
rect 7748 4548 7800 4554
rect 8298 4519 8354 4528
rect 7748 4490 7800 4496
rect 7576 4236 7696 4264
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7392 2650 7420 2858
rect 7576 2802 7604 4236
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7668 3516 7696 4082
rect 7760 3618 7788 4490
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 4146 7880 4422
rect 7840 4140 7892 4146
rect 8300 4140 8352 4146
rect 7840 4082 7892 4088
rect 8220 4100 8300 4128
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8220 3618 8248 4100
rect 8300 4082 8352 4088
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 7760 3602 7880 3618
rect 7760 3596 7892 3602
rect 7760 3590 7840 3596
rect 7840 3538 7892 3544
rect 7944 3590 8248 3618
rect 7668 3488 7788 3516
rect 7567 2774 7604 2802
rect 7567 2666 7595 2774
rect 7380 2644 7432 2650
rect 7567 2638 7696 2666
rect 7380 2586 7432 2592
rect 7668 480 7696 2638
rect 7760 1442 7788 3488
rect 7944 2990 7972 3590
rect 8128 3398 8156 3590
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8036 3210 8064 3334
rect 8036 3182 8340 3210
rect 8312 3126 8340 3182
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8404 2650 8432 3946
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 7760 1414 8064 1442
rect 8036 480 8064 1414
rect 8496 480 8524 6038
rect 8680 5710 8708 6598
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 4758 8708 5510
rect 8772 5166 8800 6122
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8772 4622 8800 5102
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8864 4282 8892 9415
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 2650 8616 3878
rect 8680 3670 8708 4014
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8772 3670 8800 3878
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8680 2446 8708 2790
rect 8956 2582 8984 2790
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9048 1170 9076 9998
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9140 3942 9168 8366
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9232 6390 9260 6666
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9324 6322 9352 7210
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9218 4584 9274 4593
rect 9218 4519 9274 4528
rect 9232 3942 9260 4519
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9232 2582 9260 3130
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 8956 1142 9076 1170
rect 8956 480 8984 1142
rect 9416 480 9444 11018
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9784 10062 9812 10678
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10266 9904 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9784 9518 9812 9998
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9692 8974 9720 9454
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9692 8430 9720 8910
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 7410 9720 8366
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9680 6112 9732 6118
rect 9864 6112 9916 6118
rect 9732 6060 9812 6066
rect 9680 6054 9812 6060
rect 9864 6054 9916 6060
rect 9692 6038 9812 6054
rect 9784 5710 9812 6038
rect 9876 5914 9904 6054
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9862 5808 9918 5817
rect 9862 5743 9864 5752
rect 9916 5743 9918 5752
rect 9864 5714 9916 5720
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9508 4826 9628 4842
rect 9508 4820 9640 4826
rect 9508 4814 9588 4820
rect 9508 4729 9536 4814
rect 9588 4762 9640 4768
rect 9784 4758 9812 5646
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9876 4865 9904 5578
rect 9862 4856 9918 4865
rect 9862 4791 9918 4800
rect 9772 4752 9824 4758
rect 9494 4720 9550 4729
rect 9772 4694 9824 4700
rect 9494 4655 9550 4664
rect 9496 4616 9548 4622
rect 9968 4570 9996 12174
rect 10336 11064 10364 13330
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10244 11036 10364 11064
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10152 6798 10180 7958
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10060 5642 10088 6122
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9496 4558 9548 4564
rect 9508 4078 9536 4558
rect 9692 4542 9996 4570
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9508 3534 9536 4014
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9692 1170 9720 4542
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4078 10088 4422
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10152 3924 10180 6734
rect 9968 3896 10180 3924
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9876 3194 9904 3334
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9784 2650 9812 2790
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9968 2582 9996 3896
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10152 3058 10180 3538
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10138 2952 10194 2961
rect 10138 2887 10194 2896
rect 10152 2854 10180 2887
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10152 2310 10180 2382
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 9692 1142 9812 1170
rect 9784 480 9812 1142
rect 10244 480 10272 11036
rect 10796 10470 10824 12718
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10336 7546 10364 10066
rect 10796 8634 10824 10406
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10428 6186 10456 6258
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10428 3534 10456 3606
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10428 2446 10456 2994
rect 10520 2922 10548 7142
rect 10796 7002 10824 7210
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6322 10824 6598
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10704 5234 10732 5782
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10600 5092 10652 5098
rect 10600 5034 10652 5040
rect 10612 3602 10640 5034
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10612 2310 10640 3538
rect 10704 3058 10732 4490
rect 10796 3466 10824 4558
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10888 2650 10916 14758
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 11354 11100 11562
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11164 10674 11192 11154
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11624 10674 11652 10950
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10980 8634 11008 8978
rect 11072 8634 11100 10542
rect 11164 9722 11192 10610
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11348 10266 11376 10474
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10980 7886 11008 8570
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11072 7342 11100 8570
rect 11164 7954 11192 9522
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8430 11652 10202
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11716 8090 11744 8298
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11716 7886 11744 8026
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10980 6798 11008 7278
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11716 6934 11744 7142
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 10968 6792 11020 6798
rect 11716 6780 11744 6870
rect 10968 6734 11020 6740
rect 11624 6752 11744 6780
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11624 6322 11652 6752
rect 11704 6384 11756 6390
rect 11702 6352 11704 6361
rect 11756 6352 11758 6361
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11612 6316 11664 6322
rect 11702 6287 11758 6296
rect 11612 6258 11664 6264
rect 11348 6118 11376 6258
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 10980 2854 11008 6054
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11624 4282 11652 4558
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11164 3670 11192 3878
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11624 3074 11652 4014
rect 11532 3046 11652 3074
rect 11532 2854 11560 3046
rect 11808 2972 11836 15302
rect 11624 2944 11836 2972
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10704 480 10732 2586
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 11164 480 11192 1362
rect 11624 480 11652 2944
rect 11900 1426 11928 15574
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 18602 11248 18658 11257
rect 18602 11183 18604 11192
rect 18656 11183 18658 11192
rect 18604 11154 18656 11160
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 6390 12020 6598
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 12084 4078 12112 9046
rect 14384 7206 14412 9862
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14660 7342 14688 7754
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6458 12388 6598
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12452 6322 12480 6802
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12452 3942 12480 6258
rect 12636 6254 12664 6734
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 13188 5914 13216 7142
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13924 6458 13952 6802
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 6186 13584 6258
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 13556 5914 13584 6122
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13188 5778 13216 5850
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13004 5234 13032 5714
rect 13740 5234 13768 6054
rect 13924 5710 13952 6394
rect 14200 5846 14228 7142
rect 14476 6186 14504 7210
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 15028 6798 15056 7822
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15212 6866 15240 7346
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14554 6352 14610 6361
rect 14554 6287 14610 6296
rect 14568 6254 14596 6287
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14292 5914 14320 6054
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 15028 5574 15056 6734
rect 15580 6118 15608 7142
rect 15672 6254 15700 7414
rect 15764 6644 15792 7958
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 15936 6656 15988 6662
rect 15764 6616 15936 6644
rect 15764 6322 15792 6616
rect 15936 6598 15988 6604
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15290 5808 15346 5817
rect 15290 5743 15292 5752
rect 15344 5743 15346 5752
rect 15292 5714 15344 5720
rect 15948 5710 15976 6190
rect 16040 6118 16068 6802
rect 16960 6458 16988 6802
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 17420 5914 17448 6122
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13832 5166 13860 5510
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 14280 5092 14332 5098
rect 14280 5034 14332 5040
rect 14556 5092 14608 5098
rect 14556 5034 14608 5040
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 4078 12664 4966
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 12624 4072 12676 4078
rect 13360 4072 13412 4078
rect 12624 4014 12676 4020
rect 13358 4040 13360 4049
rect 13412 4040 13414 4049
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12900 4004 12952 4010
rect 13358 3975 13414 3984
rect 12900 3946 12952 3952
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 3398 12296 3538
rect 12452 3534 12480 3878
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12268 3058 12296 3334
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11888 1420 11940 1426
rect 11888 1362 11940 1368
rect 11992 480 12020 2858
rect 12452 2582 12480 2926
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12544 2514 12572 3946
rect 12912 2990 12940 3946
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3398 13584 3878
rect 13648 3754 13676 4558
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13648 3726 13768 3754
rect 13924 3738 13952 3946
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 13188 2514 13216 2858
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13556 2650 13584 2790
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13740 2514 13768 3726
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13924 3058 13952 3674
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 12452 480 12480 2246
rect 12912 480 12940 2246
rect 13372 480 13400 2246
rect 13740 480 13768 2246
rect 14200 480 14228 2790
rect 14292 2514 14320 5034
rect 14370 4856 14426 4865
rect 14370 4791 14426 4800
rect 14384 3602 14412 4791
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14568 2514 14596 5034
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15028 4622 15056 5510
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 14752 4282 14780 4558
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 15028 4078 15056 4558
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15016 4072 15068 4078
rect 15014 4040 15016 4049
rect 15068 4040 15070 4049
rect 15014 3975 15070 3984
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 15120 3602 15148 4490
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15488 2514 15516 5646
rect 16500 5234 16528 5782
rect 17420 5234 17448 5850
rect 17696 5778 17724 6734
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16224 4690 16252 4966
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16132 4282 16160 4626
rect 16500 4486 16528 5170
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16684 4282 16712 4966
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16132 3534 16160 4218
rect 16868 4214 16896 4422
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 17236 3602 17264 4558
rect 17788 3602 17816 7210
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 15856 2990 15884 3470
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15936 2916 15988 2922
rect 15936 2858 15988 2864
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 14660 480 14688 2246
rect 15120 480 15148 2246
rect 15488 480 15516 2246
rect 15856 1442 15884 2790
rect 15948 2514 15976 2858
rect 16684 2514 16712 3470
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 15856 1414 15976 1442
rect 15948 480 15976 1414
rect 16408 480 16436 2246
rect 16868 480 16896 2790
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 480 17356 2246
rect 17696 480 17724 3334
rect 17880 3058 17908 7482
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18602 5808 18658 5817
rect 18602 5743 18658 5752
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17972 1986 18000 5510
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18616 4758 18644 5743
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1958 18184 1986
rect 18156 480 18184 1958
rect 18616 480 18644 3334
rect 18708 626 18736 10406
rect 18708 598 19104 626
rect 19076 480 19104 598
rect 19444 480 19472 11018
rect 19904 480 19932 11494
rect 20364 480 20392 12038
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20824 480 20852 3334
rect 21192 480 21220 3878
rect 21640 2984 21692 2990
rect 21640 2926 21692 2932
rect 21652 480 21680 2926
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22112 480 22140 2790
rect 22572 480 22600 2858
rect 3790 232 3846 241
rect 3790 167 3846 176
rect 4066 0 4122 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5446 0 5502 480
rect 5906 0 5962 480
rect 6274 0 6330 480
rect 6734 0 6790 480
rect 7194 0 7250 480
rect 7654 0 7710 480
rect 8022 0 8078 480
rect 8482 0 8538 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10230 0 10286 480
rect 10690 0 10746 480
rect 11150 0 11206 480
rect 11610 0 11666 480
rect 11978 0 12034 480
rect 12438 0 12494 480
rect 12898 0 12954 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14646 0 14702 480
rect 15106 0 15162 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16394 0 16450 480
rect 16854 0 16910 480
rect 17314 0 17370 480
rect 17682 0 17738 480
rect 18142 0 18198 480
rect 18602 0 18658 480
rect 19062 0 19118 480
rect 19430 0 19486 480
rect 19890 0 19946 480
rect 20350 0 20406 480
rect 20810 0 20866 480
rect 21178 0 21234 480
rect 21638 0 21694 480
rect 22098 0 22154 480
rect 22558 0 22614 480
<< via2 >>
rect 3606 22480 3662 22536
rect 3054 22072 3110 22128
rect 2870 21120 2926 21176
rect 2778 20576 2834 20632
rect 1950 20168 2006 20224
rect 1766 18264 1822 18320
rect 1766 17332 1822 17368
rect 1766 17312 1768 17332
rect 1768 17312 1820 17332
rect 1820 17312 1822 17332
rect 2778 18808 2834 18864
rect 3146 21528 3202 21584
rect 1950 17856 2006 17912
rect 3330 16904 3386 16960
rect 2962 16496 3018 16552
rect 1674 15952 1730 16008
rect 1674 15544 1730 15600
rect 1674 15036 1676 15056
rect 1676 15036 1728 15056
rect 1728 15036 1730 15056
rect 1674 15000 1730 15036
rect 1674 14612 1730 14648
rect 1674 14592 1676 14612
rect 1676 14592 1728 14612
rect 1728 14592 1730 14612
rect 1674 13232 1730 13288
rect 3422 14068 3478 14104
rect 3422 14048 3424 14068
rect 3424 14048 3476 14068
rect 3476 14048 3478 14068
rect 1582 2896 1638 2952
rect 1306 584 1362 640
rect 3514 13640 3570 13696
rect 3146 9968 3202 10024
rect 3054 7792 3110 7848
rect 2226 4800 2282 4856
rect 2134 3440 2190 3496
rect 2226 3304 2282 3360
rect 2962 3848 3018 3904
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 4066 19760 4122 19816
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 3790 19216 3846 19272
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 3330 7540 3386 7576
rect 3330 7520 3332 7540
rect 3332 7520 3384 7540
rect 3384 7520 3386 7540
rect 3146 3576 3202 3632
rect 3054 2488 3110 2544
rect 3422 2896 3478 2952
rect 4066 11500 4068 11520
rect 4068 11500 4120 11520
rect 4120 11500 4122 11520
rect 4066 11464 4122 11500
rect 4066 11328 4122 11384
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 3882 10784 3938 10840
rect 4066 10376 4122 10432
rect 4066 8472 4122 8528
rect 4066 8064 4122 8120
rect 3974 7112 4030 7168
rect 3698 5208 3754 5264
rect 3606 1536 3662 1592
rect 3514 992 3570 1048
rect 3882 3304 3938 3360
rect 4066 6724 4122 6760
rect 4066 6704 4068 6724
rect 4068 6704 4120 6724
rect 4120 6704 4122 6724
rect 4066 6160 4122 6216
rect 4066 5752 4122 5808
rect 4066 4256 4122 4312
rect 3974 1944 4030 2000
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4526 9560 4582 9616
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4526 7828 4528 7848
rect 4528 7828 4580 7848
rect 4580 7828 4582 7848
rect 4526 7792 4582 7828
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4710 4528 4766 4584
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5538 9560 5594 9616
rect 7102 11464 7158 11520
rect 6734 4664 6790 4720
rect 6734 3596 6790 3632
rect 6734 3576 6736 3596
rect 6736 3576 6788 3596
rect 6788 3576 6790 3596
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 8298 12688 8354 12744
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 9126 12280 9182 12336
rect 8666 11736 8722 11792
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18970 17176 19026 17232
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 9678 11192 9734 11248
rect 7838 9052 7840 9072
rect 7840 9052 7892 9072
rect 7892 9052 7894 9072
rect 7838 9016 7894 9052
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 8850 9424 8906 9480
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 8298 4564 8300 4584
rect 8300 4564 8352 4584
rect 8352 4564 8354 4584
rect 8298 4528 8354 4564
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 9218 4528 9274 4584
rect 9862 5772 9918 5808
rect 9862 5752 9864 5772
rect 9864 5752 9916 5772
rect 9916 5752 9918 5772
rect 9862 4800 9918 4856
rect 9494 4664 9550 4720
rect 10138 2896 10194 2952
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11702 6332 11704 6352
rect 11704 6332 11756 6352
rect 11756 6332 11758 6352
rect 11702 6296 11758 6332
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 18602 11212 18658 11248
rect 18602 11192 18604 11212
rect 18604 11192 18656 11212
rect 18656 11192 18658 11212
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14554 6296 14610 6352
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 15290 5772 15346 5808
rect 15290 5752 15292 5772
rect 15292 5752 15344 5772
rect 15344 5752 15346 5772
rect 13358 4020 13360 4040
rect 13360 4020 13412 4040
rect 13412 4020 13414 4040
rect 13358 3984 13414 4020
rect 14370 4800 14426 4856
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 15014 4020 15016 4040
rect 15016 4020 15068 4040
rect 15068 4020 15070 4040
rect 15014 3984 15070 4020
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18602 5752 18658 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 3790 176 3846 232
<< metal3 >>
rect 0 22538 480 22568
rect 3601 22538 3667 22541
rect 0 22536 3667 22538
rect 0 22480 3606 22536
rect 3662 22480 3667 22536
rect 0 22478 3667 22480
rect 0 22448 480 22478
rect 3601 22475 3667 22478
rect 0 22130 480 22160
rect 3049 22130 3115 22133
rect 0 22128 3115 22130
rect 0 22072 3054 22128
rect 3110 22072 3115 22128
rect 0 22070 3115 22072
rect 0 22040 480 22070
rect 3049 22067 3115 22070
rect 0 21586 480 21616
rect 3141 21586 3207 21589
rect 0 21584 3207 21586
rect 0 21528 3146 21584
rect 3202 21528 3207 21584
rect 0 21526 3207 21528
rect 0 21496 480 21526
rect 3141 21523 3207 21526
rect 0 21178 480 21208
rect 2865 21178 2931 21181
rect 0 21176 2931 21178
rect 0 21120 2870 21176
rect 2926 21120 2931 21176
rect 0 21118 2931 21120
rect 0 21088 480 21118
rect 2865 21115 2931 21118
rect 0 20634 480 20664
rect 2773 20634 2839 20637
rect 0 20632 2839 20634
rect 0 20576 2778 20632
rect 2834 20576 2839 20632
rect 0 20574 2839 20576
rect 0 20544 480 20574
rect 2773 20571 2839 20574
rect 0 20226 480 20256
rect 1945 20226 2011 20229
rect 0 20224 2011 20226
rect 0 20168 1950 20224
rect 2006 20168 2011 20224
rect 0 20166 2011 20168
rect 0 20136 480 20166
rect 1945 20163 2011 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 4061 19818 4127 19821
rect 0 19816 4127 19818
rect 0 19760 4066 19816
rect 4122 19760 4127 19816
rect 0 19758 4127 19760
rect 0 19728 480 19758
rect 4061 19755 4127 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 3785 19274 3851 19277
rect 0 19272 3851 19274
rect 0 19216 3790 19272
rect 3846 19216 3851 19272
rect 0 19214 3851 19216
rect 0 19184 480 19214
rect 3785 19211 3851 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 0 18866 480 18896
rect 2773 18866 2839 18869
rect 0 18864 2839 18866
rect 0 18808 2778 18864
rect 2834 18808 2839 18864
rect 0 18806 2839 18808
rect 0 18776 480 18806
rect 2773 18803 2839 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1761 18322 1827 18325
rect 0 18320 1827 18322
rect 0 18264 1766 18320
rect 1822 18264 1827 18320
rect 0 18262 1827 18264
rect 0 18232 480 18262
rect 1761 18259 1827 18262
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1945 17914 2011 17917
rect 0 17912 2011 17914
rect 0 17856 1950 17912
rect 2006 17856 2011 17912
rect 0 17854 2011 17856
rect 0 17824 480 17854
rect 1945 17851 2011 17854
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1761 17370 1827 17373
rect 0 17368 1827 17370
rect 0 17312 1766 17368
rect 1822 17312 1827 17368
rect 0 17310 1827 17312
rect 0 17280 480 17310
rect 1761 17307 1827 17310
rect 18965 17234 19031 17237
rect 22320 17234 22800 17264
rect 18965 17232 22800 17234
rect 18965 17176 18970 17232
rect 19026 17176 22800 17232
rect 18965 17174 22800 17176
rect 18965 17171 19031 17174
rect 22320 17144 22800 17174
rect 0 16962 480 16992
rect 3325 16962 3391 16965
rect 0 16960 3391 16962
rect 0 16904 3330 16960
rect 3386 16904 3391 16960
rect 0 16902 3391 16904
rect 0 16872 480 16902
rect 3325 16899 3391 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 0 16554 480 16584
rect 2957 16554 3023 16557
rect 0 16552 3023 16554
rect 0 16496 2962 16552
rect 3018 16496 3023 16552
rect 0 16494 3023 16496
rect 0 16464 480 16494
rect 2957 16491 3023 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 1669 16010 1735 16013
rect 0 16008 1735 16010
rect 0 15952 1674 16008
rect 1730 15952 1735 16008
rect 0 15950 1735 15952
rect 0 15920 480 15950
rect 1669 15947 1735 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 1669 15602 1735 15605
rect 0 15600 1735 15602
rect 0 15544 1674 15600
rect 1730 15544 1735 15600
rect 0 15542 1735 15544
rect 0 15512 480 15542
rect 1669 15539 1735 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 1669 15058 1735 15061
rect 0 15056 1735 15058
rect 0 15000 1674 15056
rect 1730 15000 1735 15056
rect 0 14998 1735 15000
rect 0 14968 480 14998
rect 1669 14995 1735 14998
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 1669 14650 1735 14653
rect 0 14648 1735 14650
rect 0 14592 1674 14648
rect 1730 14592 1735 14648
rect 0 14590 1735 14592
rect 0 14560 480 14590
rect 1669 14587 1735 14590
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 3417 14106 3483 14109
rect 0 14104 3483 14106
rect 0 14048 3422 14104
rect 3478 14048 3483 14104
rect 0 14046 3483 14048
rect 0 14016 480 14046
rect 3417 14043 3483 14046
rect 0 13698 480 13728
rect 3509 13698 3575 13701
rect 0 13696 3575 13698
rect 0 13640 3514 13696
rect 3570 13640 3575 13696
rect 0 13638 3575 13640
rect 0 13608 480 13638
rect 3509 13635 3575 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 0 13290 480 13320
rect 1669 13290 1735 13293
rect 0 13288 1735 13290
rect 0 13232 1674 13288
rect 1730 13232 1735 13288
rect 0 13230 1735 13232
rect 0 13200 480 13230
rect 1669 13227 1735 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12746 480 12776
rect 8293 12746 8359 12749
rect 0 12744 8359 12746
rect 0 12688 8298 12744
rect 8354 12688 8359 12744
rect 0 12686 8359 12688
rect 0 12656 480 12686
rect 8293 12683 8359 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 9121 12338 9187 12341
rect 0 12336 9187 12338
rect 0 12280 9126 12336
rect 9182 12280 9187 12336
rect 0 12278 9187 12280
rect 0 12248 480 12278
rect 9121 12275 9187 12278
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 480 11824
rect 8661 11794 8727 11797
rect 0 11792 8727 11794
rect 0 11736 8666 11792
rect 8722 11736 8727 11792
rect 0 11734 8727 11736
rect 0 11704 480 11734
rect 8661 11731 8727 11734
rect 4061 11522 4127 11525
rect 7097 11522 7163 11525
rect 4061 11520 7163 11522
rect 4061 11464 4066 11520
rect 4122 11464 7102 11520
rect 7158 11464 7163 11520
rect 4061 11462 7163 11464
rect 4061 11459 4127 11462
rect 7097 11459 7163 11462
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 4061 11386 4127 11389
rect 0 11384 4127 11386
rect 0 11328 4066 11384
rect 4122 11328 4127 11384
rect 0 11326 4127 11328
rect 0 11296 480 11326
rect 4061 11323 4127 11326
rect 9673 11250 9739 11253
rect 18597 11250 18663 11253
rect 9673 11248 18663 11250
rect 9673 11192 9678 11248
rect 9734 11192 18602 11248
rect 18658 11192 18663 11248
rect 9673 11190 18663 11192
rect 9673 11187 9739 11190
rect 18597 11187 18663 11190
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 3877 10842 3943 10845
rect 0 10840 3943 10842
rect 0 10784 3882 10840
rect 3938 10784 3943 10840
rect 0 10782 3943 10784
rect 0 10752 480 10782
rect 3877 10779 3943 10782
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 0 10026 480 10056
rect 3141 10026 3207 10029
rect 0 10024 3207 10026
rect 0 9968 3146 10024
rect 3202 9968 3207 10024
rect 0 9966 3207 9968
rect 0 9936 480 9966
rect 3141 9963 3207 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 4521 9618 4587 9621
rect 5533 9618 5599 9621
rect 4521 9616 5599 9618
rect 4521 9560 4526 9616
rect 4582 9560 5538 9616
rect 5594 9560 5599 9616
rect 4521 9558 5599 9560
rect 4521 9555 4587 9558
rect 5533 9555 5599 9558
rect 0 9482 480 9512
rect 8845 9482 8911 9485
rect 0 9480 8911 9482
rect 0 9424 8850 9480
rect 8906 9424 8911 9480
rect 0 9422 8911 9424
rect 0 9392 480 9422
rect 8845 9419 8911 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 7833 9074 7899 9077
rect 0 9072 7899 9074
rect 0 9016 7838 9072
rect 7894 9016 7899 9072
rect 0 9014 7899 9016
rect 0 8984 480 9014
rect 7833 9011 7899 9014
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 480 8560
rect 4061 8530 4127 8533
rect 0 8528 4127 8530
rect 0 8472 4066 8528
rect 4122 8472 4127 8528
rect 0 8470 4127 8472
rect 0 8440 480 8470
rect 4061 8467 4127 8470
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 480 8062
rect 4061 8059 4127 8062
rect 3049 7850 3115 7853
rect 4521 7850 4587 7853
rect 3049 7848 4587 7850
rect 3049 7792 3054 7848
rect 3110 7792 4526 7848
rect 4582 7792 4587 7848
rect 3049 7790 4587 7792
rect 3049 7787 3115 7790
rect 4521 7787 4587 7790
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 3325 7578 3391 7581
rect 0 7576 3391 7578
rect 0 7520 3330 7576
rect 3386 7520 3391 7576
rect 0 7518 3391 7520
rect 0 7488 480 7518
rect 3325 7515 3391 7518
rect 0 7170 480 7200
rect 3969 7170 4035 7173
rect 0 7168 4035 7170
rect 0 7112 3974 7168
rect 4030 7112 4035 7168
rect 0 7110 4035 7112
rect 0 7080 480 7110
rect 3969 7107 4035 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 0 6762 480 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 480 6702
rect 4061 6699 4127 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 11697 6354 11763 6357
rect 14549 6354 14615 6357
rect 11697 6352 14615 6354
rect 11697 6296 11702 6352
rect 11758 6296 14554 6352
rect 14610 6296 14615 6352
rect 11697 6294 14615 6296
rect 11697 6291 11763 6294
rect 14549 6291 14615 6294
rect 0 6218 480 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 480 6158
rect 4061 6155 4127 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 480 5750
rect 4061 5747 4127 5750
rect 9857 5810 9923 5813
rect 15285 5810 15351 5813
rect 9857 5808 15351 5810
rect 9857 5752 9862 5808
rect 9918 5752 15290 5808
rect 15346 5752 15351 5808
rect 9857 5750 15351 5752
rect 9857 5747 9923 5750
rect 15285 5747 15351 5750
rect 18597 5810 18663 5813
rect 22320 5810 22800 5840
rect 18597 5808 22800 5810
rect 18597 5752 18602 5808
rect 18658 5752 22800 5808
rect 18597 5750 22800 5752
rect 18597 5747 18663 5750
rect 22320 5720 22800 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 3693 5266 3759 5269
rect 0 5264 3759 5266
rect 0 5208 3698 5264
rect 3754 5208 3759 5264
rect 0 5206 3759 5208
rect 0 5176 480 5206
rect 3693 5203 3759 5206
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 2221 4858 2287 4861
rect 0 4856 2287 4858
rect 0 4800 2226 4856
rect 2282 4800 2287 4856
rect 0 4798 2287 4800
rect 0 4768 480 4798
rect 2221 4795 2287 4798
rect 9857 4858 9923 4861
rect 14365 4858 14431 4861
rect 9857 4856 14431 4858
rect 9857 4800 9862 4856
rect 9918 4800 14370 4856
rect 14426 4800 14431 4856
rect 9857 4798 14431 4800
rect 9857 4795 9923 4798
rect 14365 4795 14431 4798
rect 6729 4722 6795 4725
rect 9489 4722 9555 4725
rect 6729 4720 9555 4722
rect 6729 4664 6734 4720
rect 6790 4664 9494 4720
rect 9550 4664 9555 4720
rect 6729 4662 9555 4664
rect 6729 4659 6795 4662
rect 9489 4659 9555 4662
rect 4705 4586 4771 4589
rect 8293 4586 8359 4589
rect 9213 4586 9279 4589
rect 4705 4584 9279 4586
rect 4705 4528 4710 4584
rect 4766 4528 8298 4584
rect 8354 4528 9218 4584
rect 9274 4528 9279 4584
rect 4705 4526 9279 4528
rect 4705 4523 4771 4526
rect 8293 4523 8359 4526
rect 9213 4523 9279 4526
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 4061 4314 4127 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 0 4224 480 4254
rect 4061 4251 4127 4254
rect 13353 4042 13419 4045
rect 15009 4042 15075 4045
rect 13353 4040 15075 4042
rect 13353 3984 13358 4040
rect 13414 3984 15014 4040
rect 15070 3984 15075 4040
rect 13353 3982 15075 3984
rect 13353 3979 13419 3982
rect 15009 3979 15075 3982
rect 0 3906 480 3936
rect 2957 3906 3023 3909
rect 0 3904 3023 3906
rect 0 3848 2962 3904
rect 3018 3848 3023 3904
rect 0 3846 3023 3848
rect 0 3816 480 3846
rect 2957 3843 3023 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 3141 3634 3207 3637
rect 6729 3634 6795 3637
rect 3141 3632 6795 3634
rect 3141 3576 3146 3632
rect 3202 3576 6734 3632
rect 6790 3576 6795 3632
rect 3141 3574 6795 3576
rect 3141 3571 3207 3574
rect 6729 3571 6795 3574
rect 0 3498 480 3528
rect 2129 3498 2195 3501
rect 0 3496 2195 3498
rect 0 3440 2134 3496
rect 2190 3440 2195 3496
rect 0 3438 2195 3440
rect 0 3408 480 3438
rect 2129 3435 2195 3438
rect 2221 3362 2287 3365
rect 3877 3362 3943 3365
rect 2221 3360 3943 3362
rect 2221 3304 2226 3360
rect 2282 3304 3882 3360
rect 3938 3304 3943 3360
rect 2221 3302 3943 3304
rect 2221 3299 2287 3302
rect 3877 3299 3943 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 480 2984
rect 1577 2954 1643 2957
rect 0 2952 1643 2954
rect 0 2896 1582 2952
rect 1638 2896 1643 2952
rect 0 2894 1643 2896
rect 0 2864 480 2894
rect 1577 2891 1643 2894
rect 3417 2954 3483 2957
rect 10133 2954 10199 2957
rect 3417 2952 10199 2954
rect 3417 2896 3422 2952
rect 3478 2896 10138 2952
rect 10194 2896 10199 2952
rect 3417 2894 10199 2896
rect 3417 2891 3483 2894
rect 10133 2891 10199 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 3049 2546 3115 2549
rect 0 2544 3115 2546
rect 0 2488 3054 2544
rect 3110 2488 3115 2544
rect 0 2486 3115 2488
rect 0 2456 480 2486
rect 3049 2483 3115 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 3969 2002 4035 2005
rect 0 2000 4035 2002
rect 0 1944 3974 2000
rect 4030 1944 4035 2000
rect 0 1942 4035 1944
rect 0 1912 480 1942
rect 3969 1939 4035 1942
rect 0 1594 480 1624
rect 3601 1594 3667 1597
rect 0 1592 3667 1594
rect 0 1536 3606 1592
rect 3662 1536 3667 1592
rect 0 1534 3667 1536
rect 0 1504 480 1534
rect 3601 1531 3667 1534
rect 0 1050 480 1080
rect 3509 1050 3575 1053
rect 0 1048 3575 1050
rect 0 992 3514 1048
rect 3570 992 3575 1048
rect 0 990 3575 992
rect 0 960 480 990
rect 3509 987 3575 990
rect 0 642 480 672
rect 1301 642 1367 645
rect 0 640 1367 642
rect 0 584 1306 640
rect 1362 584 1367 640
rect 0 582 1367 584
rect 0 552 480 582
rect 1301 579 1367 582
rect 0 234 480 264
rect 3785 234 3851 237
rect 0 232 3851 234
rect 0 176 3790 232
rect 3846 176 3851 232
rect 0 174 3851 176
rect 0 144 480 174
rect 3785 171 3851 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2116 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1932 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 3864 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1606256979
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40
timestamp 1606256979
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp 1606256979
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4968 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51
timestamp 1606256979
transform 1 0 5796 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1606256979
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606256979
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7268 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp 1606256979
transform 1 0 7728 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1606256979
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _057_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9936 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8924 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_84
timestamp 1606256979
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1606256979
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1606256979
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94
timestamp 1606256979
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1606256979
transform 1 0 10764 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_111
timestamp 1606256979
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10764 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _110_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11500 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606256979
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606256979
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1606256979
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1606256979
transform 1 0 12052 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_133
timestamp 1606256979
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1606256979
transform 1 0 12972 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1606256979
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13432 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606256979
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1606256979
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1606256979
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1606256979
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606256979
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606256979
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606256979
transform 1 0 14444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_149
timestamp 1606256979
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1606256979
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14996 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606256979
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_157
timestamp 1606256979
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1606256979
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15732 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_165
timestamp 1606256979
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_166
timestamp 1606256979
transform 1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1606256979
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606256979
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_177
timestamp 1606256979
transform 1 0 17388 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_171
timestamp 1606256979
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606256979
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606256979
transform 1 0 17020 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606256979
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1606256979
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_173
timestamp 1606256979
transform 1 0 17020 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606256979
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1606256979
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp 1606256979
transform 1 0 20240 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606256979
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606256979
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606256979
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1606256979
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1606256979
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1564 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4508 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_21
timestamp 1606256979
transform 1 0 3036 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1606256979
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_35
timestamp 1606256979
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 6348 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1606256979
transform 1 0 5980 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7728 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_2_66
timestamp 1606256979
transform 1 0 7176 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9844 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1606256979
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_104
timestamp 1606256979
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10856 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12512 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_122
timestamp 1606256979
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14352 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_140
timestamp 1606256979
transform 1 0 13984 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15456 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1606256979
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_165
timestamp 1606256979
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1606256979
transform 1 0 18308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606256979
transform 1 0 17756 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606256979
transform 1 0 17204 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16468 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1606256979
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_179
timestamp 1606256979
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_185
timestamp 1606256979
transform 1 0 18124 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606256979
transform 1 0 19964 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1606256979
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_202
timestamp 1606256979
transform 1 0 19688 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1606256979
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1606256979
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606256979
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606256979
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2944 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1932 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1606256979
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_36
timestamp 1606256979
transform 1 0 4416 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5060 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_42
timestamp 1606256979
transform 1 0 4968 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606256979
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7728 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_65
timestamp 1606256979
transform 1 0 7084 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_71
timestamp 1606256979
transform 1 0 7636 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1606256979
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9752 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1606256979
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11408 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12604 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1606256979
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1606256979
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13340 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1606256979
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 14996 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1606256979
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16652 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_167
timestamp 1606256979
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1606256979
transform 1 0 17480 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1606256979
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1606256979
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1606256979
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1840 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_6
timestamp 1606256979
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4508 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_24
timestamp 1606256979
transform 1 0 3312 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1606256979
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1606256979
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5520 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6532 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_46
timestamp 1606256979
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_57
timestamp 1606256979
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7820 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1606256979
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_72
timestamp 1606256979
transform 1 0 7728 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_82
timestamp 1606256979
transform 1 0 8648 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1606256979
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1606256979
transform 1 0 11316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12420 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_109
timestamp 1606256979
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_114
timestamp 1606256979
transform 1 0 11592 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_122
timestamp 1606256979
transform 1 0 12328 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13708 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_129
timestamp 1606256979
transform 1 0 12972 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15456 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_146
timestamp 1606256979
transform 1 0 14536 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1606256979
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18032 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17112 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_172
timestamp 1606256979
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1606256979
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_200
timestamp 1606256979
transform 1 0 19504 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606256979
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606256979
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606256979
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 2760 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1748 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_16
timestamp 1606256979
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4232 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_27
timestamp 1606256979
transform 1 0 3588 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_33
timestamp 1606256979
transform 1 0 4140 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_43
timestamp 1606256979
transform 1 0 5060 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_49
timestamp 1606256979
transform 1 0 5612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8740 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1606256979
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1606256979
transform 1 0 8648 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_99
timestamp 1606256979
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606256979
transform 1 0 11868 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_110
timestamp 1606256979
transform 1 0 11224 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_116
timestamp 1606256979
transform 1 0 11776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606256979
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13616 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14352 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1606256979
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_142
timestamp 1606256979
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15180 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_150
timestamp 1606256979
transform 1 0 14904 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1606256979
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1606256979
transform 1 0 17204 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_173
timestamp 1606256979
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1606256979
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1606256979
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1606256979
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1606256979
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 2484 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1472 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_13
timestamp 1606256979
transform 1 0 2300 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1606256979
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606256979
transform 1 0 3036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 3588 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_24
timestamp 1606256979
transform 1 0 3312 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1606256979
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_41
timestamp 1606256979
transform 1 0 4876 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp 1606256979
transform 1 0 3312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5520 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5612 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_47
timestamp 1606256979
transform 1 0 5428 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_43
timestamp 1606256979
transform 1 0 5060 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1606256979
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8188 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1606256979
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_75
timestamp 1606256979
transform 1 0 8004 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_71
timestamp 1606256979
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10488 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10212 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1606256979
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_96
timestamp 1606256979
transform 1 0 9936 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_93
timestamp 1606256979
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_104
timestamp 1606256979
transform 1 0 10672 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12144 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12512 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11040 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_118
timestamp 1606256979
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1606256979
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1606256979
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13800 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_136
timestamp 1606256979
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1606256979
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1606256979
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1606256979
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_147
timestamp 1606256979
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15180 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_162
timestamp 1606256979
transform 1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_160
timestamp 1606256979
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16284 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16008 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606256979
transform 1 0 17664 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1606256979
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1606256979
transform 1 0 18032 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606256979
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1606256979
transform 1 0 19136 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1606256979
transform 1 0 20240 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1606256979
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1606256979
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606256979
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606256979
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1932 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_25
timestamp 1606256979
transform 1 0 3404 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 1606256979
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5428 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 5152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7084 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_63
timestamp 1606256979
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_81
timestamp 1606256979
transform 1 0 8556 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9936 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1606256979
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1606256979
transform 1 0 12604 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10948 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1606256979
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_123
timestamp 1606256979
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13064 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1606256979
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_146
timestamp 1606256979
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1606256979
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16928 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1606256979
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1606256979
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1606256979
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1606256979
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606256979
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606256979
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2944 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1932 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_18
timestamp 1606256979
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4416 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_29
timestamp 1606256979
transform 1 0 3772 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_35
timestamp 1606256979
transform 1 0 4324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1606256979
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1606256979
transform 1 0 5888 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606256979
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8096 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_71
timestamp 1606256979
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_75
timestamp 1606256979
transform 1 0 8004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10304 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_85
timestamp 1606256979
transform 1 0 8924 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_97
timestamp 1606256979
transform 1 0 10028 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 11960 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_116
timestamp 1606256979
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1606256979
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1606256979
transform 1 0 13616 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14260 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_135
timestamp 1606256979
transform 1 0 13524 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1606256979
transform 1 0 13892 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1606256979
transform 1 0 15548 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_152
timestamp 1606256979
transform 1 0 15088 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_156
timestamp 1606256979
transform 1 0 15456 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_160
timestamp 1606256979
transform 1 0 15824 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16928 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1606256979
transform 1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1606256979
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1606256979
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1606256979
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 2208 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1606256979
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1606256979
transform 1 0 3036 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1606256979
transform 1 0 3588 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp 1606256979
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5152 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_60
timestamp 1606256979
transform 1 0 6624 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 6900 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7912 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1606256979
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_83
timestamp 1606256979
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10120 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1606256979
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp 1606256979
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11132 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1606256979
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_118
timestamp 1606256979
transform 1 0 11960 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_130
timestamp 1606256979
transform 1 0 13064 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_142
timestamp 1606256979
transform 1 0 14168 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1606256979
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_170
timestamp 1606256979
transform 1 0 16744 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_182
timestamp 1606256979
transform 1 0 17848 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_194
timestamp 1606256979
transform 1 0 18952 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_206
timestamp 1606256979
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606256979
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606256979
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2760 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1748 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1606256979
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4416 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1606256979
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_45
timestamp 1606256979
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606256979
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7268 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_65
timestamp 1606256979
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_83
timestamp 1606256979
transform 1 0 8740 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9568 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 9200 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 1606256979
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_91
timestamp 1606256979
transform 1 0 9476 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 11224 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_108
timestamp 1606256979
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1606256979
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1606256979
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1606256979
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1606256979
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1606256979
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1606256979
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1606256979
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1606256979
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1606256979
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606256979
transform 1 0 3036 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1606256979
transform 1 0 3496 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_24
timestamp 1606256979
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606256979
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1606256979
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1606256979
transform 1 0 6072 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1606256979
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8096 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 7084 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1606256979
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_71
timestamp 1606256979
transform 1 0 7636 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_75
timestamp 1606256979
transform 1 0 8004 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9844 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1606256979
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1606256979
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_111
timestamp 1606256979
transform 1 0 11316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1606256979
transform 1 0 12420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_135
timestamp 1606256979
transform 1 0 13524 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_147
timestamp 1606256979
transform 1 0 14628 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1606256979
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1606256979
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1606256979
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1606256979
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606256979
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606256979
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1564 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_15
timestamp 1606256979
transform 1 0 2484 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4324 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 3496 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1606256979
transform 1 0 3036 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_25
timestamp 1606256979
transform 1 0 3404 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606256979
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_32
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1606256979
transform 1 0 5796 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_42
timestamp 1606256979
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_59
timestamp 1606256979
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606256979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1606256979
transform 1 0 5980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606256979
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7820 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1606256979
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1606256979
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_78
timestamp 1606256979
transform 1 0 8280 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8832 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9844 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606256979
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_109
timestamp 1606256979
transform 1 0 11132 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1606256979
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_115
timestamp 1606256979
transform 1 0 11684 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1606256979
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_127
timestamp 1606256979
transform 1 0 12788 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_139
timestamp 1606256979
transform 1 0 13892 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1606256979
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1606256979
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606256979
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1606256979
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1606256979
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1606256979
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1606256979
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1606256979
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1606256979
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1606256979
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606256979
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606256979
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1564 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_21
timestamp 1606256979
transform 1 0 3036 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1606256979
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_37
timestamp 1606256979
transform 1 0 4508 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5060 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606256979
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7728 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_69
timestamp 1606256979
transform 1 0 7452 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606256979
transform 1 0 10396 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9384 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_88
timestamp 1606256979
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1606256979
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_104
timestamp 1606256979
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 10856 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_109
timestamp 1606256979
transform 1 0 11132 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1606256979
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1606256979
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1606256979
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1606256979
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606256979
transform 1 0 18216 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1606256979
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_190
timestamp 1606256979
transform 1 0 18584 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_202
timestamp 1606256979
transform 1 0 19688 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_214
timestamp 1606256979
transform 1 0 20792 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_12
timestamp 1606256979
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4416 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1606256979
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606256979
transform 1 0 6440 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5428 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp 1606256979
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_56
timestamp 1606256979
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_61
timestamp 1606256979
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6900 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_72
timestamp 1606256979
transform 1 0 7728 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_80
timestamp 1606256979
transform 1 0 8464 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606256979
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1606256979
transform 1 0 11132 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1606256979
transform 1 0 12236 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_133
timestamp 1606256979
transform 1 0 13340 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1606256979
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1606256979
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1606256979
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606256979
transform 1 0 18584 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_194
timestamp 1606256979
transform 1 0 18952 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1606256979
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606256979
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606256979
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2024 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1606256979
transform 1 0 1932 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 3680 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_26
timestamp 1606256979
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_37
timestamp 1606256979
transform 1 0 4508 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5060 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606256979
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606256979
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7636 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 6992 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_67
timestamp 1606256979
transform 1 0 7268 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_80
timestamp 1606256979
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9292 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1606256979
transform 1 0 8924 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_105
timestamp 1606256979
transform 1 0 10764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1606256979
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606256979
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1606256979
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1606256979
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1606256979
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1606256979
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_184
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606256979
transform 1 0 19044 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_192
timestamp 1606256979
transform 1 0 18768 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_199
timestamp 1606256979
transform 1 0 19412 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_211
timestamp 1606256979
transform 1 0 20516 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 1606256979
transform 1 0 21252 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606256979
transform 1 0 1472 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2024 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_8
timestamp 1606256979
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_19
timestamp 1606256979
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606256979
transform 1 0 3036 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4508 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_24
timestamp 1606256979
transform 1 0 3312 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1606256979
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5520 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1606256979
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7268 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_64
timestamp 1606256979
transform 1 0 6992 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_83
timestamp 1606256979
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1606256979
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_102
timestamp 1606256979
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_114
timestamp 1606256979
transform 1 0 11592 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_126
timestamp 1606256979
transform 1 0 12696 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_138
timestamp 1606256979
transform 1 0 13800 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1606256979
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1606256979
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1606256979
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606256979
transform 1 0 19504 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_190
timestamp 1606256979
transform 1 0 18584 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1606256979
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_204
timestamp 1606256979
transform 1 0 19872 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606256979
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1606256979
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1606256979
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1606256979
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1840 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1748 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_14
timestamp 1606256979
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_13
timestamp 1606256979
transform 1 0 2300 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2576 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2852 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606256979
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4600 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_35
timestamp 1606256979
transform 1 0 4324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_22
timestamp 1606256979
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1606256979
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606256979
transform 1 0 6256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5704 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1606256979
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606256979
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1606256979
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_59
timestamp 1606256979
transform 1 0 6532 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606256979
transform 1 0 7176 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7636 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7544 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 7084 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1606256979
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_68
timestamp 1606256979
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1606256979
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 10028 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_87
timestamp 1606256979
transform 1 0 9108 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1606256979
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_100
timestamp 1606256979
transform 1 0 10304 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1606256979
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_102
timestamp 1606256979
transform 1 0 10488 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_112
timestamp 1606256979
transform 1 0 11408 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1606256979
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_114
timestamp 1606256979
transform 1 0 11592 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1606256979
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_126
timestamp 1606256979
transform 1 0 12696 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_138
timestamp 1606256979
transform 1 0 13800 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1606256979
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1606256979
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1606256979
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1606256979
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1606256979
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1606256979
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1606256979
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1606256979
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1606256979
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1606256979
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606256979
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606256979
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1748 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2484 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_13
timestamp 1606256979
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606256979
transform 1 0 3772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606256979
transform 1 0 3220 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4232 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1606256979
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_27
timestamp 1606256979
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_32
timestamp 1606256979
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606256979
transform 1 0 5888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_50
timestamp 1606256979
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_55
timestamp 1606256979
transform 1 0 6164 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8556 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_78
timestamp 1606256979
transform 1 0 8280 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606256979
transform 1 0 10212 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1606256979
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_102
timestamp 1606256979
transform 1 0 10488 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1606256979
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1606256979
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1606256979
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1606256979
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1606256979
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1606256979
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1606256979
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606256979
transform 1 0 1472 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2024 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_8
timestamp 1606256979
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4416 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_26
timestamp 1606256979
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1606256979
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606256979
transform 1 0 5888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6348 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_45
timestamp 1606256979
transform 1 0 5244 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_51
timestamp 1606256979
transform 1 0 5796 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1606256979
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1606256979
transform 1 0 7820 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1606256979
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1606256979
transform 1 0 11132 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1606256979
transform 1 0 12236 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_133
timestamp 1606256979
transform 1 0 13340 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1606256979
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1606256979
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1606256979
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1606256979
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1606256979
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606256979
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606256979
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606256979
transform 1 0 1472 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2760 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2024 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_8
timestamp 1606256979
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_16
timestamp 1606256979
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4600 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1606256979
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 1606256979
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606256979
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6992 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8004 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606256979
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9200 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606256979
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_86
timestamp 1606256979
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_104
timestamp 1606256979
transform 1 0 10672 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_116
timestamp 1606256979
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1606256979
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1606256979
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1606256979
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1606256979
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1606256979
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1606256979
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1606256979
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606256979
transform 1 0 1472 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2024 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_8
timestamp 1606256979
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_16
timestamp 1606256979
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4232 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606256979
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5888 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1606256979
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_45
timestamp 1606256979
transform 1 0 5244 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_51
timestamp 1606256979
transform 1 0 5796 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7544 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1606256979
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606256979
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_86
timestamp 1606256979
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_104
timestamp 1606256979
transform 1 0 10672 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10948 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606256979
transform 1 0 11776 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_118
timestamp 1606256979
transform 1 0 11960 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_130
timestamp 1606256979
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_142
timestamp 1606256979
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1606256979
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1606256979
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1606256979
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1606256979
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1606256979
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606256979
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606256979
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606256979
transform 1 0 2760 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606256979
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2024 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1606256979
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1606256979
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 3496 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_22
timestamp 1606256979
transform 1 0 3128 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606256979
transform 1 0 6164 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_42
timestamp 1606256979
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1606256979
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1606256979
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8188 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7176 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_75
timestamp 1606256979
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10120 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1606256979
transform 1 0 9660 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_97
timestamp 1606256979
transform 1 0 10028 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_114
timestamp 1606256979
transform 1 0 11592 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1606256979
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1606256979
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1606256979
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1606256979
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606256979
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1606256979
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1606256979
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1656 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606256979
transform 1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1606256979
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_12
timestamp 1606256979
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2116 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1606256979
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_20
timestamp 1606256979
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2852 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2392 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606256979
transform 1 0 3956 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606256979
transform 1 0 3128 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4324 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_26
timestamp 1606256979
transform 1 0 3496 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1606256979
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_32
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_25
timestamp 1606256979
transform 1 0 3404 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_34
timestamp 1606256979
transform 1 0 4232 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5980 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5520 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_51
timestamp 1606256979
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_46
timestamp 1606256979
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1606256979
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606256979
transform 1 0 7912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8372 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1606256979
transform 1 0 7452 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_73
timestamp 1606256979
transform 1 0 7820 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_77
timestamp 1606256979
transform 1 0 8188 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_74
timestamp 1606256979
transform 1 0 7912 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_78
timestamp 1606256979
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606256979
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9108 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1606256979
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1606256979
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1606256979
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_96
timestamp 1606256979
transform 1 0 9936 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606256979
transform 1 0 11684 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11316 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1606256979
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1606256979
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1606256979
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_127
timestamp 1606256979
transform 1 0 12788 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_139
timestamp 1606256979
transform 1 0 13892 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1606256979
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1606256979
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1606256979
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1606256979
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1606256979
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1606256979
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1606256979
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1606256979
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1606256979
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1606256979
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1606256979
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1606256979
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606256979
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606256979
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606256979
transform 1 0 2944 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606256979
transform 1 0 1656 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2208 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1606256979
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1606256979
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_18
timestamp 1606256979
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_24
timestamp 1606256979
transform 1 0 3312 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1606256979
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606256979
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606256979
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606256979
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 7728 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1606256979
transform 1 0 7360 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_78
timestamp 1606256979
transform 1 0 8280 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 10028 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606256979
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1606256979
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_103
timestamp 1606256979
transform 1 0 10580 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_115
timestamp 1606256979
transform 1 0 11684 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_127
timestamp 1606256979
transform 1 0 12788 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_139
timestamp 1606256979
transform 1 0 13892 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1606256979
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1606256979
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1606256979
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1606256979
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1606256979
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1606256979
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606256979
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606256979
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606256979
transform 1 0 2852 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606256979
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606256979
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1606256979
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1606256979
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1606256979
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1606256979
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_47
timestamp 1606256979
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606256979
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1606256979
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 6992 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1606256979
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1606256979
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1606256979
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_106
timestamp 1606256979
transform 1 0 10856 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1606256979
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1606256979
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1606256979
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1606256979
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1606256979
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1606256979
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606256979
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1606256979
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1606256979
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2116 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2852 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1606256979
transform 1 0 1380 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1606256979
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_25
timestamp 1606256979
transform 1 0 3404 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606256979
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1606256979
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_56
timestamp 1606256979
transform 1 0 6256 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606256979
transform 1 0 7268 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_64
timestamp 1606256979
transform 1 0 6992 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_71
timestamp 1606256979
transform 1 0 7636 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_83
timestamp 1606256979
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1606256979
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1606256979
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1606256979
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1606256979
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1606256979
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1606256979
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1606256979
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1606256979
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1606256979
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1606256979
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1606256979
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606256979
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606256979
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606256979
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1606256979
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1606256979
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_17
timestamp 1606256979
transform 1 0 2668 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1606256979
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_41
timestamp 1606256979
transform 1 0 4876 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606256979
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1606256979
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_66
timestamp 1606256979
transform 1 0 7176 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_78
timestamp 1606256979
transform 1 0 8280 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_90
timestamp 1606256979
transform 1 0 9384 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_102
timestamp 1606256979
transform 1 0 10488 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_114
timestamp 1606256979
transform 1 0 11592 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1606256979
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1606256979
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1606256979
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1606256979
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1606256979
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1606256979
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1606256979
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1606256979
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606256979
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1606256979
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1606256979
transform 1 0 2116 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1606256979
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606256979
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606256979
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606256979
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606256979
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1606256979
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606256979
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1606256979
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1606256979
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1606256979
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1606256979
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1606256979
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1606256979
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1606256979
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1606256979
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1606256979
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1606256979
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1606256979
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1606256979
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606256979
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 21638 0 21694 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 22098 0 22154 480 6 SC_OUT_BOT
port 1 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 2 nsew default input
rlabel metal2 s 570 0 626 480 6 bottom_left_grid_pin_43_
port 3 nsew default input
rlabel metal2 s 1030 0 1086 480 6 bottom_left_grid_pin_44_
port 4 nsew default input
rlabel metal2 s 1490 0 1546 480 6 bottom_left_grid_pin_45_
port 5 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_46_
port 6 nsew default input
rlabel metal2 s 2318 0 2374 480 6 bottom_left_grid_pin_47_
port 7 nsew default input
rlabel metal2 s 2778 0 2834 480 6 bottom_left_grid_pin_48_
port 8 nsew default input
rlabel metal2 s 3238 0 3294 480 6 bottom_left_grid_pin_49_
port 9 nsew default input
rlabel metal2 s 21178 0 21234 480 6 bottom_right_grid_pin_1_
port 10 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 ccff_head
port 11 nsew default input
rlabel metal3 s 22320 17144 22800 17264 6 ccff_tail
port 12 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 13 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[10]
port 14 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[11]
port 15 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[12]
port 16 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[13]
port 17 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[14]
port 18 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[15]
port 19 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[16]
port 20 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[17]
port 21 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[18]
port 22 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[19]
port 23 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[1]
port 24 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[2]
port 25 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[3]
port 26 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[4]
port 27 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[5]
port 28 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[6]
port 29 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[7]
port 30 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 31 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[9]
port 32 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[0]
port 33 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[10]
port 34 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[11]
port 35 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[12]
port 36 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[13]
port 37 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[14]
port 38 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[15]
port 39 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[16]
port 40 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[17]
port 41 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[18]
port 42 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[19]
port 43 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[1]
port 44 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[2]
port 45 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[3]
port 46 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[4]
port 47 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[5]
port 48 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[6]
port 49 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[7]
port 50 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[8]
port 51 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[9]
port 52 nsew default tristate
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[0]
port 53 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[10]
port 54 nsew default input
rlabel metal2 s 8482 0 8538 480 6 chany_bottom_in[11]
port 55 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[12]
port 56 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[13]
port 57 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[14]
port 58 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[15]
port 59 nsew default input
rlabel metal2 s 10690 0 10746 480 6 chany_bottom_in[16]
port 60 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[17]
port 61 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[18]
port 62 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[19]
port 63 nsew default input
rlabel metal2 s 4066 0 4122 480 6 chany_bottom_in[1]
port 64 nsew default input
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[2]
port 65 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[3]
port 66 nsew default input
rlabel metal2 s 5446 0 5502 480 6 chany_bottom_in[4]
port 67 nsew default input
rlabel metal2 s 5906 0 5962 480 6 chany_bottom_in[5]
port 68 nsew default input
rlabel metal2 s 6274 0 6330 480 6 chany_bottom_in[6]
port 69 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[7]
port 70 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[8]
port 71 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[9]
port 72 nsew default input
rlabel metal2 s 12438 0 12494 480 6 chany_bottom_out[0]
port 73 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chany_bottom_out[10]
port 74 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[11]
port 75 nsew default tristate
rlabel metal2 s 17682 0 17738 480 6 chany_bottom_out[12]
port 76 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 chany_bottom_out[13]
port 77 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[14]
port 78 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[15]
port 79 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 chany_bottom_out[16]
port 80 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[17]
port 81 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_out[18]
port 82 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[19]
port 83 nsew default tristate
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_out[1]
port 84 nsew default tristate
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_out[2]
port 85 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[3]
port 86 nsew default tristate
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_out[4]
port 87 nsew default tristate
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_out[5]
port 88 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_out[6]
port 89 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[7]
port 90 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[8]
port 91 nsew default tristate
rlabel metal2 s 16394 0 16450 480 6 chany_bottom_out[9]
port 92 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 93 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 94 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_36_
port 95 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 96 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_38_
port 97 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 98 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_40_
port 99 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 100 nsew default input
rlabel metal3 s 0 22448 480 22568 6 left_top_grid_pin_1_
port 101 nsew default input
rlabel metal2 s 22558 0 22614 480 6 prog_clk_0_S_in
port 102 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 103 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 104 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22568
<< end >>
