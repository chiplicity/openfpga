magic
tech EFS8A
magscale 1 2
timestamp 1604399152
<< locali >>
rect 22017 16983 22051 17221
rect 14933 10523 14967 10693
rect 15393 10523 15427 10761
rect 15209 6239 15243 6409
rect 22845 5083 22879 5185
rect 17693 4063 17727 4165
rect 22569 3451 22603 3621
<< viali >>
rect 14473 25449 14507 25483
rect 15669 25449 15703 25483
rect 16865 25449 16899 25483
rect 19625 25449 19659 25483
rect 22201 25449 22235 25483
rect 14289 25313 14323 25347
rect 15485 25313 15519 25347
rect 16681 25313 16715 25347
rect 19441 25313 19475 25347
rect 22017 25313 22051 25347
rect 18153 25245 18187 25279
rect 18337 25245 18371 25279
rect 16129 25109 16163 25143
rect 22017 24837 22051 24871
rect 15945 24769 15979 24803
rect 16129 24769 16163 24803
rect 17509 24769 17543 24803
rect 18705 24769 18739 24803
rect 12817 24701 12851 24735
rect 13921 24701 13955 24735
rect 14381 24701 14415 24735
rect 15025 24701 15059 24735
rect 15853 24701 15887 24735
rect 18429 24701 18463 24735
rect 19993 24701 20027 24735
rect 20545 24701 20579 24735
rect 21097 24701 21131 24735
rect 21649 24701 21683 24735
rect 22201 24701 22235 24735
rect 22753 24701 22787 24735
rect 15393 24633 15427 24667
rect 17877 24633 17911 24667
rect 18521 24633 18555 24667
rect 13001 24565 13035 24599
rect 13369 24565 13403 24599
rect 14289 24565 14323 24599
rect 14565 24565 14599 24599
rect 15485 24565 15519 24599
rect 16773 24565 16807 24599
rect 18061 24565 18095 24599
rect 19441 24565 19475 24599
rect 20177 24565 20211 24599
rect 21281 24565 21315 24599
rect 22385 24565 22419 24599
rect 12357 24361 12391 24395
rect 16313 24361 16347 24395
rect 19809 24361 19843 24395
rect 23673 24361 23707 24395
rect 24777 24361 24811 24395
rect 12265 24225 12299 24259
rect 13369 24225 13403 24259
rect 13829 24225 13863 24259
rect 13921 24225 13955 24259
rect 15485 24225 15519 24259
rect 16221 24225 16255 24259
rect 17325 24225 17359 24259
rect 18153 24225 18187 24259
rect 19625 24225 19659 24259
rect 21281 24225 21315 24259
rect 23489 24225 23523 24259
rect 24593 24225 24627 24259
rect 12541 24157 12575 24191
rect 14013 24157 14047 24191
rect 16405 24157 16439 24191
rect 18245 24157 18279 24191
rect 18429 24157 18463 24191
rect 21373 24157 21407 24191
rect 21557 24157 21591 24191
rect 22477 24157 22511 24191
rect 13001 24089 13035 24123
rect 15853 24089 15887 24123
rect 17601 24089 17635 24123
rect 11897 24021 11931 24055
rect 13461 24021 13495 24055
rect 14933 24021 14967 24055
rect 17785 24021 17819 24055
rect 18981 24021 19015 24055
rect 20913 24021 20947 24055
rect 11529 23817 11563 23851
rect 11989 23817 12023 23851
rect 14933 23817 14967 23851
rect 16037 23817 16071 23851
rect 16313 23817 16347 23851
rect 17049 23817 17083 23851
rect 21281 23817 21315 23851
rect 22661 23817 22695 23851
rect 24777 23817 24811 23851
rect 15577 23681 15611 23715
rect 25145 23681 25179 23715
rect 12449 23613 12483 23647
rect 12716 23613 12750 23647
rect 16865 23613 16899 23647
rect 18981 23613 19015 23647
rect 22477 23613 22511 23647
rect 24593 23613 24627 23647
rect 11253 23545 11287 23579
rect 14749 23545 14783 23579
rect 15393 23545 15427 23579
rect 17417 23545 17451 23579
rect 17877 23545 17911 23579
rect 18521 23545 18555 23579
rect 19248 23545 19282 23579
rect 13829 23477 13863 23511
rect 14381 23477 14415 23511
rect 15301 23477 15335 23511
rect 16681 23477 16715 23511
rect 18797 23477 18831 23511
rect 20361 23477 20395 23511
rect 21005 23477 21039 23511
rect 21465 23477 21499 23511
rect 21925 23477 21959 23511
rect 23121 23477 23155 23511
rect 23857 23477 23891 23511
rect 24409 23477 24443 23511
rect 13185 23273 13219 23307
rect 13645 23273 13679 23307
rect 15577 23273 15611 23307
rect 17233 23273 17267 23307
rect 18153 23273 18187 23307
rect 19717 23273 19751 23307
rect 21373 23273 21407 23307
rect 23305 23273 23339 23307
rect 23949 23273 23983 23307
rect 24685 23273 24719 23307
rect 16120 23205 16154 23239
rect 18582 23205 18616 23239
rect 11060 23137 11094 23171
rect 13737 23137 13771 23171
rect 18337 23137 18371 23171
rect 21281 23137 21315 23171
rect 24501 23137 24535 23171
rect 10793 23069 10827 23103
rect 13829 23069 13863 23103
rect 14381 23069 14415 23103
rect 15853 23069 15887 23103
rect 21465 23069 21499 23103
rect 23397 23069 23431 23103
rect 23581 23069 23615 23103
rect 12817 23001 12851 23035
rect 20913 23001 20947 23035
rect 12173 22933 12207 22967
rect 13277 22933 13311 22967
rect 14933 22933 14967 22967
rect 22937 22933 22971 22967
rect 24317 22933 24351 22967
rect 10793 22729 10827 22763
rect 11253 22729 11287 22763
rect 13829 22729 13863 22763
rect 14381 22729 14415 22763
rect 15945 22729 15979 22763
rect 16405 22729 16439 22763
rect 17049 22729 17083 22763
rect 17509 22729 17543 22763
rect 17785 22729 17819 22763
rect 18061 22729 18095 22763
rect 21557 22729 21591 22763
rect 22937 22729 22971 22763
rect 25421 22729 25455 22763
rect 12173 22661 12207 22695
rect 22661 22661 22695 22695
rect 12449 22593 12483 22627
rect 15577 22593 15611 22627
rect 18521 22593 18555 22627
rect 18613 22593 18647 22627
rect 22201 22593 22235 22627
rect 24225 22593 24259 22627
rect 16865 22525 16899 22559
rect 18429 22525 18463 22559
rect 19441 22525 19475 22559
rect 20177 22525 20211 22559
rect 24041 22525 24075 22559
rect 12716 22457 12750 22491
rect 14841 22457 14875 22491
rect 20422 22457 20456 22491
rect 24133 22457 24167 22491
rect 14933 22389 14967 22423
rect 15301 22389 15335 22423
rect 15393 22389 15427 22423
rect 19165 22389 19199 22423
rect 20085 22389 20119 22423
rect 23489 22389 23523 22423
rect 23673 22389 23707 22423
rect 24777 22389 24811 22423
rect 11437 22185 11471 22219
rect 12909 22185 12943 22219
rect 13277 22185 13311 22219
rect 17325 22185 17359 22219
rect 18429 22185 18463 22219
rect 18889 22185 18923 22219
rect 20269 22185 20303 22219
rect 20729 22185 20763 22219
rect 21649 22185 21683 22219
rect 22661 22185 22695 22219
rect 23029 22185 23063 22219
rect 12173 22049 12207 22083
rect 12541 22049 12575 22083
rect 15761 22049 15795 22083
rect 21005 22049 21039 22083
rect 22109 22049 22143 22083
rect 23388 22049 23422 22083
rect 11529 21981 11563 22015
rect 11713 21981 11747 22015
rect 13369 21981 13403 22015
rect 13553 21981 13587 22015
rect 15025 21981 15059 22015
rect 15853 21981 15887 22015
rect 15945 21981 15979 22015
rect 17417 21981 17451 22015
rect 17601 21981 17635 22015
rect 18981 21981 19015 22015
rect 19073 21981 19107 22015
rect 22017 21981 22051 22015
rect 23121 21981 23155 22015
rect 15393 21913 15427 21947
rect 21189 21913 21223 21947
rect 11069 21845 11103 21879
rect 13921 21845 13955 21879
rect 16405 21845 16439 21879
rect 16957 21845 16991 21879
rect 18521 21845 18555 21879
rect 19533 21845 19567 21879
rect 22293 21845 22327 21879
rect 24501 21845 24535 21879
rect 11069 21641 11103 21675
rect 13553 21641 13587 21675
rect 15945 21641 15979 21675
rect 16589 21641 16623 21675
rect 18889 21641 18923 21675
rect 20361 21641 20395 21675
rect 22017 21641 22051 21675
rect 21925 21573 21959 21607
rect 13001 21505 13035 21539
rect 14381 21505 14415 21539
rect 15393 21505 15427 21539
rect 16957 21505 16991 21539
rect 18981 21505 19015 21539
rect 21557 21505 21591 21539
rect 22477 21505 22511 21539
rect 22569 21505 22603 21539
rect 14749 21437 14783 21471
rect 15209 21437 15243 21471
rect 16405 21437 16439 21471
rect 19248 21437 19282 21471
rect 22385 21437 22419 21471
rect 24133 21437 24167 21471
rect 24389 21437 24423 21471
rect 10793 21369 10827 21403
rect 12909 21369 12943 21403
rect 15301 21369 15335 21403
rect 17417 21369 17451 21403
rect 11529 21301 11563 21335
rect 11805 21301 11839 21335
rect 12173 21301 12207 21335
rect 12449 21301 12483 21335
rect 12817 21301 12851 21335
rect 13921 21301 13955 21335
rect 14841 21301 14875 21335
rect 16221 21301 16255 21335
rect 17785 21301 17819 21335
rect 18429 21301 18463 21335
rect 21097 21301 21131 21335
rect 23213 21301 23247 21335
rect 23949 21301 23983 21335
rect 25513 21301 25547 21335
rect 13461 21097 13495 21131
rect 14013 21097 14047 21131
rect 15117 21097 15151 21131
rect 17693 21097 17727 21131
rect 18613 21097 18647 21131
rect 21741 21097 21775 21131
rect 23213 21097 23247 21131
rect 23765 21097 23799 21131
rect 15761 21029 15795 21063
rect 16681 21029 16715 21063
rect 17601 21029 17635 21063
rect 1409 20961 1443 20995
rect 11785 20961 11819 20995
rect 15669 20961 15703 20995
rect 19165 20961 19199 20995
rect 19809 20961 19843 20995
rect 21833 20961 21867 20995
rect 22100 20961 22134 20995
rect 24685 20961 24719 20995
rect 11529 20893 11563 20927
rect 15853 20893 15887 20927
rect 17877 20893 17911 20927
rect 19257 20893 19291 20927
rect 19441 20893 19475 20927
rect 24777 20893 24811 20927
rect 24961 20893 24995 20927
rect 1593 20825 1627 20859
rect 13829 20825 13863 20859
rect 12909 20757 12943 20791
rect 14749 20757 14783 20791
rect 15301 20757 15335 20791
rect 17049 20757 17083 20791
rect 17233 20757 17267 20791
rect 18797 20757 18831 20791
rect 20545 20757 20579 20791
rect 24133 20757 24167 20791
rect 24317 20757 24351 20791
rect 11253 20553 11287 20587
rect 11805 20553 11839 20587
rect 12449 20553 12483 20587
rect 16037 20553 16071 20587
rect 16957 20553 16991 20587
rect 19441 20553 19475 20587
rect 20085 20553 20119 20587
rect 21833 20553 21867 20587
rect 22201 20553 22235 20587
rect 23489 20553 23523 20587
rect 25513 20553 25547 20587
rect 25881 20553 25915 20587
rect 16589 20485 16623 20519
rect 10333 20417 10367 20451
rect 13001 20417 13035 20451
rect 13461 20417 13495 20451
rect 17877 20417 17911 20451
rect 18061 20417 18095 20451
rect 21097 20417 21131 20451
rect 24777 20417 24811 20451
rect 1409 20349 1443 20383
rect 14657 20349 14691 20383
rect 20453 20349 20487 20383
rect 21005 20349 21039 20383
rect 22569 20349 22603 20383
rect 24501 20349 24535 20383
rect 12909 20281 12943 20315
rect 13829 20281 13863 20315
rect 14902 20281 14936 20315
rect 17509 20281 17543 20315
rect 18328 20281 18362 20315
rect 24593 20281 24627 20315
rect 1593 20213 1627 20247
rect 1961 20213 1995 20247
rect 11345 20213 11379 20247
rect 12265 20213 12299 20247
rect 12817 20213 12851 20247
rect 14473 20213 14507 20247
rect 20545 20213 20579 20247
rect 20913 20213 20947 20247
rect 23949 20213 23983 20247
rect 24133 20213 24167 20247
rect 25145 20213 25179 20247
rect 13921 20009 13955 20043
rect 17693 20009 17727 20043
rect 18429 20009 18463 20043
rect 18613 20009 18647 20043
rect 22293 20009 22327 20043
rect 23857 20009 23891 20043
rect 12808 19941 12842 19975
rect 15660 19941 15694 19975
rect 19073 19941 19107 19975
rect 21158 19941 21192 19975
rect 24216 19941 24250 19975
rect 10057 19873 10091 19907
rect 10313 19873 10347 19907
rect 12541 19873 12575 19907
rect 14749 19873 14783 19907
rect 15393 19873 15427 19907
rect 18981 19873 19015 19907
rect 20913 19873 20947 19907
rect 17417 19805 17451 19839
rect 19257 19805 19291 19839
rect 23949 19805 23983 19839
rect 19809 19737 19843 19771
rect 1593 19669 1627 19703
rect 11437 19669 11471 19703
rect 16773 19669 16807 19703
rect 18153 19669 18187 19703
rect 20177 19669 20211 19703
rect 20637 19669 20671 19703
rect 22845 19669 22879 19703
rect 25329 19669 25363 19703
rect 9781 19465 9815 19499
rect 11805 19465 11839 19499
rect 16497 19465 16531 19499
rect 19165 19465 19199 19499
rect 20913 19465 20947 19499
rect 22293 19465 22327 19499
rect 25053 19465 25087 19499
rect 18061 19397 18095 19431
rect 19717 19397 19751 19431
rect 10885 19329 10919 19363
rect 11253 19329 11287 19363
rect 13001 19329 13035 19363
rect 14105 19329 14139 19363
rect 14197 19329 14231 19363
rect 17509 19329 17543 19363
rect 18705 19329 18739 19363
rect 20269 19329 20303 19363
rect 21925 19329 21959 19363
rect 24593 19329 24627 19363
rect 9413 19261 9447 19295
rect 10057 19261 10091 19295
rect 10609 19261 10643 19295
rect 12817 19261 12851 19295
rect 16957 19261 16991 19295
rect 18429 19261 18463 19295
rect 21649 19261 21683 19295
rect 23121 19261 23155 19295
rect 24317 19261 24351 19295
rect 25513 19261 25547 19295
rect 26065 19261 26099 19295
rect 12265 19193 12299 19227
rect 13737 19193 13771 19227
rect 14442 19193 14476 19227
rect 20085 19193 20119 19227
rect 23489 19193 23523 19227
rect 24409 19193 24443 19227
rect 25329 19193 25363 19227
rect 10241 19125 10275 19159
rect 10701 19125 10735 19159
rect 12449 19125 12483 19159
rect 12909 19125 12943 19159
rect 15577 19125 15611 19159
rect 16221 19125 16255 19159
rect 17877 19125 17911 19159
rect 18521 19125 18555 19159
rect 19533 19125 19567 19159
rect 20177 19125 20211 19159
rect 21281 19125 21315 19159
rect 21741 19125 21775 19159
rect 22661 19125 22695 19159
rect 23949 19125 23983 19159
rect 25697 19125 25731 19159
rect 12909 18921 12943 18955
rect 13277 18921 13311 18955
rect 13645 18921 13679 18955
rect 14013 18921 14047 18955
rect 14105 18921 14139 18955
rect 15117 18921 15151 18955
rect 15761 18921 15795 18955
rect 19349 18921 19383 18955
rect 21189 18921 21223 18955
rect 21557 18921 21591 18955
rect 22569 18921 22603 18955
rect 23673 18921 23707 18955
rect 15853 18853 15887 18887
rect 19073 18853 19107 18887
rect 24124 18853 24158 18887
rect 10865 18785 10899 18819
rect 17316 18785 17350 18819
rect 19809 18785 19843 18819
rect 22293 18785 22327 18819
rect 10609 18717 10643 18751
rect 14197 18717 14231 18751
rect 16037 18717 16071 18751
rect 17049 18717 17083 18751
rect 21649 18717 21683 18751
rect 21741 18717 21775 18751
rect 22845 18717 22879 18751
rect 23857 18717 23891 18751
rect 18429 18649 18463 18683
rect 20729 18649 20763 18683
rect 10333 18581 10367 18615
rect 11989 18581 12023 18615
rect 12633 18581 12667 18615
rect 14657 18581 14691 18615
rect 15393 18581 15427 18615
rect 16865 18581 16899 18615
rect 19993 18581 20027 18615
rect 25237 18581 25271 18615
rect 10333 18377 10367 18411
rect 10609 18377 10643 18411
rect 14197 18377 14231 18411
rect 15761 18377 15795 18411
rect 16405 18377 16439 18411
rect 17693 18377 17727 18411
rect 18613 18377 18647 18411
rect 20453 18377 20487 18411
rect 21557 18377 21591 18411
rect 23397 18377 23431 18411
rect 24685 18377 24719 18411
rect 25145 18377 25179 18411
rect 10793 18309 10827 18343
rect 11805 18309 11839 18343
rect 13829 18309 13863 18343
rect 16681 18309 16715 18343
rect 11253 18241 11287 18275
rect 11437 18241 11471 18275
rect 13277 18241 13311 18275
rect 22017 18241 22051 18275
rect 22201 18241 22235 18275
rect 24133 18241 24167 18275
rect 24317 18241 24351 18275
rect 9965 18173 9999 18207
rect 13369 18173 13403 18207
rect 14381 18173 14415 18207
rect 14648 18173 14682 18207
rect 16865 18173 16899 18207
rect 18061 18173 18095 18207
rect 19073 18173 19107 18207
rect 22937 18173 22971 18207
rect 24041 18173 24075 18207
rect 25237 18173 25271 18207
rect 25789 18173 25823 18207
rect 17325 18105 17359 18139
rect 18889 18105 18923 18139
rect 19340 18105 19374 18139
rect 21925 18105 21959 18139
rect 22569 18105 22603 18139
rect 11161 18037 11195 18071
rect 13553 18037 13587 18071
rect 17049 18037 17083 18071
rect 18245 18037 18279 18071
rect 21281 18037 21315 18071
rect 23673 18037 23707 18071
rect 25421 18037 25455 18071
rect 13369 17833 13403 17867
rect 13645 17833 13679 17867
rect 15761 17833 15795 17867
rect 16681 17833 16715 17867
rect 19993 17833 20027 17867
rect 20361 17833 20395 17867
rect 20913 17833 20947 17867
rect 21373 17833 21407 17867
rect 23121 17833 23155 17867
rect 23673 17833 23707 17867
rect 24225 17833 24259 17867
rect 11428 17765 11462 17799
rect 14013 17765 14047 17799
rect 14105 17765 14139 17799
rect 14749 17765 14783 17799
rect 17224 17765 17258 17799
rect 11161 17697 11195 17731
rect 15669 17697 15703 17731
rect 19809 17697 19843 17731
rect 21281 17697 21315 17731
rect 23581 17697 23615 17731
rect 24777 17697 24811 17731
rect 14289 17629 14323 17663
rect 15025 17629 15059 17663
rect 15853 17629 15887 17663
rect 16313 17629 16347 17663
rect 16957 17629 16991 17663
rect 21465 17629 21499 17663
rect 23765 17629 23799 17663
rect 23213 17561 23247 17595
rect 10885 17493 10919 17527
rect 12541 17493 12575 17527
rect 15301 17493 15335 17527
rect 18337 17493 18371 17527
rect 19165 17493 19199 17527
rect 20729 17493 20763 17527
rect 22017 17493 22051 17527
rect 24961 17493 24995 17527
rect 11805 17289 11839 17323
rect 12173 17289 12207 17323
rect 14749 17289 14783 17323
rect 16313 17289 16347 17323
rect 22569 17289 22603 17323
rect 25053 17289 25087 17323
rect 25605 17289 25639 17323
rect 22017 17221 22051 17255
rect 22293 17221 22327 17255
rect 10333 17153 10367 17187
rect 11437 17153 11471 17187
rect 12449 17153 12483 17187
rect 14933 17153 14967 17187
rect 21833 17153 21867 17187
rect 10701 17085 10735 17119
rect 12705 17085 12739 17119
rect 17417 17085 17451 17119
rect 18705 17085 18739 17119
rect 11161 17017 11195 17051
rect 15178 17017 15212 17051
rect 18972 17017 19006 17051
rect 21005 17017 21039 17051
rect 21557 17017 21591 17051
rect 23489 17085 23523 17119
rect 23673 17085 23707 17119
rect 23940 17085 23974 17119
rect 10793 16949 10827 16983
rect 11253 16949 11287 16983
rect 13829 16949 13863 16983
rect 14381 16949 14415 16983
rect 16957 16949 16991 16983
rect 18521 16949 18555 16983
rect 20085 16949 20119 16983
rect 21189 16949 21223 16983
rect 21649 16949 21683 16983
rect 22017 16949 22051 16983
rect 23029 16949 23063 16983
rect 11253 16745 11287 16779
rect 12541 16745 12575 16779
rect 13737 16745 13771 16779
rect 14105 16745 14139 16779
rect 15117 16745 15151 16779
rect 16405 16745 16439 16779
rect 18889 16745 18923 16779
rect 19809 16745 19843 16779
rect 20361 16745 20395 16779
rect 20729 16745 20763 16779
rect 22293 16745 22327 16779
rect 22937 16745 22971 16779
rect 23489 16745 23523 16779
rect 24593 16745 24627 16779
rect 25237 16745 25271 16779
rect 11713 16677 11747 16711
rect 14657 16677 14691 16711
rect 15761 16677 15795 16711
rect 21158 16677 21192 16711
rect 23213 16677 23247 16711
rect 10885 16609 10919 16643
rect 15669 16609 15703 16643
rect 16865 16609 16899 16643
rect 17132 16609 17166 16643
rect 20913 16609 20947 16643
rect 23857 16609 23891 16643
rect 25053 16609 25087 16643
rect 11805 16541 11839 16575
rect 11989 16541 12023 16575
rect 14197 16541 14231 16575
rect 15853 16541 15887 16575
rect 23949 16541 23983 16575
rect 24133 16541 24167 16575
rect 15301 16473 15335 16507
rect 11345 16405 11379 16439
rect 18245 16405 18279 16439
rect 11161 16201 11195 16235
rect 11897 16201 11931 16235
rect 14197 16201 14231 16235
rect 14657 16201 14691 16235
rect 15761 16201 15795 16235
rect 18521 16201 18555 16235
rect 21189 16201 21223 16235
rect 23489 16201 23523 16235
rect 24225 16201 24259 16235
rect 25513 16201 25547 16235
rect 12173 16133 12207 16167
rect 21741 16133 21775 16167
rect 11345 16065 11379 16099
rect 15209 16065 15243 16099
rect 17049 16065 17083 16099
rect 17877 16065 17911 16099
rect 19073 16065 19107 16099
rect 19165 16065 19199 16099
rect 19717 16065 19751 16099
rect 20729 16065 20763 16099
rect 21557 16065 21591 16099
rect 22293 16065 22327 16099
rect 12449 15997 12483 16031
rect 12909 15997 12943 16031
rect 15025 15997 15059 16031
rect 16773 15997 16807 16031
rect 18981 15997 19015 16031
rect 20637 15997 20671 16031
rect 22109 15997 22143 16031
rect 24593 15997 24627 16031
rect 25145 15997 25179 16031
rect 16313 15929 16347 15963
rect 16865 15929 16899 15963
rect 22201 15929 22235 15963
rect 22753 15929 22787 15963
rect 12633 15861 12667 15895
rect 14473 15861 14507 15895
rect 15117 15861 15151 15895
rect 16405 15861 16439 15895
rect 17417 15861 17451 15895
rect 18613 15861 18647 15895
rect 20085 15861 20119 15895
rect 20177 15861 20211 15895
rect 20545 15861 20579 15895
rect 23857 15861 23891 15895
rect 24777 15861 24811 15895
rect 14657 15657 14691 15691
rect 15117 15657 15151 15691
rect 16681 15657 16715 15691
rect 17049 15657 17083 15691
rect 19165 15657 19199 15691
rect 20269 15657 20303 15691
rect 21373 15657 21407 15691
rect 21833 15657 21867 15691
rect 23305 15657 23339 15691
rect 14197 15521 14231 15555
rect 15945 15521 15979 15555
rect 17408 15521 17442 15555
rect 20913 15521 20947 15555
rect 21925 15521 21959 15555
rect 22192 15521 22226 15555
rect 24593 15521 24627 15555
rect 16037 15453 16071 15487
rect 16221 15453 16255 15487
rect 17141 15453 17175 15487
rect 19625 15453 19659 15487
rect 14381 15385 14415 15419
rect 24777 15385 24811 15419
rect 15577 15317 15611 15351
rect 18521 15317 18555 15351
rect 21097 15317 21131 15351
rect 14289 15113 14323 15147
rect 14749 15113 14783 15147
rect 15761 15113 15795 15147
rect 16221 15113 16255 15147
rect 20821 15113 20855 15147
rect 21925 15113 21959 15147
rect 22293 15113 22327 15147
rect 22753 15113 22787 15147
rect 24501 15113 24535 15147
rect 16681 14977 16715 15011
rect 16773 14977 16807 15011
rect 13001 14909 13035 14943
rect 13461 14909 13495 14943
rect 16129 14909 16163 14943
rect 17601 14909 17635 14943
rect 18521 14909 18555 14943
rect 18777 14909 18811 14943
rect 21005 14909 21039 14943
rect 22569 14909 22603 14943
rect 24593 14909 24627 14943
rect 25145 14909 25179 14943
rect 15117 14841 15151 14875
rect 21465 14841 21499 14875
rect 13185 14773 13219 14807
rect 15209 14773 15243 14807
rect 16589 14773 16623 14807
rect 17233 14773 17267 14807
rect 18337 14773 18371 14807
rect 19901 14773 19935 14807
rect 21189 14773 21223 14807
rect 23121 14773 23155 14807
rect 24777 14773 24811 14807
rect 15761 14569 15795 14603
rect 17417 14569 17451 14603
rect 18153 14569 18187 14603
rect 18613 14569 18647 14603
rect 19073 14569 19107 14603
rect 19441 14569 19475 14603
rect 25421 14569 25455 14603
rect 15117 14501 15151 14535
rect 16282 14501 16316 14535
rect 13093 14433 13127 14467
rect 14105 14433 14139 14467
rect 16037 14433 16071 14467
rect 20913 14433 20947 14467
rect 23020 14433 23054 14467
rect 25237 14433 25271 14467
rect 18981 14365 19015 14399
rect 19533 14365 19567 14399
rect 19625 14365 19659 14399
rect 22753 14365 22787 14399
rect 14289 14297 14323 14331
rect 20085 14297 20119 14331
rect 13277 14229 13311 14263
rect 21097 14229 21131 14263
rect 24133 14229 24167 14263
rect 13093 14025 13127 14059
rect 14657 14025 14691 14059
rect 15761 14025 15795 14059
rect 17141 14025 17175 14059
rect 18061 14025 18095 14059
rect 19165 14025 19199 14059
rect 21557 14025 21591 14059
rect 23029 14025 23063 14059
rect 23673 14025 23707 14059
rect 25789 14025 25823 14059
rect 14381 13957 14415 13991
rect 15301 13957 15335 13991
rect 23397 13957 23431 13991
rect 25421 13957 25455 13991
rect 16221 13889 16255 13923
rect 16405 13889 16439 13923
rect 18613 13889 18647 13923
rect 24225 13889 24259 13923
rect 25053 13889 25087 13923
rect 14013 13821 14047 13855
rect 14197 13821 14231 13855
rect 15577 13821 15611 13855
rect 16129 13821 16163 13855
rect 16865 13821 16899 13855
rect 18521 13821 18555 13855
rect 19533 13821 19567 13855
rect 19625 13821 19659 13855
rect 19881 13821 19915 13855
rect 25237 13821 25271 13855
rect 17785 13753 17819 13787
rect 18429 13753 18463 13787
rect 22477 13753 22511 13787
rect 21005 13685 21039 13719
rect 22569 13685 22603 13719
rect 24041 13685 24075 13719
rect 24133 13685 24167 13719
rect 14105 13481 14139 13515
rect 15485 13481 15519 13515
rect 16865 13481 16899 13515
rect 17417 13481 17451 13515
rect 18061 13481 18095 13515
rect 19165 13481 19199 13515
rect 19625 13481 19659 13515
rect 22201 13481 22235 13515
rect 23029 13481 23063 13515
rect 23121 13481 23155 13515
rect 23765 13481 23799 13515
rect 24777 13481 24811 13515
rect 16589 13413 16623 13447
rect 17509 13413 17543 13447
rect 14013 13345 14047 13379
rect 15853 13345 15887 13379
rect 21281 13345 21315 13379
rect 24593 13345 24627 13379
rect 14289 13277 14323 13311
rect 15945 13277 15979 13311
rect 16037 13277 16071 13311
rect 17693 13277 17727 13311
rect 19717 13277 19751 13311
rect 19809 13277 19843 13311
rect 21373 13277 21407 13311
rect 21465 13277 21499 13311
rect 23305 13277 23339 13311
rect 15117 13209 15151 13243
rect 17049 13209 17083 13243
rect 18797 13209 18831 13243
rect 19257 13209 19291 13243
rect 22661 13209 22695 13243
rect 24041 13209 24075 13243
rect 13645 13141 13679 13175
rect 14657 13141 14691 13175
rect 20729 13141 20763 13175
rect 20913 13141 20947 13175
rect 13093 12937 13127 12971
rect 16129 12937 16163 12971
rect 16865 12937 16899 12971
rect 18613 12937 18647 12971
rect 20177 12937 20211 12971
rect 20545 12937 20579 12971
rect 23029 12937 23063 12971
rect 24501 12937 24535 12971
rect 13737 12869 13771 12903
rect 18245 12869 18279 12903
rect 22385 12869 22419 12903
rect 17877 12801 17911 12835
rect 18889 12801 18923 12835
rect 19625 12801 19659 12835
rect 21281 12801 21315 12835
rect 22753 12801 22787 12835
rect 14197 12733 14231 12767
rect 14464 12733 14498 12767
rect 16681 12733 16715 12767
rect 17233 12733 17267 12767
rect 18061 12733 18095 12767
rect 19533 12733 19567 12767
rect 21649 12733 21683 12767
rect 22201 12733 22235 12767
rect 24593 12733 24627 12767
rect 25145 12733 25179 12767
rect 14105 12665 14139 12699
rect 19441 12665 19475 12699
rect 13185 12597 13219 12631
rect 15577 12597 15611 12631
rect 16589 12597 16623 12631
rect 19073 12597 19107 12631
rect 20637 12597 20671 12631
rect 21005 12597 21039 12631
rect 21097 12597 21131 12631
rect 22109 12597 22143 12631
rect 23489 12597 23523 12631
rect 24777 12597 24811 12631
rect 12449 12393 12483 12427
rect 13645 12393 13679 12427
rect 15025 12393 15059 12427
rect 17049 12393 17083 12427
rect 19165 12393 19199 12427
rect 20729 12393 20763 12427
rect 23765 12393 23799 12427
rect 12541 12325 12575 12359
rect 18153 12325 18187 12359
rect 20361 12325 20395 12359
rect 21364 12325 21398 12359
rect 13185 12257 13219 12291
rect 14013 12257 14047 12291
rect 15925 12257 15959 12291
rect 19625 12257 19659 12291
rect 23581 12257 23615 12291
rect 24409 12257 24443 12291
rect 24593 12257 24627 12291
rect 12725 12189 12759 12223
rect 13553 12189 13587 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 15676 12189 15710 12223
rect 19717 12189 19751 12223
rect 19901 12189 19935 12223
rect 21097 12189 21131 12223
rect 12081 12121 12115 12155
rect 18061 12121 18095 12155
rect 19257 12121 19291 12155
rect 14657 12053 14691 12087
rect 15485 12053 15519 12087
rect 17601 12053 17635 12087
rect 18613 12053 18647 12087
rect 22477 12053 22511 12087
rect 24133 12053 24167 12087
rect 24777 12053 24811 12087
rect 11437 11849 11471 11883
rect 12173 11849 12207 11883
rect 13185 11849 13219 11883
rect 15025 11849 15059 11883
rect 15669 11849 15703 11883
rect 17141 11849 17175 11883
rect 19441 11849 19475 11883
rect 21925 11849 21959 11883
rect 23489 11849 23523 11883
rect 24685 11849 24719 11883
rect 11805 11713 11839 11747
rect 13553 11713 13587 11747
rect 13645 11713 13679 11747
rect 16681 11713 16715 11747
rect 24133 11713 24167 11747
rect 24225 11713 24259 11747
rect 16497 11645 16531 11679
rect 18061 11645 18095 11679
rect 20545 11645 20579 11679
rect 12817 11577 12851 11611
rect 13890 11577 13924 11611
rect 18306 11577 18340 11611
rect 20812 11577 20846 11611
rect 24041 11577 24075 11611
rect 16129 11509 16163 11543
rect 16589 11509 16623 11543
rect 17785 11509 17819 11543
rect 20085 11509 20119 11543
rect 20453 11509 20487 11543
rect 22477 11509 22511 11543
rect 23029 11509 23063 11543
rect 23673 11509 23707 11543
rect 12081 11305 12115 11339
rect 13645 11305 13679 11339
rect 14657 11305 14691 11339
rect 15117 11305 15151 11339
rect 15761 11305 15795 11339
rect 18337 11305 18371 11339
rect 18981 11305 19015 11339
rect 19809 11305 19843 11339
rect 21465 11305 21499 11339
rect 25237 11305 25271 11339
rect 17202 11237 17236 11271
rect 12449 11169 12483 11203
rect 13553 11169 13587 11203
rect 14013 11169 14047 11203
rect 15669 11169 15703 11203
rect 21281 11169 21315 11203
rect 22560 11169 22594 11203
rect 25145 11169 25179 11203
rect 11621 11101 11655 11135
rect 12541 11101 12575 11135
rect 12633 11101 12667 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 15853 11101 15887 11135
rect 16957 11101 16991 11135
rect 21741 11101 21775 11135
rect 22293 11101 22327 11135
rect 25421 11101 25455 11135
rect 15301 11033 15335 11067
rect 16313 11033 16347 11067
rect 16681 11033 16715 11067
rect 19441 11033 19475 11067
rect 21189 11033 21223 11067
rect 24777 11033 24811 11067
rect 1593 10965 1627 10999
rect 11897 10965 11931 10999
rect 13093 10965 13127 10999
rect 20545 10965 20579 10999
rect 23673 10965 23707 10999
rect 24225 10965 24259 10999
rect 11529 10761 11563 10795
rect 11897 10761 11931 10795
rect 14105 10761 14139 10795
rect 15209 10761 15243 10795
rect 15393 10761 15427 10795
rect 16957 10761 16991 10795
rect 17325 10761 17359 10795
rect 18245 10761 18279 10795
rect 22845 10761 22879 10795
rect 25973 10761 26007 10795
rect 10885 10693 10919 10727
rect 11253 10693 11287 10727
rect 12449 10693 12483 10727
rect 14933 10693 14967 10727
rect 12909 10625 12943 10659
rect 13001 10625 13035 10659
rect 14657 10625 14691 10659
rect 1409 10557 1443 10591
rect 1676 10557 1710 10591
rect 11345 10557 11379 10591
rect 12265 10557 12299 10591
rect 13645 10557 13679 10591
rect 12817 10489 12851 10523
rect 14013 10489 14047 10523
rect 14473 10489 14507 10523
rect 14933 10489 14967 10523
rect 18797 10693 18831 10727
rect 16221 10625 16255 10659
rect 18981 10625 19015 10659
rect 22017 10625 22051 10659
rect 15577 10557 15611 10591
rect 16037 10557 16071 10591
rect 19237 10557 19271 10591
rect 21373 10557 21407 10591
rect 21925 10557 21959 10591
rect 23673 10557 23707 10591
rect 15393 10489 15427 10523
rect 16129 10489 16163 10523
rect 20913 10489 20947 10523
rect 21833 10489 21867 10523
rect 23918 10489 23952 10523
rect 2789 10421 2823 10455
rect 14565 10421 14599 10455
rect 15669 10421 15703 10455
rect 20361 10421 20395 10455
rect 21465 10421 21499 10455
rect 22569 10421 22603 10455
rect 23397 10421 23431 10455
rect 25053 10421 25087 10455
rect 25605 10421 25639 10455
rect 1685 10217 1719 10251
rect 11069 10217 11103 10251
rect 12633 10217 12667 10251
rect 13737 10217 13771 10251
rect 14381 10217 14415 10251
rect 15301 10217 15335 10251
rect 16313 10217 16347 10251
rect 16681 10217 16715 10251
rect 16865 10217 16899 10251
rect 18429 10217 18463 10251
rect 18797 10217 18831 10251
rect 19533 10217 19567 10251
rect 20913 10217 20947 10251
rect 21925 10217 21959 10251
rect 22477 10217 22511 10251
rect 23029 10217 23063 10251
rect 25421 10217 25455 10251
rect 12173 10149 12207 10183
rect 13001 10149 13035 10183
rect 14105 10149 14139 10183
rect 15761 10149 15795 10183
rect 23734 10149 23768 10183
rect 11437 10081 11471 10115
rect 13093 10081 13127 10115
rect 14197 10081 14231 10115
rect 15669 10081 15703 10115
rect 17233 10081 17267 10115
rect 18889 10081 18923 10115
rect 21281 10081 21315 10115
rect 10977 10013 11011 10047
rect 11529 10013 11563 10047
rect 11713 10013 11747 10047
rect 13185 10013 13219 10047
rect 15945 10013 15979 10047
rect 17325 10013 17359 10047
rect 17417 10013 17451 10047
rect 18981 10013 19015 10047
rect 21373 10013 21407 10047
rect 21465 10013 21499 10047
rect 23489 10013 23523 10047
rect 12541 9877 12575 9911
rect 14749 9877 14783 9911
rect 15025 9877 15059 9911
rect 18153 9877 18187 9911
rect 24869 9877 24903 9911
rect 16037 9673 16071 9707
rect 19901 9673 19935 9707
rect 20729 9673 20763 9707
rect 22109 9673 22143 9707
rect 11253 9605 11287 9639
rect 12449 9605 12483 9639
rect 14565 9605 14599 9639
rect 17417 9605 17451 9639
rect 17877 9605 17911 9639
rect 18061 9605 18095 9639
rect 21741 9605 21775 9639
rect 13001 9537 13035 9571
rect 13461 9537 13495 9571
rect 16681 9537 16715 9571
rect 18521 9537 18555 9571
rect 18705 9537 18739 9571
rect 19441 9537 19475 9571
rect 21281 9537 21315 9571
rect 22477 9537 22511 9571
rect 9873 9469 9907 9503
rect 10140 9469 10174 9503
rect 12817 9469 12851 9503
rect 14657 9469 14691 9503
rect 20637 9469 20671 9503
rect 21097 9469 21131 9503
rect 21189 9469 21223 9503
rect 24133 9469 24167 9503
rect 24400 9469 24434 9503
rect 14924 9401 14958 9435
rect 18429 9401 18463 9435
rect 20269 9401 20303 9435
rect 9689 9333 9723 9367
rect 11805 9333 11839 9367
rect 12265 9333 12299 9367
rect 12909 9333 12943 9367
rect 13921 9333 13955 9367
rect 16957 9333 16991 9367
rect 19073 9333 19107 9367
rect 23029 9333 23063 9367
rect 23397 9333 23431 9367
rect 23949 9333 23983 9367
rect 25513 9333 25547 9367
rect 9965 9129 9999 9163
rect 12633 9129 12667 9163
rect 13185 9129 13219 9163
rect 14289 9129 14323 9163
rect 16681 9129 16715 9163
rect 17785 9129 17819 9163
rect 18245 9129 18279 9163
rect 19993 9129 20027 9163
rect 21097 9129 21131 9163
rect 23121 9129 23155 9163
rect 23673 9129 23707 9163
rect 24225 9129 24259 9163
rect 11161 9061 11195 9095
rect 11520 9061 11554 9095
rect 15117 9061 15151 9095
rect 21465 9061 21499 9095
rect 23029 9061 23063 9095
rect 24133 9061 24167 9095
rect 11253 8993 11287 9027
rect 15568 8993 15602 9027
rect 17601 8993 17635 9027
rect 18153 8993 18187 9027
rect 24593 8993 24627 9027
rect 24685 8993 24719 9027
rect 25237 8993 25271 9027
rect 15301 8925 15335 8959
rect 18337 8925 18371 8959
rect 19533 8925 19567 8959
rect 20729 8925 20763 8959
rect 21557 8925 21591 8959
rect 21741 8925 21775 8959
rect 23305 8925 23339 8959
rect 24777 8925 24811 8959
rect 17233 8857 17267 8891
rect 22661 8857 22695 8891
rect 14749 8789 14783 8823
rect 18797 8789 18831 8823
rect 22201 8789 22235 8823
rect 22477 8789 22511 8823
rect 11161 8585 11195 8619
rect 11805 8585 11839 8619
rect 12173 8585 12207 8619
rect 17049 8585 17083 8619
rect 17509 8585 17543 8619
rect 18061 8585 18095 8619
rect 21281 8585 21315 8619
rect 22201 8585 22235 8619
rect 22937 8585 22971 8619
rect 21833 8517 21867 8551
rect 22569 8517 22603 8551
rect 11345 8449 11379 8483
rect 12449 8449 12483 8483
rect 18705 8449 18739 8483
rect 14749 8381 14783 8415
rect 14933 8381 14967 8415
rect 17785 8381 17819 8415
rect 18521 8381 18555 8415
rect 19901 8381 19935 8415
rect 20157 8381 20191 8415
rect 22385 8381 22419 8415
rect 24133 8381 24167 8415
rect 12694 8313 12728 8347
rect 14473 8313 14507 8347
rect 15200 8313 15234 8347
rect 18429 8313 18463 8347
rect 19073 8313 19107 8347
rect 24041 8313 24075 8347
rect 24400 8313 24434 8347
rect 13829 8245 13863 8279
rect 16313 8245 16347 8279
rect 19809 8245 19843 8279
rect 23397 8245 23431 8279
rect 25513 8245 25547 8279
rect 12909 8041 12943 8075
rect 13921 8041 13955 8075
rect 14933 8041 14967 8075
rect 15301 8041 15335 8075
rect 16589 8041 16623 8075
rect 16957 8041 16991 8075
rect 17877 8041 17911 8075
rect 18153 8041 18187 8075
rect 19441 8041 19475 8075
rect 21097 8041 21131 8075
rect 24961 8041 24995 8075
rect 15853 7973 15887 8007
rect 21557 7973 21591 8007
rect 24593 7973 24627 8007
rect 12265 7905 12299 7939
rect 13829 7905 13863 7939
rect 17049 7905 17083 7939
rect 18521 7905 18555 7939
rect 21465 7905 21499 7939
rect 22928 7905 22962 7939
rect 12357 7837 12391 7871
rect 12449 7837 12483 7871
rect 14105 7837 14139 7871
rect 17233 7837 17267 7871
rect 18613 7837 18647 7871
rect 18705 7837 18739 7871
rect 19809 7837 19843 7871
rect 20729 7837 20763 7871
rect 21741 7837 21775 7871
rect 22661 7837 22695 7871
rect 11897 7701 11931 7735
rect 13461 7701 13495 7735
rect 16497 7701 16531 7735
rect 22385 7701 22419 7735
rect 24041 7701 24075 7735
rect 11989 7497 12023 7531
rect 12725 7497 12759 7531
rect 17785 7497 17819 7531
rect 18337 7497 18371 7531
rect 18889 7497 18923 7531
rect 21465 7497 21499 7531
rect 21833 7497 21867 7531
rect 13093 7429 13127 7463
rect 16405 7429 16439 7463
rect 23673 7429 23707 7463
rect 11621 7361 11655 7395
rect 14473 7361 14507 7395
rect 14933 7361 14967 7395
rect 16865 7361 16899 7395
rect 16957 7361 16991 7395
rect 19349 7361 19383 7395
rect 22477 7361 22511 7395
rect 22661 7361 22695 7395
rect 23489 7361 23523 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 25053 7361 25087 7395
rect 13461 7293 13495 7327
rect 14381 7293 14415 7327
rect 16313 7293 16347 7327
rect 18429 7293 18463 7327
rect 19441 7293 19475 7327
rect 22385 7293 22419 7327
rect 23029 7293 23063 7327
rect 14289 7225 14323 7259
rect 15945 7225 15979 7259
rect 16773 7225 16807 7259
rect 19686 7225 19720 7259
rect 24041 7225 24075 7259
rect 24777 7225 24811 7259
rect 25237 7225 25271 7259
rect 13737 7157 13771 7191
rect 13921 7157 13955 7191
rect 17509 7157 17543 7191
rect 18613 7157 18647 7191
rect 20821 7157 20855 7191
rect 22017 7157 22051 7191
rect 11989 6953 12023 6987
rect 13645 6953 13679 6987
rect 16957 6953 16991 6987
rect 17325 6953 17359 6987
rect 22661 6953 22695 6987
rect 24133 6953 24167 6987
rect 15761 6885 15795 6919
rect 16865 6885 16899 6919
rect 21557 6885 21591 6919
rect 13093 6817 13127 6851
rect 13553 6817 13587 6851
rect 15117 6817 15151 6851
rect 17417 6817 17451 6851
rect 18889 6817 18923 6851
rect 19809 6817 19843 6851
rect 22753 6817 22787 6851
rect 23020 6817 23054 6851
rect 25237 6817 25271 6851
rect 13737 6749 13771 6783
rect 15853 6749 15887 6783
rect 15945 6749 15979 6783
rect 17601 6749 17635 6783
rect 18981 6749 19015 6783
rect 19073 6749 19107 6783
rect 21649 6749 21683 6783
rect 21741 6749 21775 6783
rect 12725 6681 12759 6715
rect 18521 6681 18555 6715
rect 21189 6681 21223 6715
rect 13185 6613 13219 6647
rect 14197 6613 14231 6647
rect 15393 6613 15427 6647
rect 16497 6613 16531 6647
rect 18429 6613 18463 6647
rect 20729 6613 20763 6647
rect 22201 6613 22235 6647
rect 25421 6613 25455 6647
rect 15209 6409 15243 6443
rect 15301 6409 15335 6443
rect 17417 6409 17451 6443
rect 17785 6409 17819 6443
rect 18613 6409 18647 6443
rect 21833 6409 21867 6443
rect 22017 6409 22051 6443
rect 23029 6409 23063 6443
rect 24041 6409 24075 6443
rect 25237 6409 25271 6443
rect 13645 6273 13679 6307
rect 14105 6273 14139 6307
rect 14657 6273 14691 6307
rect 22477 6273 22511 6307
rect 22661 6273 22695 6307
rect 24685 6273 24719 6307
rect 24869 6273 24903 6307
rect 13553 6205 13587 6239
rect 15209 6205 15243 6239
rect 15485 6205 15519 6239
rect 15752 6205 15786 6239
rect 19533 6205 19567 6239
rect 19800 6205 19834 6239
rect 12265 6137 12299 6171
rect 13461 6137 13495 6171
rect 14933 6137 14967 6171
rect 19349 6137 19383 6171
rect 22385 6137 22419 6171
rect 23489 6137 23523 6171
rect 24593 6137 24627 6171
rect 12909 6069 12943 6103
rect 13093 6069 13127 6103
rect 16865 6069 16899 6103
rect 18061 6069 18095 6103
rect 18889 6069 18923 6103
rect 20913 6069 20947 6103
rect 21557 6069 21591 6103
rect 24225 6069 24259 6103
rect 14013 5865 14047 5899
rect 15117 5865 15151 5899
rect 19533 5865 19567 5899
rect 20729 5865 20763 5899
rect 22385 5865 22419 5899
rect 25237 5865 25271 5899
rect 12326 5797 12360 5831
rect 15669 5797 15703 5831
rect 16589 5797 16623 5831
rect 16957 5797 16991 5831
rect 17316 5797 17350 5831
rect 19073 5797 19107 5831
rect 21373 5797 21407 5831
rect 15761 5729 15795 5763
rect 19717 5729 19751 5763
rect 21281 5729 21315 5763
rect 22477 5729 22511 5763
rect 24041 5729 24075 5763
rect 12081 5661 12115 5695
rect 15945 5661 15979 5695
rect 17049 5661 17083 5695
rect 21465 5661 21499 5695
rect 24133 5661 24167 5695
rect 24317 5661 24351 5695
rect 13461 5593 13495 5627
rect 15301 5593 15335 5627
rect 22661 5593 22695 5627
rect 23581 5593 23615 5627
rect 11989 5525 12023 5559
rect 18429 5525 18463 5559
rect 19901 5525 19935 5559
rect 20361 5525 20395 5559
rect 20913 5525 20947 5559
rect 22017 5525 22051 5559
rect 23121 5525 23155 5559
rect 23673 5525 23707 5559
rect 24777 5525 24811 5559
rect 25053 5525 25087 5559
rect 12081 5321 12115 5355
rect 15485 5321 15519 5355
rect 16129 5321 16163 5355
rect 19901 5321 19935 5355
rect 21005 5321 21039 5355
rect 21373 5321 21407 5355
rect 22017 5321 22051 5355
rect 23029 5321 23063 5355
rect 25789 5321 25823 5355
rect 11253 5253 11287 5287
rect 18337 5253 18371 5287
rect 19993 5253 20027 5287
rect 25237 5253 25271 5287
rect 11345 5185 11379 5219
rect 13185 5185 13219 5219
rect 13553 5185 13587 5219
rect 17417 5185 17451 5219
rect 19073 5185 19107 5219
rect 20637 5185 20671 5219
rect 21925 5185 21959 5219
rect 22661 5185 22695 5219
rect 22845 5185 22879 5219
rect 12909 5117 12943 5151
rect 14013 5117 14047 5151
rect 14105 5117 14139 5151
rect 16865 5117 16899 5151
rect 18889 5117 18923 5151
rect 20361 5117 20395 5151
rect 22477 5117 22511 5151
rect 23857 5117 23891 5151
rect 13001 5049 13035 5083
rect 14350 5049 14384 5083
rect 17785 5049 17819 5083
rect 20453 5049 20487 5083
rect 22385 5049 22419 5083
rect 22845 5049 22879 5083
rect 24102 5049 24136 5083
rect 12541 4981 12575 5015
rect 16681 4981 16715 5015
rect 17049 4981 17083 5015
rect 18429 4981 18463 5015
rect 18797 4981 18831 5015
rect 19533 4981 19567 5015
rect 23397 4981 23431 5015
rect 12081 4777 12115 4811
rect 13553 4777 13587 4811
rect 14197 4777 14231 4811
rect 15117 4777 15151 4811
rect 16865 4777 16899 4811
rect 17325 4777 17359 4811
rect 18153 4777 18187 4811
rect 18889 4777 18923 4811
rect 19993 4777 20027 4811
rect 20729 4777 20763 4811
rect 22937 4777 22971 4811
rect 17417 4709 17451 4743
rect 12173 4641 12207 4675
rect 12440 4641 12474 4675
rect 15853 4641 15887 4675
rect 18981 4641 19015 4675
rect 21169 4641 21203 4675
rect 23653 4641 23687 4675
rect 17509 4573 17543 4607
rect 19073 4573 19107 4607
rect 20913 4573 20947 4607
rect 23397 4573 23431 4607
rect 16497 4505 16531 4539
rect 18521 4505 18555 4539
rect 22293 4505 22327 4539
rect 14749 4437 14783 4471
rect 15577 4437 15611 4471
rect 16037 4437 16071 4471
rect 16957 4437 16991 4471
rect 19717 4437 19751 4471
rect 23213 4437 23247 4471
rect 24777 4437 24811 4471
rect 12173 4233 12207 4267
rect 12633 4233 12667 4267
rect 15853 4233 15887 4267
rect 17233 4233 17267 4267
rect 21005 4233 21039 4267
rect 21925 4233 21959 4267
rect 25053 4233 25087 4267
rect 17693 4165 17727 4199
rect 17785 4165 17819 4199
rect 18061 4165 18095 4199
rect 21557 4165 21591 4199
rect 23397 4165 23431 4199
rect 15577 4097 15611 4131
rect 16681 4097 16715 4131
rect 18521 4097 18555 4131
rect 18613 4097 18647 4131
rect 23673 4097 23707 4131
rect 11345 4029 11379 4063
rect 13185 4029 13219 4063
rect 13369 4029 13403 4063
rect 16589 4029 16623 4063
rect 17693 4029 17727 4063
rect 18429 4029 18463 4063
rect 19165 4029 19199 4063
rect 19625 4029 19659 4063
rect 22201 4029 22235 4063
rect 22753 4029 22787 4063
rect 11897 3961 11931 3995
rect 13614 3961 13648 3995
rect 16497 3961 16531 3995
rect 19892 3961 19926 3995
rect 23918 3961 23952 3995
rect 11529 3893 11563 3927
rect 14749 3893 14783 3927
rect 16129 3893 16163 3927
rect 19441 3893 19475 3927
rect 22385 3893 22419 3927
rect 12725 3689 12759 3723
rect 13461 3689 13495 3723
rect 14105 3689 14139 3723
rect 18613 3689 18647 3723
rect 19257 3689 19291 3723
rect 19901 3689 19935 3723
rect 20729 3689 20763 3723
rect 21281 3689 21315 3723
rect 22109 3689 22143 3723
rect 22477 3689 22511 3723
rect 23305 3689 23339 3723
rect 24869 3689 24903 3723
rect 25237 3689 25271 3723
rect 14657 3621 14691 3655
rect 22569 3621 22603 3655
rect 22753 3621 22787 3655
rect 23213 3621 23247 3655
rect 10425 3553 10459 3587
rect 11437 3553 11471 3587
rect 12541 3553 12575 3587
rect 14013 3553 14047 3587
rect 15301 3553 15335 3587
rect 16129 3553 16163 3587
rect 16405 3553 16439 3587
rect 16672 3553 16706 3587
rect 14289 3485 14323 3519
rect 19349 3485 19383 3519
rect 19441 3485 19475 3519
rect 21373 3485 21407 3519
rect 21557 3485 21591 3519
rect 23673 3553 23707 3587
rect 23765 3485 23799 3519
rect 23949 3485 23983 3519
rect 25329 3485 25363 3519
rect 25513 3485 25547 3519
rect 13645 3417 13679 3451
rect 20913 3417 20947 3451
rect 22569 3417 22603 3451
rect 24409 3417 24443 3451
rect 10609 3349 10643 3383
rect 11621 3349 11655 3383
rect 15025 3349 15059 3383
rect 15485 3349 15519 3383
rect 17785 3349 17819 3383
rect 18889 3349 18923 3383
rect 20361 3349 20395 3383
rect 10149 3145 10183 3179
rect 10701 3145 10735 3179
rect 11161 3145 11195 3179
rect 13001 3145 13035 3179
rect 13369 3145 13403 3179
rect 14105 3145 14139 3179
rect 16497 3145 16531 3179
rect 17049 3145 17083 3179
rect 20729 3145 20763 3179
rect 21741 3145 21775 3179
rect 23305 3145 23339 3179
rect 23857 3145 23891 3179
rect 25145 3145 25179 3179
rect 25881 3145 25915 3179
rect 10425 3077 10459 3111
rect 11437 3077 11471 3111
rect 15945 3077 15979 3111
rect 19625 3077 19659 3111
rect 22109 3077 22143 3111
rect 24409 3077 24443 3111
rect 9781 3009 9815 3043
rect 12449 3009 12483 3043
rect 14381 3009 14415 3043
rect 14565 3009 14599 3043
rect 17785 3009 17819 3043
rect 18245 3009 18279 3043
rect 20269 3009 20303 3043
rect 21281 3009 21315 3043
rect 25513 3009 25547 3043
rect 9229 2941 9263 2975
rect 10241 2941 10275 2975
rect 11253 2941 11287 2975
rect 13461 2941 13495 2975
rect 20545 2941 20579 2975
rect 21097 2941 21131 2975
rect 22477 2941 22511 2975
rect 24593 2941 24627 2975
rect 11805 2873 11839 2907
rect 14832 2873 14866 2907
rect 18490 2873 18524 2907
rect 21189 2873 21223 2907
rect 9413 2805 9447 2839
rect 13645 2805 13679 2839
rect 17417 2805 17451 2839
rect 22661 2805 22695 2839
rect 24777 2805 24811 2839
rect 2973 2601 3007 2635
rect 5733 2601 5767 2635
rect 8309 2601 8343 2635
rect 10885 2601 10919 2635
rect 13093 2601 13127 2635
rect 16037 2601 16071 2635
rect 16497 2601 16531 2635
rect 17141 2601 17175 2635
rect 19073 2601 19107 2635
rect 19533 2601 19567 2635
rect 19901 2601 19935 2635
rect 20821 2601 20855 2635
rect 22661 2601 22695 2635
rect 23857 2601 23891 2635
rect 13737 2533 13771 2567
rect 14197 2533 14231 2567
rect 15761 2533 15795 2567
rect 16405 2533 16439 2567
rect 18061 2533 18095 2567
rect 2789 2465 2823 2499
rect 3341 2465 3375 2499
rect 5549 2465 5583 2499
rect 6101 2465 6135 2499
rect 8125 2465 8159 2499
rect 10333 2465 10367 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 13185 2465 13219 2499
rect 14289 2465 14323 2499
rect 14933 2465 14967 2499
rect 17785 2465 17819 2499
rect 18429 2465 18463 2499
rect 19441 2465 19475 2499
rect 21741 2465 21775 2499
rect 22293 2465 22327 2499
rect 22845 2465 22879 2499
rect 23397 2465 23431 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 12449 2397 12483 2431
rect 16589 2397 16623 2431
rect 19993 2397 20027 2431
rect 20085 2397 20119 2431
rect 14473 2329 14507 2363
rect 15301 2329 15335 2363
rect 18613 2329 18647 2363
rect 21373 2329 21407 2363
rect 23029 2329 23063 2363
rect 24777 2329 24811 2363
rect 8677 2261 8711 2295
rect 10517 2261 10551 2295
rect 11621 2261 11655 2295
rect 13369 2261 13403 2295
rect 21925 2261 21959 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 14461 25483 14519 25489
rect 14461 25449 14473 25483
rect 14507 25480 14519 25483
rect 15286 25480 15292 25492
rect 14507 25452 15292 25480
rect 14507 25449 14519 25452
rect 14461 25443 14519 25449
rect 15286 25440 15292 25452
rect 15344 25440 15350 25492
rect 15657 25483 15715 25489
rect 15657 25449 15669 25483
rect 15703 25480 15715 25483
rect 16574 25480 16580 25492
rect 15703 25452 16580 25480
rect 15703 25449 15715 25452
rect 15657 25443 15715 25449
rect 16574 25440 16580 25452
rect 16632 25440 16638 25492
rect 16853 25483 16911 25489
rect 16853 25449 16865 25483
rect 16899 25480 16911 25483
rect 17954 25480 17960 25492
rect 16899 25452 17960 25480
rect 16899 25449 16911 25452
rect 16853 25443 16911 25449
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 19613 25483 19671 25489
rect 19613 25449 19625 25483
rect 19659 25480 19671 25483
rect 20070 25480 20076 25492
rect 19659 25452 20076 25480
rect 19659 25449 19671 25452
rect 19613 25443 19671 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 22189 25483 22247 25489
rect 22189 25449 22201 25483
rect 22235 25480 22247 25483
rect 22738 25480 22744 25492
rect 22235 25452 22744 25480
rect 22235 25449 22247 25452
rect 22189 25443 22247 25449
rect 22738 25440 22744 25452
rect 22796 25440 22802 25492
rect 14277 25347 14335 25353
rect 14277 25313 14289 25347
rect 14323 25344 14335 25347
rect 14366 25344 14372 25356
rect 14323 25316 14372 25344
rect 14323 25313 14335 25316
rect 14277 25307 14335 25313
rect 14366 25304 14372 25316
rect 14424 25304 14430 25356
rect 15473 25347 15531 25353
rect 15473 25313 15485 25347
rect 15519 25344 15531 25347
rect 15562 25344 15568 25356
rect 15519 25316 15568 25344
rect 15519 25313 15531 25316
rect 15473 25307 15531 25313
rect 15562 25304 15568 25316
rect 15620 25304 15626 25356
rect 16666 25344 16672 25356
rect 16627 25316 16672 25344
rect 16666 25304 16672 25316
rect 16724 25304 16730 25356
rect 19334 25304 19340 25356
rect 19392 25344 19398 25356
rect 19429 25347 19487 25353
rect 19429 25344 19441 25347
rect 19392 25316 19441 25344
rect 19392 25304 19398 25316
rect 19429 25313 19441 25316
rect 19475 25313 19487 25347
rect 22002 25344 22008 25356
rect 21963 25316 22008 25344
rect 19429 25307 19487 25313
rect 22002 25304 22008 25316
rect 22060 25304 22066 25356
rect 18141 25279 18199 25285
rect 18141 25245 18153 25279
rect 18187 25276 18199 25279
rect 18325 25279 18383 25285
rect 18325 25276 18337 25279
rect 18187 25248 18337 25276
rect 18187 25245 18199 25248
rect 18141 25239 18199 25245
rect 18325 25245 18337 25248
rect 18371 25276 18383 25279
rect 18414 25276 18420 25288
rect 18371 25248 18420 25276
rect 18371 25245 18383 25248
rect 18325 25239 18383 25245
rect 18414 25236 18420 25248
rect 18472 25236 18478 25288
rect 16117 25143 16175 25149
rect 16117 25109 16129 25143
rect 16163 25140 16175 25143
rect 16390 25140 16396 25152
rect 16163 25112 16396 25140
rect 16163 25109 16175 25112
rect 16117 25103 16175 25109
rect 16390 25100 16396 25112
rect 16448 25100 16454 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 18874 24896 18880 24948
rect 18932 24936 18938 24948
rect 24762 24936 24768 24948
rect 18932 24908 24768 24936
rect 18932 24896 18938 24908
rect 24762 24896 24768 24908
rect 24820 24896 24826 24948
rect 17512 24840 19380 24868
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 9582 24800 9588 24812
rect 8444 24772 9588 24800
rect 8444 24760 8450 24772
rect 9582 24760 9588 24772
rect 9640 24760 9646 24812
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 15933 24803 15991 24809
rect 15933 24800 15945 24803
rect 15436 24772 15945 24800
rect 15436 24760 15442 24772
rect 15933 24769 15945 24772
rect 15979 24769 15991 24803
rect 15933 24763 15991 24769
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24800 16175 24803
rect 16390 24800 16396 24812
rect 16163 24772 16396 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 16390 24760 16396 24772
rect 16448 24800 16454 24812
rect 17512 24809 17540 24840
rect 18708 24809 18736 24840
rect 17497 24803 17555 24809
rect 17497 24800 17509 24803
rect 16448 24772 17509 24800
rect 16448 24760 16454 24772
rect 17497 24769 17509 24772
rect 17543 24769 17555 24803
rect 17497 24763 17555 24769
rect 18693 24803 18751 24809
rect 18693 24769 18705 24803
rect 18739 24769 18751 24803
rect 19352 24800 19380 24840
rect 21450 24828 21456 24880
rect 21508 24868 21514 24880
rect 22002 24868 22008 24880
rect 21508 24840 22008 24868
rect 21508 24828 21514 24840
rect 22002 24828 22008 24840
rect 22060 24828 22066 24880
rect 23658 24868 23664 24880
rect 22112 24840 23664 24868
rect 19352 24772 20760 24800
rect 18693 24763 18751 24769
rect 12805 24735 12863 24741
rect 12805 24701 12817 24735
rect 12851 24732 12863 24735
rect 13909 24735 13967 24741
rect 12851 24704 13308 24732
rect 12851 24701 12863 24704
rect 12805 24695 12863 24701
rect 13280 24608 13308 24704
rect 13909 24701 13921 24735
rect 13955 24732 13967 24735
rect 14369 24735 14427 24741
rect 14369 24732 14381 24735
rect 13955 24704 14381 24732
rect 13955 24701 13967 24704
rect 13909 24695 13967 24701
rect 14369 24701 14381 24704
rect 14415 24732 14427 24735
rect 14642 24732 14648 24744
rect 14415 24704 14648 24732
rect 14415 24701 14427 24704
rect 14369 24695 14427 24701
rect 14642 24692 14648 24704
rect 14700 24692 14706 24744
rect 15010 24732 15016 24744
rect 14923 24704 15016 24732
rect 15010 24692 15016 24704
rect 15068 24732 15074 24744
rect 15841 24735 15899 24741
rect 15841 24732 15853 24735
rect 15068 24704 15853 24732
rect 15068 24692 15074 24704
rect 15841 24701 15853 24704
rect 15887 24701 15899 24735
rect 18414 24732 18420 24744
rect 18375 24704 18420 24732
rect 15841 24695 15899 24701
rect 18414 24692 18420 24704
rect 18472 24692 18478 24744
rect 19978 24732 19984 24744
rect 19939 24704 19984 24732
rect 19978 24692 19984 24704
rect 20036 24732 20042 24744
rect 20533 24735 20591 24741
rect 20533 24732 20545 24735
rect 20036 24704 20545 24732
rect 20036 24692 20042 24704
rect 20533 24701 20545 24704
rect 20579 24701 20591 24735
rect 20533 24695 20591 24701
rect 15381 24667 15439 24673
rect 15381 24633 15393 24667
rect 15427 24664 15439 24667
rect 15562 24664 15568 24676
rect 15427 24636 15568 24664
rect 15427 24633 15439 24636
rect 15381 24627 15439 24633
rect 15562 24624 15568 24636
rect 15620 24624 15626 24676
rect 17494 24624 17500 24676
rect 17552 24664 17558 24676
rect 17865 24667 17923 24673
rect 17865 24664 17877 24667
rect 17552 24636 17877 24664
rect 17552 24624 17558 24636
rect 17865 24633 17877 24636
rect 17911 24664 17923 24667
rect 18509 24667 18567 24673
rect 18509 24664 18521 24667
rect 17911 24636 18521 24664
rect 17911 24633 17923 24636
rect 17865 24627 17923 24633
rect 18509 24633 18521 24636
rect 18555 24633 18567 24667
rect 20732 24664 20760 24772
rect 21174 24760 21180 24812
rect 21232 24800 21238 24812
rect 22112 24800 22140 24840
rect 23658 24828 23664 24840
rect 23716 24828 23722 24880
rect 21232 24772 22140 24800
rect 21232 24760 21238 24772
rect 21082 24732 21088 24744
rect 21043 24704 21088 24732
rect 21082 24692 21088 24704
rect 21140 24732 21146 24744
rect 21637 24735 21695 24741
rect 21637 24732 21649 24735
rect 21140 24704 21649 24732
rect 21140 24692 21146 24704
rect 21637 24701 21649 24704
rect 21683 24701 21695 24735
rect 21637 24695 21695 24701
rect 21726 24692 21732 24744
rect 21784 24732 21790 24744
rect 22189 24735 22247 24741
rect 22189 24732 22201 24735
rect 21784 24704 22201 24732
rect 21784 24692 21790 24704
rect 22189 24701 22201 24704
rect 22235 24732 22247 24735
rect 22741 24735 22799 24741
rect 22741 24732 22753 24735
rect 22235 24704 22753 24732
rect 22235 24701 22247 24704
rect 22189 24695 22247 24701
rect 22741 24701 22753 24704
rect 22787 24701 22799 24735
rect 22741 24695 22799 24701
rect 21818 24664 21824 24676
rect 20732 24636 21824 24664
rect 18509 24627 18567 24633
rect 21818 24624 21824 24636
rect 21876 24624 21882 24676
rect 12986 24596 12992 24608
rect 12947 24568 12992 24596
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 13262 24556 13268 24608
rect 13320 24596 13326 24608
rect 13357 24599 13415 24605
rect 13357 24596 13369 24599
rect 13320 24568 13369 24596
rect 13320 24556 13326 24568
rect 13357 24565 13369 24568
rect 13403 24565 13415 24599
rect 13357 24559 13415 24565
rect 14277 24599 14335 24605
rect 14277 24565 14289 24599
rect 14323 24596 14335 24599
rect 14366 24596 14372 24608
rect 14323 24568 14372 24596
rect 14323 24565 14335 24568
rect 14277 24559 14335 24565
rect 14366 24556 14372 24568
rect 14424 24556 14430 24608
rect 14550 24596 14556 24608
rect 14511 24568 14556 24596
rect 14550 24556 14556 24568
rect 14608 24556 14614 24608
rect 15470 24596 15476 24608
rect 15431 24568 15476 24596
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 16666 24556 16672 24608
rect 16724 24596 16730 24608
rect 16761 24599 16819 24605
rect 16761 24596 16773 24599
rect 16724 24568 16773 24596
rect 16724 24556 16730 24568
rect 16761 24565 16773 24568
rect 16807 24596 16819 24599
rect 17126 24596 17132 24608
rect 16807 24568 17132 24596
rect 16807 24565 16819 24568
rect 16761 24559 16819 24565
rect 17126 24556 17132 24568
rect 17184 24556 17190 24608
rect 18049 24599 18107 24605
rect 18049 24565 18061 24599
rect 18095 24596 18107 24599
rect 18322 24596 18328 24608
rect 18095 24568 18328 24596
rect 18095 24565 18107 24568
rect 18049 24559 18107 24565
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 19334 24556 19340 24608
rect 19392 24596 19398 24608
rect 19429 24599 19487 24605
rect 19429 24596 19441 24599
rect 19392 24568 19441 24596
rect 19392 24556 19398 24568
rect 19429 24565 19441 24568
rect 19475 24565 19487 24599
rect 20162 24596 20168 24608
rect 20123 24568 20168 24596
rect 19429 24559 19487 24565
rect 20162 24556 20168 24568
rect 20220 24556 20226 24608
rect 21266 24596 21272 24608
rect 21227 24568 21272 24596
rect 21266 24556 21272 24568
rect 21324 24556 21330 24608
rect 22373 24599 22431 24605
rect 22373 24565 22385 24599
rect 22419 24596 22431 24599
rect 24118 24596 24124 24608
rect 22419 24568 24124 24596
rect 22419 24565 22431 24568
rect 22373 24559 22431 24565
rect 24118 24556 24124 24568
rect 24176 24556 24182 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 12342 24392 12348 24404
rect 12303 24364 12348 24392
rect 12342 24352 12348 24364
rect 12400 24352 12406 24404
rect 15470 24352 15476 24404
rect 15528 24392 15534 24404
rect 16298 24392 16304 24404
rect 15528 24364 16304 24392
rect 15528 24352 15534 24364
rect 16298 24352 16304 24364
rect 16356 24352 16362 24404
rect 19797 24395 19855 24401
rect 19797 24361 19809 24395
rect 19843 24392 19855 24395
rect 20622 24392 20628 24404
rect 19843 24364 20628 24392
rect 19843 24361 19855 24364
rect 19797 24355 19855 24361
rect 20622 24352 20628 24364
rect 20680 24352 20686 24404
rect 23658 24392 23664 24404
rect 23619 24364 23664 24392
rect 23658 24352 23664 24364
rect 23716 24352 23722 24404
rect 24762 24392 24768 24404
rect 24723 24364 24768 24392
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 11514 24216 11520 24268
rect 11572 24256 11578 24268
rect 12253 24259 12311 24265
rect 12253 24256 12265 24259
rect 11572 24228 12265 24256
rect 11572 24216 11578 24228
rect 12253 24225 12265 24228
rect 12299 24225 12311 24259
rect 12253 24219 12311 24225
rect 13357 24259 13415 24265
rect 13357 24225 13369 24259
rect 13403 24256 13415 24259
rect 13814 24256 13820 24268
rect 13403 24228 13820 24256
rect 13403 24225 13415 24228
rect 13357 24219 13415 24225
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 13909 24259 13967 24265
rect 13909 24225 13921 24259
rect 13955 24256 13967 24259
rect 14458 24256 14464 24268
rect 13955 24228 14464 24256
rect 13955 24225 13967 24228
rect 13909 24219 13967 24225
rect 14458 24216 14464 24228
rect 14516 24216 14522 24268
rect 15378 24216 15384 24268
rect 15436 24256 15442 24268
rect 15473 24259 15531 24265
rect 15473 24256 15485 24259
rect 15436 24228 15485 24256
rect 15436 24216 15442 24228
rect 15473 24225 15485 24228
rect 15519 24225 15531 24259
rect 15473 24219 15531 24225
rect 16022 24216 16028 24268
rect 16080 24256 16086 24268
rect 16209 24259 16267 24265
rect 16209 24256 16221 24259
rect 16080 24228 16221 24256
rect 16080 24216 16086 24228
rect 16209 24225 16221 24228
rect 16255 24225 16267 24259
rect 16209 24219 16267 24225
rect 17313 24259 17371 24265
rect 17313 24225 17325 24259
rect 17359 24256 17371 24259
rect 18046 24256 18052 24268
rect 17359 24228 18052 24256
rect 17359 24225 17371 24228
rect 17313 24219 17371 24225
rect 18046 24216 18052 24228
rect 18104 24256 18110 24268
rect 18141 24259 18199 24265
rect 18141 24256 18153 24259
rect 18104 24228 18153 24256
rect 18104 24216 18110 24228
rect 18141 24225 18153 24228
rect 18187 24225 18199 24259
rect 18141 24219 18199 24225
rect 18598 24216 18604 24268
rect 18656 24256 18662 24268
rect 19613 24259 19671 24265
rect 19613 24256 19625 24259
rect 18656 24228 19625 24256
rect 18656 24216 18662 24228
rect 19613 24225 19625 24228
rect 19659 24225 19671 24259
rect 21266 24256 21272 24268
rect 21227 24228 21272 24256
rect 19613 24219 19671 24225
rect 21266 24216 21272 24228
rect 21324 24216 21330 24268
rect 23477 24259 23535 24265
rect 23477 24225 23489 24259
rect 23523 24256 23535 24259
rect 23842 24256 23848 24268
rect 23523 24228 23848 24256
rect 23523 24225 23535 24228
rect 23477 24219 23535 24225
rect 23842 24216 23848 24228
rect 23900 24216 23906 24268
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24176 24228 24593 24256
rect 24176 24216 24182 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 12710 24188 12716 24200
rect 12575 24160 12716 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 12710 24148 12716 24160
rect 12768 24188 12774 24200
rect 13998 24188 14004 24200
rect 12768 24160 13032 24188
rect 13959 24160 14004 24188
rect 12768 24148 12774 24160
rect 13004 24129 13032 24160
rect 13998 24148 14004 24160
rect 14056 24148 14062 24200
rect 16114 24148 16120 24200
rect 16172 24188 16178 24200
rect 16393 24191 16451 24197
rect 16393 24188 16405 24191
rect 16172 24160 16405 24188
rect 16172 24148 16178 24160
rect 16393 24157 16405 24160
rect 16439 24188 16451 24191
rect 16482 24188 16488 24200
rect 16439 24160 16488 24188
rect 16439 24157 16451 24160
rect 16393 24151 16451 24157
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24157 18291 24191
rect 18414 24188 18420 24200
rect 18375 24160 18420 24188
rect 18233 24151 18291 24157
rect 12989 24123 13047 24129
rect 12989 24089 13001 24123
rect 13035 24120 13047 24123
rect 13035 24092 14504 24120
rect 13035 24089 13047 24092
rect 12989 24083 13047 24089
rect 11885 24055 11943 24061
rect 11885 24021 11897 24055
rect 11931 24052 11943 24055
rect 12342 24052 12348 24064
rect 11931 24024 12348 24052
rect 11931 24021 11943 24024
rect 11885 24015 11943 24021
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 13446 24052 13452 24064
rect 13407 24024 13452 24052
rect 13446 24012 13452 24024
rect 13504 24012 13510 24064
rect 14476 24052 14504 24092
rect 14550 24080 14556 24132
rect 14608 24120 14614 24132
rect 15010 24120 15016 24132
rect 14608 24092 15016 24120
rect 14608 24080 14614 24092
rect 15010 24080 15016 24092
rect 15068 24080 15074 24132
rect 15841 24123 15899 24129
rect 15841 24089 15853 24123
rect 15887 24120 15899 24123
rect 17589 24123 17647 24129
rect 17589 24120 17601 24123
rect 15887 24092 17601 24120
rect 15887 24089 15899 24092
rect 15841 24083 15899 24089
rect 17589 24089 17601 24092
rect 17635 24120 17647 24123
rect 18248 24120 18276 24151
rect 18414 24148 18420 24160
rect 18472 24148 18478 24200
rect 21174 24148 21180 24200
rect 21232 24188 21238 24200
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 21232 24160 21373 24188
rect 21232 24148 21238 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 21545 24191 21603 24197
rect 21545 24157 21557 24191
rect 21591 24188 21603 24191
rect 21818 24188 21824 24200
rect 21591 24160 21824 24188
rect 21591 24157 21603 24160
rect 21545 24151 21603 24157
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 22465 24191 22523 24197
rect 22465 24157 22477 24191
rect 22511 24188 22523 24191
rect 23566 24188 23572 24200
rect 22511 24160 23572 24188
rect 22511 24157 22523 24160
rect 22465 24151 22523 24157
rect 23566 24148 23572 24160
rect 23624 24148 23630 24200
rect 17635 24092 18276 24120
rect 17635 24089 17647 24092
rect 17589 24083 17647 24089
rect 14921 24055 14979 24061
rect 14921 24052 14933 24055
rect 14476 24024 14933 24052
rect 14921 24021 14933 24024
rect 14967 24052 14979 24055
rect 15654 24052 15660 24064
rect 14967 24024 15660 24052
rect 14967 24021 14979 24024
rect 14921 24015 14979 24021
rect 15654 24012 15660 24024
rect 15712 24012 15718 24064
rect 17770 24052 17776 24064
rect 17731 24024 17776 24052
rect 17770 24012 17776 24024
rect 17828 24012 17834 24064
rect 18966 24052 18972 24064
rect 18927 24024 18972 24052
rect 18966 24012 18972 24024
rect 19024 24012 19030 24064
rect 20898 24052 20904 24064
rect 20859 24024 20904 24052
rect 20898 24012 20904 24024
rect 20956 24012 20962 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 11514 23848 11520 23860
rect 11475 23820 11520 23848
rect 11514 23808 11520 23820
rect 11572 23808 11578 23860
rect 11977 23851 12035 23857
rect 11977 23817 11989 23851
rect 12023 23848 12035 23851
rect 12250 23848 12256 23860
rect 12023 23820 12256 23848
rect 12023 23817 12035 23820
rect 11977 23811 12035 23817
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 13814 23808 13820 23860
rect 13872 23848 13878 23860
rect 14921 23851 14979 23857
rect 14921 23848 14933 23851
rect 13872 23820 14933 23848
rect 13872 23808 13878 23820
rect 14921 23817 14933 23820
rect 14967 23817 14979 23851
rect 14921 23811 14979 23817
rect 16025 23851 16083 23857
rect 16025 23817 16037 23851
rect 16071 23848 16083 23851
rect 16114 23848 16120 23860
rect 16071 23820 16120 23848
rect 16071 23817 16083 23820
rect 16025 23811 16083 23817
rect 16114 23808 16120 23820
rect 16172 23808 16178 23860
rect 16298 23848 16304 23860
rect 16259 23820 16304 23848
rect 16298 23808 16304 23820
rect 16356 23808 16362 23860
rect 17034 23848 17040 23860
rect 16995 23820 17040 23848
rect 17034 23808 17040 23820
rect 17092 23808 17098 23860
rect 20990 23808 20996 23860
rect 21048 23848 21054 23860
rect 21266 23848 21272 23860
rect 21048 23820 21272 23848
rect 21048 23808 21054 23820
rect 21266 23808 21272 23820
rect 21324 23808 21330 23860
rect 22646 23848 22652 23860
rect 22607 23820 22652 23848
rect 22646 23808 22652 23820
rect 22704 23808 22710 23860
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23712 15623 23715
rect 15654 23712 15660 23724
rect 15611 23684 15660 23712
rect 15611 23681 15623 23684
rect 15565 23675 15623 23681
rect 15654 23672 15660 23684
rect 15712 23672 15718 23724
rect 24118 23672 24124 23724
rect 24176 23712 24182 23724
rect 25133 23715 25191 23721
rect 25133 23712 25145 23715
rect 24176 23684 25145 23712
rect 24176 23672 24182 23684
rect 25133 23681 25145 23684
rect 25179 23681 25191 23715
rect 25133 23675 25191 23681
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 12710 23653 12716 23656
rect 12704 23644 12716 23653
rect 12492 23616 12537 23644
rect 12636 23616 12716 23644
rect 12492 23604 12498 23616
rect 11241 23579 11299 23585
rect 11241 23545 11253 23579
rect 11287 23576 11299 23579
rect 12636 23576 12664 23616
rect 12704 23607 12716 23616
rect 12710 23604 12716 23607
rect 12768 23604 12774 23656
rect 16853 23647 16911 23653
rect 16853 23613 16865 23647
rect 16899 23613 16911 23647
rect 18966 23644 18972 23656
rect 18927 23616 18972 23644
rect 16853 23607 16911 23613
rect 11287 23548 12664 23576
rect 11287 23545 11299 23548
rect 11241 23539 11299 23545
rect 14274 23536 14280 23588
rect 14332 23576 14338 23588
rect 14737 23579 14795 23585
rect 14737 23576 14749 23579
rect 14332 23548 14749 23576
rect 14332 23536 14338 23548
rect 14737 23545 14749 23548
rect 14783 23576 14795 23579
rect 15381 23579 15439 23585
rect 15381 23576 15393 23579
rect 14783 23548 15393 23576
rect 14783 23545 14795 23548
rect 14737 23539 14795 23545
rect 15381 23545 15393 23548
rect 15427 23576 15439 23579
rect 16868 23576 16896 23607
rect 18966 23604 18972 23616
rect 19024 23604 19030 23656
rect 22465 23647 22523 23653
rect 22465 23613 22477 23647
rect 22511 23644 22523 23647
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 22511 23616 23152 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 17405 23579 17463 23585
rect 17405 23576 17417 23579
rect 15427 23548 17417 23576
rect 15427 23545 15439 23548
rect 15381 23539 15439 23545
rect 17405 23545 17417 23548
rect 17451 23545 17463 23579
rect 17405 23539 17463 23545
rect 17865 23579 17923 23585
rect 17865 23545 17877 23579
rect 17911 23576 17923 23579
rect 18414 23576 18420 23588
rect 17911 23548 18420 23576
rect 17911 23545 17923 23548
rect 17865 23539 17923 23545
rect 18414 23536 18420 23548
rect 18472 23576 18478 23588
rect 18509 23579 18567 23585
rect 18509 23576 18521 23579
rect 18472 23548 18521 23576
rect 18472 23536 18478 23548
rect 18509 23545 18521 23548
rect 18555 23576 18567 23579
rect 19236 23579 19294 23585
rect 19236 23576 19248 23579
rect 18555 23548 19248 23576
rect 18555 23545 18567 23548
rect 18509 23539 18567 23545
rect 19236 23545 19248 23548
rect 19282 23576 19294 23579
rect 19426 23576 19432 23588
rect 19282 23548 19432 23576
rect 19282 23545 19294 23548
rect 19236 23539 19294 23545
rect 19426 23536 19432 23548
rect 19484 23536 19490 23588
rect 23124 23520 23152 23616
rect 24412 23616 24593 23644
rect 13814 23508 13820 23520
rect 13775 23480 13820 23508
rect 13814 23468 13820 23480
rect 13872 23508 13878 23520
rect 13998 23508 14004 23520
rect 13872 23480 14004 23508
rect 13872 23468 13878 23480
rect 13998 23468 14004 23480
rect 14056 23508 14062 23520
rect 14369 23511 14427 23517
rect 14369 23508 14381 23511
rect 14056 23480 14381 23508
rect 14056 23468 14062 23480
rect 14369 23477 14381 23480
rect 14415 23477 14427 23511
rect 15286 23508 15292 23520
rect 15247 23480 15292 23508
rect 14369 23471 14427 23477
rect 15286 23468 15292 23480
rect 15344 23468 15350 23520
rect 16022 23468 16028 23520
rect 16080 23508 16086 23520
rect 16669 23511 16727 23517
rect 16669 23508 16681 23511
rect 16080 23480 16681 23508
rect 16080 23468 16086 23480
rect 16669 23477 16681 23480
rect 16715 23477 16727 23511
rect 16669 23471 16727 23477
rect 18598 23468 18604 23520
rect 18656 23508 18662 23520
rect 18785 23511 18843 23517
rect 18785 23508 18797 23511
rect 18656 23480 18797 23508
rect 18656 23468 18662 23480
rect 18785 23477 18797 23480
rect 18831 23477 18843 23511
rect 18785 23471 18843 23477
rect 20349 23511 20407 23517
rect 20349 23477 20361 23511
rect 20395 23508 20407 23511
rect 20622 23508 20628 23520
rect 20395 23480 20628 23508
rect 20395 23477 20407 23480
rect 20349 23471 20407 23477
rect 20622 23468 20628 23480
rect 20680 23468 20686 23520
rect 20993 23511 21051 23517
rect 20993 23477 21005 23511
rect 21039 23508 21051 23511
rect 21174 23508 21180 23520
rect 21039 23480 21180 23508
rect 21039 23477 21051 23480
rect 20993 23471 21051 23477
rect 21174 23468 21180 23480
rect 21232 23468 21238 23520
rect 21453 23511 21511 23517
rect 21453 23477 21465 23511
rect 21499 23508 21511 23511
rect 21542 23508 21548 23520
rect 21499 23480 21548 23508
rect 21499 23477 21511 23480
rect 21453 23471 21511 23477
rect 21542 23468 21548 23480
rect 21600 23468 21606 23520
rect 21818 23468 21824 23520
rect 21876 23508 21882 23520
rect 21913 23511 21971 23517
rect 21913 23508 21925 23511
rect 21876 23480 21925 23508
rect 21876 23468 21882 23480
rect 21913 23477 21925 23480
rect 21959 23477 21971 23511
rect 23106 23508 23112 23520
rect 23067 23480 23112 23508
rect 21913 23471 21971 23477
rect 23106 23468 23112 23480
rect 23164 23468 23170 23520
rect 23842 23508 23848 23520
rect 23803 23480 23848 23508
rect 23842 23468 23848 23480
rect 23900 23468 23906 23520
rect 24026 23468 24032 23520
rect 24084 23508 24090 23520
rect 24412 23517 24440 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24084 23480 24409 23508
rect 24084 23468 24090 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 13173 23307 13231 23313
rect 13173 23273 13185 23307
rect 13219 23304 13231 23307
rect 13446 23304 13452 23316
rect 13219 23276 13452 23304
rect 13219 23273 13231 23276
rect 13173 23267 13231 23273
rect 13446 23264 13452 23276
rect 13504 23304 13510 23316
rect 13633 23307 13691 23313
rect 13633 23304 13645 23307
rect 13504 23276 13645 23304
rect 13504 23264 13510 23276
rect 13633 23273 13645 23276
rect 13679 23273 13691 23307
rect 13633 23267 13691 23273
rect 15565 23307 15623 23313
rect 15565 23273 15577 23307
rect 15611 23304 15623 23307
rect 15654 23304 15660 23316
rect 15611 23276 15660 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 17221 23307 17279 23313
rect 17221 23304 17233 23307
rect 16632 23276 17233 23304
rect 16632 23264 16638 23276
rect 17221 23273 17233 23276
rect 17267 23304 17279 23307
rect 17770 23304 17776 23316
rect 17267 23276 17776 23304
rect 17267 23273 17279 23276
rect 17221 23267 17279 23273
rect 17770 23264 17776 23276
rect 17828 23264 17834 23316
rect 18138 23304 18144 23316
rect 18099 23276 18144 23304
rect 18138 23264 18144 23276
rect 18196 23264 18202 23316
rect 19426 23264 19432 23316
rect 19484 23304 19490 23316
rect 19705 23307 19763 23313
rect 19705 23304 19717 23307
rect 19484 23276 19717 23304
rect 19484 23264 19490 23276
rect 19705 23273 19717 23276
rect 19751 23273 19763 23307
rect 19705 23267 19763 23273
rect 21361 23307 21419 23313
rect 21361 23273 21373 23307
rect 21407 23304 21419 23307
rect 21634 23304 21640 23316
rect 21407 23276 21640 23304
rect 21407 23273 21419 23276
rect 21361 23267 21419 23273
rect 21634 23264 21640 23276
rect 21692 23304 21698 23316
rect 23290 23304 23296 23316
rect 21692 23276 23296 23304
rect 21692 23264 21698 23276
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 23566 23264 23572 23316
rect 23624 23304 23630 23316
rect 23937 23307 23995 23313
rect 23937 23304 23949 23307
rect 23624 23276 23949 23304
rect 23624 23264 23630 23276
rect 15930 23196 15936 23248
rect 15988 23236 15994 23248
rect 16108 23239 16166 23245
rect 16108 23236 16120 23239
rect 15988 23208 16120 23236
rect 15988 23196 15994 23208
rect 16108 23205 16120 23208
rect 16154 23236 16166 23239
rect 16390 23236 16396 23248
rect 16154 23208 16396 23236
rect 16154 23205 16166 23208
rect 16108 23199 16166 23205
rect 16390 23196 16396 23208
rect 16448 23196 16454 23248
rect 17788 23236 17816 23264
rect 23860 23248 23888 23276
rect 23937 23273 23949 23276
rect 23983 23273 23995 23307
rect 24670 23304 24676 23316
rect 24631 23276 24676 23304
rect 23937 23267 23995 23273
rect 24670 23264 24676 23276
rect 24728 23264 24734 23316
rect 18570 23239 18628 23245
rect 18570 23236 18582 23239
rect 17788 23208 18582 23236
rect 18570 23205 18582 23208
rect 18616 23205 18628 23239
rect 18570 23199 18628 23205
rect 23842 23196 23848 23248
rect 23900 23196 23906 23248
rect 11054 23177 11060 23180
rect 11048 23168 11060 23177
rect 11015 23140 11060 23168
rect 11048 23131 11060 23140
rect 11054 23128 11060 23131
rect 11112 23128 11118 23180
rect 12894 23128 12900 23180
rect 12952 23168 12958 23180
rect 13446 23168 13452 23180
rect 12952 23140 13452 23168
rect 12952 23128 12958 23140
rect 13446 23128 13452 23140
rect 13504 23168 13510 23180
rect 13725 23171 13783 23177
rect 13725 23168 13737 23171
rect 13504 23140 13737 23168
rect 13504 23128 13510 23140
rect 13725 23137 13737 23140
rect 13771 23137 13783 23171
rect 13725 23131 13783 23137
rect 18325 23171 18383 23177
rect 18325 23137 18337 23171
rect 18371 23168 18383 23171
rect 18966 23168 18972 23180
rect 18371 23140 18972 23168
rect 18371 23137 18383 23140
rect 18325 23131 18383 23137
rect 18966 23128 18972 23140
rect 19024 23128 19030 23180
rect 21266 23168 21272 23180
rect 21227 23140 21272 23168
rect 21266 23128 21272 23140
rect 21324 23128 21330 23180
rect 24489 23171 24547 23177
rect 24489 23137 24501 23171
rect 24535 23168 24547 23171
rect 24762 23168 24768 23180
rect 24535 23140 24768 23168
rect 24535 23137 24547 23140
rect 24489 23131 24547 23137
rect 24762 23128 24768 23140
rect 24820 23128 24826 23180
rect 10778 23100 10784 23112
rect 10739 23072 10784 23100
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 13814 23100 13820 23112
rect 13775 23072 13820 23100
rect 13814 23060 13820 23072
rect 13872 23060 13878 23112
rect 14369 23103 14427 23109
rect 14369 23069 14381 23103
rect 14415 23100 14427 23103
rect 14458 23100 14464 23112
rect 14415 23072 14464 23100
rect 14415 23069 14427 23072
rect 14369 23063 14427 23069
rect 14458 23060 14464 23072
rect 14516 23060 14522 23112
rect 15838 23100 15844 23112
rect 15799 23072 15844 23100
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21453 23103 21511 23109
rect 21453 23100 21465 23103
rect 20864 23072 21465 23100
rect 20864 23060 20870 23072
rect 21453 23069 21465 23072
rect 21499 23069 21511 23103
rect 21453 23063 21511 23069
rect 22922 23060 22928 23112
rect 22980 23100 22986 23112
rect 23385 23103 23443 23109
rect 23385 23100 23397 23103
rect 22980 23072 23397 23100
rect 22980 23060 22986 23072
rect 23385 23069 23397 23072
rect 23431 23069 23443 23103
rect 23385 23063 23443 23069
rect 23569 23103 23627 23109
rect 23569 23069 23581 23103
rect 23615 23100 23627 23103
rect 23615 23072 24256 23100
rect 23615 23069 23627 23072
rect 23569 23063 23627 23069
rect 12434 22992 12440 23044
rect 12492 23032 12498 23044
rect 12805 23035 12863 23041
rect 12805 23032 12817 23035
rect 12492 23004 12817 23032
rect 12492 22992 12498 23004
rect 12805 23001 12817 23004
rect 12851 23032 12863 23035
rect 15856 23032 15884 23060
rect 12851 23004 15884 23032
rect 12851 23001 12863 23004
rect 12805 22995 12863 23001
rect 20714 22992 20720 23044
rect 20772 23032 20778 23044
rect 20901 23035 20959 23041
rect 20901 23032 20913 23035
rect 20772 23004 20913 23032
rect 20772 22992 20778 23004
rect 20901 23001 20913 23004
rect 20947 23001 20959 23035
rect 20901 22995 20959 23001
rect 24228 22976 24256 23072
rect 11790 22924 11796 22976
rect 11848 22964 11854 22976
rect 12161 22967 12219 22973
rect 12161 22964 12173 22967
rect 11848 22936 12173 22964
rect 11848 22924 11854 22936
rect 12161 22933 12173 22936
rect 12207 22933 12219 22967
rect 12161 22927 12219 22933
rect 13078 22924 13084 22976
rect 13136 22964 13142 22976
rect 13265 22967 13323 22973
rect 13265 22964 13277 22967
rect 13136 22936 13277 22964
rect 13136 22924 13142 22936
rect 13265 22933 13277 22936
rect 13311 22933 13323 22967
rect 13265 22927 13323 22933
rect 14826 22924 14832 22976
rect 14884 22964 14890 22976
rect 14921 22967 14979 22973
rect 14921 22964 14933 22967
rect 14884 22936 14933 22964
rect 14884 22924 14890 22936
rect 14921 22933 14933 22936
rect 14967 22964 14979 22967
rect 15286 22964 15292 22976
rect 14967 22936 15292 22964
rect 14967 22933 14979 22936
rect 14921 22927 14979 22933
rect 15286 22924 15292 22936
rect 15344 22924 15350 22976
rect 22462 22924 22468 22976
rect 22520 22964 22526 22976
rect 22925 22967 22983 22973
rect 22925 22964 22937 22967
rect 22520 22936 22937 22964
rect 22520 22924 22526 22936
rect 22925 22933 22937 22936
rect 22971 22933 22983 22967
rect 22925 22927 22983 22933
rect 24210 22924 24216 22976
rect 24268 22964 24274 22976
rect 24305 22967 24363 22973
rect 24305 22964 24317 22967
rect 24268 22936 24317 22964
rect 24268 22924 24274 22936
rect 24305 22933 24317 22936
rect 24351 22933 24363 22967
rect 24305 22927 24363 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 10778 22760 10784 22772
rect 10739 22732 10784 22760
rect 10778 22720 10784 22732
rect 10836 22720 10842 22772
rect 11054 22720 11060 22772
rect 11112 22760 11118 22772
rect 11241 22763 11299 22769
rect 11241 22760 11253 22763
rect 11112 22732 11253 22760
rect 11112 22720 11118 22732
rect 11241 22729 11253 22732
rect 11287 22760 11299 22763
rect 13814 22760 13820 22772
rect 11287 22732 13820 22760
rect 11287 22729 11299 22732
rect 11241 22723 11299 22729
rect 13814 22720 13820 22732
rect 13872 22760 13878 22772
rect 14369 22763 14427 22769
rect 14369 22760 14381 22763
rect 13872 22732 14381 22760
rect 13872 22720 13878 22732
rect 14369 22729 14381 22732
rect 14415 22729 14427 22763
rect 14369 22723 14427 22729
rect 15838 22720 15844 22772
rect 15896 22760 15902 22772
rect 15933 22763 15991 22769
rect 15933 22760 15945 22763
rect 15896 22732 15945 22760
rect 15896 22720 15902 22732
rect 15933 22729 15945 22732
rect 15979 22729 15991 22763
rect 16390 22760 16396 22772
rect 16351 22732 16396 22760
rect 15933 22723 15991 22729
rect 16390 22720 16396 22732
rect 16448 22720 16454 22772
rect 17034 22760 17040 22772
rect 16995 22732 17040 22760
rect 17034 22720 17040 22732
rect 17092 22720 17098 22772
rect 17494 22760 17500 22772
rect 17455 22732 17500 22760
rect 17494 22720 17500 22732
rect 17552 22720 17558 22772
rect 17770 22760 17776 22772
rect 17731 22732 17776 22760
rect 17770 22720 17776 22732
rect 17828 22720 17834 22772
rect 18046 22760 18052 22772
rect 18007 22732 18052 22760
rect 18046 22720 18052 22732
rect 18104 22720 18110 22772
rect 21545 22763 21603 22769
rect 21545 22729 21557 22763
rect 21591 22760 21603 22763
rect 21818 22760 21824 22772
rect 21591 22732 21824 22760
rect 21591 22729 21603 22732
rect 21545 22723 21603 22729
rect 21818 22720 21824 22732
rect 21876 22720 21882 22772
rect 22922 22760 22928 22772
rect 22883 22732 22928 22760
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 25406 22760 25412 22772
rect 25367 22732 25412 22760
rect 25406 22720 25412 22732
rect 25464 22720 25470 22772
rect 10796 22692 10824 22720
rect 11514 22692 11520 22704
rect 10796 22664 11520 22692
rect 11514 22652 11520 22664
rect 11572 22692 11578 22704
rect 12161 22695 12219 22701
rect 12161 22692 12173 22695
rect 11572 22664 12173 22692
rect 11572 22652 11578 22664
rect 12161 22661 12173 22664
rect 12207 22661 12219 22695
rect 17788 22692 17816 22720
rect 18414 22692 18420 22704
rect 17788 22664 18420 22692
rect 12161 22655 12219 22661
rect 12176 22624 12204 22655
rect 18414 22652 18420 22664
rect 18472 22692 18478 22704
rect 22649 22695 22707 22701
rect 18472 22664 18644 22692
rect 18472 22652 18478 22664
rect 12434 22624 12440 22636
rect 12176 22596 12440 22624
rect 12434 22584 12440 22596
rect 12492 22624 12498 22636
rect 15565 22627 15623 22633
rect 12492 22596 12537 22624
rect 12492 22584 12498 22596
rect 15565 22593 15577 22627
rect 15611 22624 15623 22627
rect 15654 22624 15660 22636
rect 15611 22596 15660 22624
rect 15611 22593 15623 22596
rect 15565 22587 15623 22593
rect 15654 22584 15660 22596
rect 15712 22584 15718 22636
rect 18138 22584 18144 22636
rect 18196 22624 18202 22636
rect 18616 22633 18644 22664
rect 22649 22661 22661 22695
rect 22695 22692 22707 22695
rect 23290 22692 23296 22704
rect 22695 22664 23296 22692
rect 22695 22661 22707 22664
rect 22649 22655 22707 22661
rect 23290 22652 23296 22664
rect 23348 22652 23354 22704
rect 18509 22627 18567 22633
rect 18509 22624 18521 22627
rect 18196 22596 18521 22624
rect 18196 22584 18202 22596
rect 18509 22593 18521 22596
rect 18555 22593 18567 22627
rect 18509 22587 18567 22593
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 21266 22584 21272 22636
rect 21324 22624 21330 22636
rect 22189 22627 22247 22633
rect 22189 22624 22201 22627
rect 21324 22596 22201 22624
rect 21324 22584 21330 22596
rect 22189 22593 22201 22596
rect 22235 22624 22247 22627
rect 23198 22624 23204 22636
rect 22235 22596 23204 22624
rect 22235 22593 22247 22596
rect 22189 22587 22247 22593
rect 23198 22584 23204 22596
rect 23256 22584 23262 22636
rect 23382 22584 23388 22636
rect 23440 22624 23446 22636
rect 24210 22624 24216 22636
rect 23440 22596 24216 22624
rect 23440 22584 23446 22596
rect 24210 22584 24216 22596
rect 24268 22584 24274 22636
rect 16853 22559 16911 22565
rect 16853 22525 16865 22559
rect 16899 22556 16911 22559
rect 17494 22556 17500 22568
rect 16899 22528 17500 22556
rect 16899 22525 16911 22528
rect 16853 22519 16911 22525
rect 17494 22516 17500 22528
rect 17552 22516 17558 22568
rect 18322 22516 18328 22568
rect 18380 22556 18386 22568
rect 18417 22559 18475 22565
rect 18417 22556 18429 22559
rect 18380 22528 18429 22556
rect 18380 22516 18386 22528
rect 18417 22525 18429 22528
rect 18463 22556 18475 22559
rect 19429 22559 19487 22565
rect 19429 22556 19441 22559
rect 18463 22528 19441 22556
rect 18463 22525 18475 22528
rect 18417 22519 18475 22525
rect 19429 22525 19441 22528
rect 19475 22525 19487 22559
rect 19429 22519 19487 22525
rect 20165 22559 20223 22565
rect 20165 22525 20177 22559
rect 20211 22525 20223 22559
rect 20165 22519 20223 22525
rect 12710 22497 12716 22500
rect 12704 22451 12716 22497
rect 12768 22488 12774 22500
rect 14829 22491 14887 22497
rect 12768 22460 12804 22488
rect 12710 22448 12716 22451
rect 12768 22448 12774 22460
rect 14829 22457 14841 22491
rect 14875 22488 14887 22491
rect 14875 22460 15424 22488
rect 14875 22457 14887 22460
rect 14829 22451 14887 22457
rect 15396 22432 15424 22460
rect 14918 22420 14924 22432
rect 14879 22392 14924 22420
rect 14918 22380 14924 22392
rect 14976 22380 14982 22432
rect 15286 22420 15292 22432
rect 15247 22392 15292 22420
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 15378 22380 15384 22432
rect 15436 22420 15442 22432
rect 15436 22392 15481 22420
rect 15436 22380 15442 22392
rect 18966 22380 18972 22432
rect 19024 22420 19030 22432
rect 19153 22423 19211 22429
rect 19153 22420 19165 22423
rect 19024 22392 19165 22420
rect 19024 22380 19030 22392
rect 19153 22389 19165 22392
rect 19199 22420 19211 22423
rect 20073 22423 20131 22429
rect 20073 22420 20085 22423
rect 19199 22392 20085 22420
rect 19199 22389 19211 22392
rect 19153 22383 19211 22389
rect 20073 22389 20085 22392
rect 20119 22420 20131 22423
rect 20180 22420 20208 22519
rect 23842 22516 23848 22568
rect 23900 22556 23906 22568
rect 24029 22559 24087 22565
rect 24029 22556 24041 22559
rect 23900 22528 24041 22556
rect 23900 22516 23906 22528
rect 24029 22525 24041 22528
rect 24075 22525 24087 22559
rect 24029 22519 24087 22525
rect 20254 22448 20260 22500
rect 20312 22488 20318 22500
rect 20410 22491 20468 22497
rect 20410 22488 20422 22491
rect 20312 22460 20422 22488
rect 20312 22448 20318 22460
rect 20410 22457 20422 22460
rect 20456 22457 20468 22491
rect 24121 22491 24179 22497
rect 24121 22488 24133 22491
rect 20410 22451 20468 22457
rect 23492 22460 24133 22488
rect 20714 22420 20720 22432
rect 20119 22392 20720 22420
rect 20119 22389 20131 22392
rect 20073 22383 20131 22389
rect 20714 22380 20720 22392
rect 20772 22380 20778 22432
rect 23290 22380 23296 22432
rect 23348 22420 23354 22432
rect 23492 22429 23520 22460
rect 24121 22457 24133 22460
rect 24167 22457 24179 22491
rect 24121 22451 24179 22457
rect 23477 22423 23535 22429
rect 23477 22420 23489 22423
rect 23348 22392 23489 22420
rect 23348 22380 23354 22392
rect 23477 22389 23489 22392
rect 23523 22389 23535 22423
rect 23658 22420 23664 22432
rect 23619 22392 23664 22420
rect 23477 22383 23535 22389
rect 23658 22380 23664 22392
rect 23716 22380 23722 22432
rect 24762 22420 24768 22432
rect 24723 22392 24768 22420
rect 24762 22380 24768 22392
rect 24820 22380 24826 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 11422 22216 11428 22228
rect 11383 22188 11428 22216
rect 11422 22176 11428 22188
rect 11480 22176 11486 22228
rect 12894 22216 12900 22228
rect 12855 22188 12900 22216
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 13265 22219 13323 22225
rect 13265 22185 13277 22219
rect 13311 22216 13323 22219
rect 14918 22216 14924 22228
rect 13311 22188 14924 22216
rect 13311 22185 13323 22188
rect 13265 22179 13323 22185
rect 13280 22148 13308 22179
rect 14918 22176 14924 22188
rect 14976 22176 14982 22228
rect 17313 22219 17371 22225
rect 17313 22185 17325 22219
rect 17359 22216 17371 22219
rect 17402 22216 17408 22228
rect 17359 22188 17408 22216
rect 17359 22185 17371 22188
rect 17313 22179 17371 22185
rect 17402 22176 17408 22188
rect 17460 22176 17466 22228
rect 18414 22216 18420 22228
rect 18375 22188 18420 22216
rect 18414 22176 18420 22188
rect 18472 22176 18478 22228
rect 18506 22176 18512 22228
rect 18564 22216 18570 22228
rect 18874 22216 18880 22228
rect 18564 22188 18880 22216
rect 18564 22176 18570 22188
rect 18874 22176 18880 22188
rect 18932 22176 18938 22228
rect 20254 22216 20260 22228
rect 20215 22188 20260 22216
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 20717 22219 20775 22225
rect 20717 22185 20729 22219
rect 20763 22216 20775 22219
rect 20806 22216 20812 22228
rect 20763 22188 20812 22216
rect 20763 22185 20775 22188
rect 20717 22179 20775 22185
rect 20806 22176 20812 22188
rect 20864 22176 20870 22228
rect 21634 22216 21640 22228
rect 21595 22188 21640 22216
rect 21634 22176 21640 22188
rect 21692 22176 21698 22228
rect 22649 22219 22707 22225
rect 22649 22185 22661 22219
rect 22695 22216 22707 22219
rect 23017 22219 23075 22225
rect 23017 22216 23029 22219
rect 22695 22188 23029 22216
rect 22695 22185 22707 22188
rect 22649 22179 22707 22185
rect 23017 22185 23029 22188
rect 23063 22216 23075 22219
rect 23382 22216 23388 22228
rect 23063 22188 23388 22216
rect 23063 22185 23075 22188
rect 23017 22179 23075 22185
rect 23382 22176 23388 22188
rect 23440 22176 23446 22228
rect 23658 22148 23664 22160
rect 12360 22120 13308 22148
rect 23216 22120 23664 22148
rect 12161 22083 12219 22089
rect 12161 22049 12173 22083
rect 12207 22080 12219 22083
rect 12360 22080 12388 22120
rect 12207 22052 12388 22080
rect 12529 22083 12587 22089
rect 12207 22049 12219 22052
rect 12161 22043 12219 22049
rect 12529 22049 12541 22083
rect 12575 22080 12587 22083
rect 12710 22080 12716 22092
rect 12575 22052 12716 22080
rect 12575 22049 12587 22052
rect 12529 22043 12587 22049
rect 12710 22040 12716 22052
rect 12768 22080 12774 22092
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 12768 22052 13584 22080
rect 12768 22040 12774 22052
rect 11054 21972 11060 22024
rect 11112 22012 11118 22024
rect 11517 22015 11575 22021
rect 11517 22012 11529 22015
rect 11112 21984 11529 22012
rect 11112 21972 11118 21984
rect 11517 21981 11529 21984
rect 11563 21981 11575 22015
rect 11517 21975 11575 21981
rect 11701 22015 11759 22021
rect 11701 21981 11713 22015
rect 11747 22012 11759 22015
rect 11790 22012 11796 22024
rect 11747 21984 11796 22012
rect 11747 21981 11759 21984
rect 11701 21975 11759 21981
rect 11790 21972 11796 21984
rect 11848 21972 11854 22024
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 13354 22012 13360 22024
rect 12492 21984 13360 22012
rect 12492 21972 12498 21984
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 13556 22021 13584 22052
rect 15672 22052 15761 22080
rect 15672 22024 15700 22052
rect 15749 22049 15761 22052
rect 15795 22049 15807 22083
rect 20993 22083 21051 22089
rect 15749 22043 15807 22049
rect 17696 22052 19104 22080
rect 17696 22024 17724 22052
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 13722 22012 13728 22024
rect 13587 21984 13728 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 13722 21972 13728 21984
rect 13780 21972 13786 22024
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 22012 15071 22015
rect 15286 22012 15292 22024
rect 15059 21984 15292 22012
rect 15059 21981 15071 21984
rect 15013 21975 15071 21981
rect 15286 21972 15292 21984
rect 15344 21972 15350 22024
rect 15654 21972 15660 22024
rect 15712 21972 15718 22024
rect 15838 22012 15844 22024
rect 15799 21984 15844 22012
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 15930 21972 15936 22024
rect 15988 22012 15994 22024
rect 15988 21984 16033 22012
rect 15988 21972 15994 21984
rect 16666 21972 16672 22024
rect 16724 22012 16730 22024
rect 17405 22015 17463 22021
rect 17405 22012 17417 22015
rect 16724 21984 17417 22012
rect 16724 21972 16730 21984
rect 17405 21981 17417 21984
rect 17451 21981 17463 22015
rect 17405 21975 17463 21981
rect 17589 22015 17647 22021
rect 17589 21981 17601 22015
rect 17635 22012 17647 22015
rect 17678 22012 17684 22024
rect 17635 21984 17684 22012
rect 17635 21981 17647 21984
rect 17589 21975 17647 21981
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 18414 21972 18420 22024
rect 18472 22012 18478 22024
rect 19076 22021 19104 22052
rect 20993 22049 21005 22083
rect 21039 22080 21051 22083
rect 21039 22052 21128 22080
rect 21039 22049 21051 22052
rect 20993 22043 21051 22049
rect 18969 22015 19027 22021
rect 18969 22012 18981 22015
rect 18472 21984 18981 22012
rect 18472 21972 18478 21984
rect 18969 21981 18981 21984
rect 19015 21981 19027 22015
rect 18969 21975 19027 21981
rect 19061 22015 19119 22021
rect 19061 21981 19073 22015
rect 19107 21981 19119 22015
rect 19061 21975 19119 21981
rect 15381 21947 15439 21953
rect 15381 21913 15393 21947
rect 15427 21944 15439 21947
rect 16022 21944 16028 21956
rect 15427 21916 16028 21944
rect 15427 21913 15439 21916
rect 15381 21907 15439 21913
rect 16022 21904 16028 21916
rect 16080 21904 16086 21956
rect 18984 21944 19012 21975
rect 21100 21956 21128 22052
rect 22094 22040 22100 22092
rect 22152 22080 22158 22092
rect 23216 22080 23244 22120
rect 23658 22108 23664 22120
rect 23716 22108 23722 22160
rect 23382 22089 23388 22092
rect 23376 22080 23388 22089
rect 22152 22052 22197 22080
rect 22572 22052 23244 22080
rect 23343 22052 23388 22080
rect 22152 22040 22158 22052
rect 22005 22015 22063 22021
rect 22005 21981 22017 22015
rect 22051 22012 22063 22015
rect 22370 22012 22376 22024
rect 22051 21984 22376 22012
rect 22051 21981 22063 21984
rect 22005 21975 22063 21981
rect 22370 21972 22376 21984
rect 22428 22012 22434 22024
rect 22572 22012 22600 22052
rect 23376 22043 23388 22052
rect 23382 22040 23388 22043
rect 23440 22040 23446 22092
rect 23106 22012 23112 22024
rect 22428 21984 22600 22012
rect 23067 21984 23112 22012
rect 22428 21972 22434 21984
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 19150 21944 19156 21956
rect 18984 21916 19156 21944
rect 19150 21904 19156 21916
rect 19208 21904 19214 21956
rect 21082 21904 21088 21956
rect 21140 21904 21146 21956
rect 21177 21947 21235 21953
rect 21177 21913 21189 21947
rect 21223 21944 21235 21947
rect 21910 21944 21916 21956
rect 21223 21916 21916 21944
rect 21223 21913 21235 21916
rect 21177 21907 21235 21913
rect 21910 21904 21916 21916
rect 21968 21904 21974 21956
rect 11057 21879 11115 21885
rect 11057 21845 11069 21879
rect 11103 21876 11115 21879
rect 12342 21876 12348 21888
rect 11103 21848 12348 21876
rect 11103 21845 11115 21848
rect 11057 21839 11115 21845
rect 12342 21836 12348 21848
rect 12400 21836 12406 21888
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 13909 21879 13967 21885
rect 13909 21876 13921 21879
rect 13504 21848 13921 21876
rect 13504 21836 13510 21848
rect 13909 21845 13921 21848
rect 13955 21845 13967 21879
rect 16390 21876 16396 21888
rect 16351 21848 16396 21876
rect 13909 21839 13967 21845
rect 16390 21836 16396 21848
rect 16448 21836 16454 21888
rect 16942 21876 16948 21888
rect 16903 21848 16948 21876
rect 16942 21836 16948 21848
rect 17000 21836 17006 21888
rect 17586 21836 17592 21888
rect 17644 21876 17650 21888
rect 18509 21879 18567 21885
rect 18509 21876 18521 21879
rect 17644 21848 18521 21876
rect 17644 21836 17650 21848
rect 18509 21845 18521 21848
rect 18555 21845 18567 21879
rect 19518 21876 19524 21888
rect 19479 21848 19524 21876
rect 18509 21839 18567 21845
rect 19518 21836 19524 21848
rect 19576 21836 19582 21888
rect 22281 21879 22339 21885
rect 22281 21845 22293 21879
rect 22327 21876 22339 21879
rect 23290 21876 23296 21888
rect 22327 21848 23296 21876
rect 22327 21845 22339 21848
rect 22281 21839 22339 21845
rect 23290 21836 23296 21848
rect 23348 21836 23354 21888
rect 24210 21836 24216 21888
rect 24268 21876 24274 21888
rect 24489 21879 24547 21885
rect 24489 21876 24501 21879
rect 24268 21848 24501 21876
rect 24268 21836 24274 21848
rect 24489 21845 24501 21848
rect 24535 21845 24547 21879
rect 24489 21839 24547 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 11054 21672 11060 21684
rect 11015 21644 11060 21672
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 13722 21672 13728 21684
rect 13587 21644 13728 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 15838 21632 15844 21684
rect 15896 21672 15902 21684
rect 15933 21675 15991 21681
rect 15933 21672 15945 21675
rect 15896 21644 15945 21672
rect 15896 21632 15902 21644
rect 15933 21641 15945 21644
rect 15979 21672 15991 21675
rect 16022 21672 16028 21684
rect 15979 21644 16028 21672
rect 15979 21641 15991 21644
rect 15933 21635 15991 21641
rect 16022 21632 16028 21644
rect 16080 21632 16086 21684
rect 16577 21675 16635 21681
rect 16577 21641 16589 21675
rect 16623 21672 16635 21675
rect 17310 21672 17316 21684
rect 16623 21644 17316 21672
rect 16623 21641 16635 21644
rect 16577 21635 16635 21641
rect 17310 21632 17316 21644
rect 17368 21632 17374 21684
rect 18877 21675 18935 21681
rect 18877 21641 18889 21675
rect 18923 21672 18935 21675
rect 18966 21672 18972 21684
rect 18923 21644 18972 21672
rect 18923 21641 18935 21644
rect 18877 21635 18935 21641
rect 18966 21632 18972 21644
rect 19024 21632 19030 21684
rect 20254 21632 20260 21684
rect 20312 21672 20318 21684
rect 20349 21675 20407 21681
rect 20349 21672 20361 21675
rect 20312 21644 20361 21672
rect 20312 21632 20318 21644
rect 20349 21641 20361 21644
rect 20395 21641 20407 21675
rect 20349 21635 20407 21641
rect 22005 21675 22063 21681
rect 22005 21641 22017 21675
rect 22051 21672 22063 21675
rect 22094 21672 22100 21684
rect 22051 21644 22100 21672
rect 22051 21641 22063 21644
rect 22005 21635 22063 21641
rect 22094 21632 22100 21644
rect 22152 21632 22158 21684
rect 12158 21564 12164 21616
rect 12216 21604 12222 21616
rect 12216 21576 13032 21604
rect 12216 21564 12222 21576
rect 11330 21496 11336 21548
rect 11388 21536 11394 21548
rect 11514 21536 11520 21548
rect 11388 21508 11520 21536
rect 11388 21496 11394 21508
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 13004 21545 13032 21576
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 14369 21539 14427 21545
rect 14369 21505 14381 21539
rect 14415 21536 14427 21539
rect 15381 21539 15439 21545
rect 15381 21536 15393 21539
rect 14415 21508 15393 21536
rect 14415 21505 14427 21508
rect 14369 21499 14427 21505
rect 15381 21505 15393 21508
rect 15427 21536 15439 21539
rect 15838 21536 15844 21548
rect 15427 21508 15844 21536
rect 15427 21505 15439 21508
rect 15381 21499 15439 21505
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 16945 21539 17003 21545
rect 16945 21536 16957 21539
rect 16632 21508 16957 21536
rect 16632 21496 16638 21508
rect 16945 21505 16957 21508
rect 16991 21505 17003 21539
rect 16945 21499 17003 21505
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18984 21545 19012 21632
rect 21913 21607 21971 21613
rect 21913 21573 21925 21607
rect 21959 21604 21971 21607
rect 21959 21576 22600 21604
rect 21959 21573 21971 21576
rect 21913 21567 21971 21573
rect 18969 21539 19027 21545
rect 18969 21536 18981 21539
rect 18104 21508 18981 21536
rect 18104 21496 18110 21508
rect 18969 21505 18981 21508
rect 19015 21505 19027 21539
rect 18969 21499 19027 21505
rect 21545 21539 21603 21545
rect 21545 21505 21557 21539
rect 21591 21536 21603 21539
rect 22462 21536 22468 21548
rect 21591 21508 22468 21536
rect 21591 21505 21603 21508
rect 21545 21499 21603 21505
rect 22462 21496 22468 21508
rect 22520 21496 22526 21548
rect 22572 21545 22600 21576
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21536 22615 21539
rect 23750 21536 23756 21548
rect 22603 21508 23756 21536
rect 22603 21505 22615 21508
rect 22557 21499 22615 21505
rect 23750 21496 23756 21508
rect 23808 21536 23814 21548
rect 23808 21508 24256 21536
rect 23808 21496 23814 21508
rect 24228 21480 24256 21508
rect 14737 21471 14795 21477
rect 14737 21437 14749 21471
rect 14783 21468 14795 21471
rect 15194 21468 15200 21480
rect 14783 21440 15200 21468
rect 14783 21437 14795 21440
rect 14737 21431 14795 21437
rect 15194 21428 15200 21440
rect 15252 21428 15258 21480
rect 16390 21468 16396 21480
rect 16351 21440 16396 21468
rect 16390 21428 16396 21440
rect 16448 21428 16454 21480
rect 19236 21471 19294 21477
rect 19236 21437 19248 21471
rect 19282 21468 19294 21471
rect 19518 21468 19524 21480
rect 19282 21440 19524 21468
rect 19282 21437 19294 21440
rect 19236 21431 19294 21437
rect 19518 21428 19524 21440
rect 19576 21428 19582 21480
rect 22370 21468 22376 21480
rect 22331 21440 22376 21468
rect 22370 21428 22376 21440
rect 22428 21428 22434 21480
rect 24121 21471 24179 21477
rect 24121 21468 24133 21471
rect 23952 21440 24133 21468
rect 10781 21403 10839 21409
rect 10781 21369 10793 21403
rect 10827 21400 10839 21403
rect 12526 21400 12532 21412
rect 10827 21372 12532 21400
rect 10827 21369 10839 21372
rect 10781 21363 10839 21369
rect 12526 21360 12532 21372
rect 12584 21400 12590 21412
rect 12897 21403 12955 21409
rect 12897 21400 12909 21403
rect 12584 21372 12909 21400
rect 12584 21360 12590 21372
rect 12897 21369 12909 21372
rect 12943 21369 12955 21403
rect 15289 21403 15347 21409
rect 15289 21400 15301 21403
rect 12897 21363 12955 21369
rect 13924 21372 15301 21400
rect 11514 21332 11520 21344
rect 11475 21304 11520 21332
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 11790 21332 11796 21344
rect 11751 21304 11796 21332
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 12158 21332 12164 21344
rect 12119 21304 12164 21332
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 12437 21335 12495 21341
rect 12437 21301 12449 21335
rect 12483 21332 12495 21335
rect 12618 21332 12624 21344
rect 12483 21304 12624 21332
rect 12483 21301 12495 21304
rect 12437 21295 12495 21301
rect 12618 21292 12624 21304
rect 12676 21292 12682 21344
rect 12802 21332 12808 21344
rect 12763 21304 12808 21332
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 13924 21341 13952 21372
rect 15289 21369 15301 21372
rect 15335 21369 15347 21403
rect 17402 21400 17408 21412
rect 17315 21372 17408 21400
rect 15289 21363 15347 21369
rect 17402 21360 17408 21372
rect 17460 21400 17466 21412
rect 17862 21400 17868 21412
rect 17460 21372 17868 21400
rect 17460 21360 17466 21372
rect 17862 21360 17868 21372
rect 17920 21360 17926 21412
rect 13909 21335 13967 21341
rect 13909 21332 13921 21335
rect 13872 21304 13921 21332
rect 13872 21292 13878 21304
rect 13909 21301 13921 21304
rect 13955 21301 13967 21335
rect 13909 21295 13967 21301
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 14792 21304 14841 21332
rect 14792 21292 14798 21304
rect 14829 21301 14841 21304
rect 14875 21301 14887 21335
rect 14829 21295 14887 21301
rect 15746 21292 15752 21344
rect 15804 21332 15810 21344
rect 16209 21335 16267 21341
rect 16209 21332 16221 21335
rect 15804 21304 16221 21332
rect 15804 21292 15810 21304
rect 16209 21301 16221 21304
rect 16255 21301 16267 21335
rect 16209 21295 16267 21301
rect 17034 21292 17040 21344
rect 17092 21332 17098 21344
rect 17678 21332 17684 21344
rect 17092 21304 17684 21332
rect 17092 21292 17098 21304
rect 17678 21292 17684 21304
rect 17736 21332 17742 21344
rect 17773 21335 17831 21341
rect 17773 21332 17785 21335
rect 17736 21304 17785 21332
rect 17736 21292 17742 21304
rect 17773 21301 17785 21304
rect 17819 21301 17831 21335
rect 17773 21295 17831 21301
rect 17954 21292 17960 21344
rect 18012 21332 18018 21344
rect 18414 21332 18420 21344
rect 18012 21304 18420 21332
rect 18012 21292 18018 21304
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 21085 21335 21143 21341
rect 21085 21301 21097 21335
rect 21131 21332 21143 21335
rect 21174 21332 21180 21344
rect 21131 21304 21180 21332
rect 21131 21301 21143 21304
rect 21085 21295 21143 21301
rect 21174 21292 21180 21304
rect 21232 21292 21238 21344
rect 23106 21292 23112 21344
rect 23164 21332 23170 21344
rect 23201 21335 23259 21341
rect 23201 21332 23213 21335
rect 23164 21304 23213 21332
rect 23164 21292 23170 21304
rect 23201 21301 23213 21304
rect 23247 21332 23259 21335
rect 23842 21332 23848 21344
rect 23247 21304 23848 21332
rect 23247 21301 23259 21304
rect 23201 21295 23259 21301
rect 23842 21292 23848 21304
rect 23900 21332 23906 21344
rect 23952 21341 23980 21440
rect 24121 21437 24133 21440
rect 24167 21437 24179 21471
rect 24121 21431 24179 21437
rect 24210 21428 24216 21480
rect 24268 21468 24274 21480
rect 24377 21471 24435 21477
rect 24377 21468 24389 21471
rect 24268 21440 24389 21468
rect 24268 21428 24274 21440
rect 24377 21437 24389 21440
rect 24423 21437 24435 21471
rect 24377 21431 24435 21437
rect 23937 21335 23995 21341
rect 23937 21332 23949 21335
rect 23900 21304 23949 21332
rect 23900 21292 23906 21304
rect 23937 21301 23949 21304
rect 23983 21301 23995 21335
rect 25498 21332 25504 21344
rect 25459 21304 25504 21332
rect 23937 21295 23995 21301
rect 25498 21292 25504 21304
rect 25556 21292 25562 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 13354 21088 13360 21140
rect 13412 21128 13418 21140
rect 13449 21131 13507 21137
rect 13449 21128 13461 21131
rect 13412 21100 13461 21128
rect 13412 21088 13418 21100
rect 13449 21097 13461 21100
rect 13495 21097 13507 21131
rect 13449 21091 13507 21097
rect 14001 21131 14059 21137
rect 14001 21097 14013 21131
rect 14047 21128 14059 21131
rect 14826 21128 14832 21140
rect 14047 21100 14832 21128
rect 14047 21097 14059 21100
rect 14001 21091 14059 21097
rect 14826 21088 14832 21100
rect 14884 21088 14890 21140
rect 15105 21131 15163 21137
rect 15105 21097 15117 21131
rect 15151 21128 15163 21131
rect 15930 21128 15936 21140
rect 15151 21100 15936 21128
rect 15151 21097 15163 21100
rect 15105 21091 15163 21097
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 16942 21088 16948 21140
rect 17000 21128 17006 21140
rect 17678 21128 17684 21140
rect 17000 21100 17684 21128
rect 17000 21088 17006 21100
rect 17678 21088 17684 21100
rect 17736 21088 17742 21140
rect 18601 21131 18659 21137
rect 18601 21097 18613 21131
rect 18647 21128 18659 21131
rect 18874 21128 18880 21140
rect 18647 21100 18880 21128
rect 18647 21097 18659 21100
rect 18601 21091 18659 21097
rect 18874 21088 18880 21100
rect 18932 21088 18938 21140
rect 21729 21131 21787 21137
rect 21729 21097 21741 21131
rect 21775 21128 21787 21131
rect 22094 21128 22100 21140
rect 21775 21100 22100 21128
rect 21775 21097 21787 21100
rect 21729 21091 21787 21097
rect 22094 21088 22100 21100
rect 22152 21088 22158 21140
rect 23201 21131 23259 21137
rect 23201 21097 23213 21131
rect 23247 21128 23259 21131
rect 23382 21128 23388 21140
rect 23247 21100 23388 21128
rect 23247 21097 23259 21100
rect 23201 21091 23259 21097
rect 23382 21088 23388 21100
rect 23440 21088 23446 21140
rect 23750 21128 23756 21140
rect 23711 21100 23756 21128
rect 23750 21088 23756 21100
rect 23808 21088 23814 21140
rect 15378 21020 15384 21072
rect 15436 21060 15442 21072
rect 15749 21063 15807 21069
rect 15749 21060 15761 21063
rect 15436 21032 15761 21060
rect 15436 21020 15442 21032
rect 15749 21029 15761 21032
rect 15795 21029 15807 21063
rect 15749 21023 15807 21029
rect 16669 21063 16727 21069
rect 16669 21029 16681 21063
rect 16715 21060 16727 21063
rect 17586 21060 17592 21072
rect 16715 21032 17592 21060
rect 16715 21029 16727 21032
rect 16669 21023 16727 21029
rect 17586 21020 17592 21032
rect 17644 21020 17650 21072
rect 19518 21060 19524 21072
rect 18340 21032 19524 21060
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 1946 20992 1952 21004
rect 1443 20964 1952 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 1946 20952 1952 20964
rect 2004 20952 2010 21004
rect 11238 20952 11244 21004
rect 11296 20992 11302 21004
rect 11790 21001 11796 21004
rect 11773 20995 11796 21001
rect 11773 20992 11785 20995
rect 11296 20964 11785 20992
rect 11296 20952 11302 20964
rect 11773 20961 11785 20964
rect 11848 20992 11854 21004
rect 15654 20992 15660 21004
rect 11848 20964 11921 20992
rect 15615 20964 15660 20992
rect 11773 20955 11796 20961
rect 11790 20952 11796 20955
rect 11848 20952 11854 20964
rect 15654 20952 15660 20964
rect 15712 20952 15718 21004
rect 11330 20884 11336 20936
rect 11388 20924 11394 20936
rect 11517 20927 11575 20933
rect 11517 20924 11529 20927
rect 11388 20896 11529 20924
rect 11388 20884 11394 20896
rect 11517 20893 11529 20896
rect 11563 20893 11575 20927
rect 15838 20924 15844 20936
rect 15799 20896 15844 20924
rect 11517 20887 11575 20893
rect 15838 20884 15844 20896
rect 15896 20884 15902 20936
rect 17865 20927 17923 20933
rect 17865 20893 17877 20927
rect 17911 20924 17923 20927
rect 18340 20924 18368 21032
rect 19518 21020 19524 21032
rect 19576 21020 19582 21072
rect 20714 21020 20720 21072
rect 20772 21060 20778 21072
rect 20898 21060 20904 21072
rect 20772 21032 20904 21060
rect 20772 21020 20778 21032
rect 20898 21020 20904 21032
rect 20956 21060 20962 21072
rect 23106 21060 23112 21072
rect 20956 21032 23112 21060
rect 20956 21020 20962 21032
rect 21836 21004 21864 21032
rect 23106 21020 23112 21032
rect 23164 21020 23170 21072
rect 23566 21020 23572 21072
rect 23624 21060 23630 21072
rect 24026 21060 24032 21072
rect 23624 21032 24032 21060
rect 23624 21020 23630 21032
rect 24026 21020 24032 21032
rect 24084 21020 24090 21072
rect 19150 20992 19156 21004
rect 19111 20964 19156 20992
rect 19150 20952 19156 20964
rect 19208 20992 19214 21004
rect 19797 20995 19855 21001
rect 19797 20992 19809 20995
rect 19208 20964 19809 20992
rect 19208 20952 19214 20964
rect 19797 20961 19809 20964
rect 19843 20961 19855 20995
rect 21818 20992 21824 21004
rect 21731 20964 21824 20992
rect 19797 20955 19855 20961
rect 21818 20952 21824 20964
rect 21876 20992 21882 21004
rect 22094 21001 22100 21004
rect 21876 20964 21901 20992
rect 21876 20952 21882 20964
rect 22088 20955 22100 21001
rect 22152 20992 22158 21004
rect 22152 20964 22188 20992
rect 22094 20952 22100 20955
rect 22152 20952 22158 20964
rect 23474 20952 23480 21004
rect 23532 20992 23538 21004
rect 24670 20992 24676 21004
rect 23532 20964 24676 20992
rect 23532 20952 23538 20964
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 17911 20896 18368 20924
rect 18432 20896 19257 20924
rect 17911 20893 17923 20896
rect 17865 20887 17923 20893
rect 1578 20856 1584 20868
rect 1539 20828 1584 20856
rect 1578 20816 1584 20828
rect 1636 20816 1642 20868
rect 12802 20816 12808 20868
rect 12860 20856 12866 20868
rect 13817 20859 13875 20865
rect 13817 20856 13829 20859
rect 12860 20828 13829 20856
rect 12860 20816 12866 20828
rect 13817 20825 13829 20828
rect 13863 20825 13875 20859
rect 13817 20819 13875 20825
rect 18432 20800 18460 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20924 19487 20927
rect 20254 20924 20260 20936
rect 19475 20896 20260 20924
rect 19475 20893 19487 20896
rect 19429 20887 19487 20893
rect 20254 20884 20260 20896
rect 20312 20884 20318 20936
rect 24210 20884 24216 20936
rect 24268 20924 24274 20936
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 24268 20896 24777 20924
rect 24268 20884 24274 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20924 25007 20927
rect 25498 20924 25504 20936
rect 24995 20896 25504 20924
rect 24995 20893 25007 20896
rect 24949 20887 25007 20893
rect 12894 20788 12900 20800
rect 12855 20760 12900 20788
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 14737 20791 14795 20797
rect 14737 20757 14749 20791
rect 14783 20788 14795 20791
rect 14826 20788 14832 20800
rect 14783 20760 14832 20788
rect 14783 20757 14795 20760
rect 14737 20751 14795 20757
rect 14826 20748 14832 20760
rect 14884 20748 14890 20800
rect 15286 20788 15292 20800
rect 15247 20760 15292 20788
rect 15286 20748 15292 20760
rect 15344 20748 15350 20800
rect 17034 20788 17040 20800
rect 16995 20760 17040 20788
rect 17034 20748 17040 20760
rect 17092 20748 17098 20800
rect 17221 20791 17279 20797
rect 17221 20757 17233 20791
rect 17267 20788 17279 20791
rect 18414 20788 18420 20800
rect 17267 20760 18420 20788
rect 17267 20757 17279 20760
rect 17221 20751 17279 20757
rect 18414 20748 18420 20760
rect 18472 20748 18478 20800
rect 18782 20788 18788 20800
rect 18743 20760 18788 20788
rect 18782 20748 18788 20760
rect 18840 20748 18846 20800
rect 20438 20748 20444 20800
rect 20496 20788 20502 20800
rect 20533 20791 20591 20797
rect 20533 20788 20545 20791
rect 20496 20760 20545 20788
rect 20496 20748 20502 20760
rect 20533 20757 20545 20760
rect 20579 20757 20591 20791
rect 24118 20788 24124 20800
rect 24079 20760 24124 20788
rect 20533 20751 20591 20757
rect 24118 20748 24124 20760
rect 24176 20748 24182 20800
rect 24210 20748 24216 20800
rect 24268 20788 24274 20800
rect 24305 20791 24363 20797
rect 24305 20788 24317 20791
rect 24268 20760 24317 20788
rect 24268 20748 24274 20760
rect 24305 20757 24317 20760
rect 24351 20757 24363 20791
rect 24780 20788 24808 20887
rect 25498 20884 25504 20896
rect 25556 20884 25562 20936
rect 24946 20788 24952 20800
rect 24780 20760 24952 20788
rect 24305 20751 24363 20757
rect 24946 20748 24952 20760
rect 25004 20748 25010 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 11238 20584 11244 20596
rect 11199 20556 11244 20584
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 11330 20544 11336 20596
rect 11388 20584 11394 20596
rect 11793 20587 11851 20593
rect 11793 20584 11805 20587
rect 11388 20556 11805 20584
rect 11388 20544 11394 20556
rect 11793 20553 11805 20556
rect 11839 20553 11851 20587
rect 11793 20547 11851 20553
rect 12437 20587 12495 20593
rect 12437 20553 12449 20587
rect 12483 20584 12495 20587
rect 12526 20584 12532 20596
rect 12483 20556 12532 20584
rect 12483 20553 12495 20556
rect 12437 20547 12495 20553
rect 10042 20476 10048 20528
rect 10100 20516 10106 20528
rect 11348 20516 11376 20544
rect 10100 20488 11376 20516
rect 11808 20516 11836 20547
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16025 20587 16083 20593
rect 16025 20584 16037 20587
rect 15896 20556 16037 20584
rect 15896 20544 15902 20556
rect 16025 20553 16037 20556
rect 16071 20584 16083 20587
rect 16945 20587 17003 20593
rect 16945 20584 16957 20587
rect 16071 20556 16957 20584
rect 16071 20553 16083 20556
rect 16025 20547 16083 20553
rect 16945 20553 16957 20556
rect 16991 20553 17003 20587
rect 16945 20547 17003 20553
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 19518 20584 19524 20596
rect 19475 20556 19524 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 20073 20587 20131 20593
rect 20073 20553 20085 20587
rect 20119 20584 20131 20587
rect 20254 20584 20260 20596
rect 20119 20556 20260 20584
rect 20119 20553 20131 20556
rect 20073 20547 20131 20553
rect 20254 20544 20260 20556
rect 20312 20544 20318 20596
rect 21818 20584 21824 20596
rect 21779 20556 21824 20584
rect 21818 20544 21824 20556
rect 21876 20544 21882 20596
rect 22094 20544 22100 20596
rect 22152 20584 22158 20596
rect 22189 20587 22247 20593
rect 22189 20584 22201 20587
rect 22152 20556 22201 20584
rect 22152 20544 22158 20556
rect 22189 20553 22201 20556
rect 22235 20553 22247 20587
rect 23474 20584 23480 20596
rect 23435 20556 23480 20584
rect 22189 20547 22247 20553
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 25498 20584 25504 20596
rect 25459 20556 25504 20584
rect 25498 20544 25504 20556
rect 25556 20584 25562 20596
rect 25869 20587 25927 20593
rect 25869 20584 25881 20587
rect 25556 20556 25881 20584
rect 25556 20544 25562 20556
rect 25869 20553 25881 20556
rect 25915 20553 25927 20587
rect 25869 20547 25927 20553
rect 13354 20516 13360 20528
rect 11808 20488 13360 20516
rect 10100 20476 10106 20488
rect 13354 20476 13360 20488
rect 13412 20476 13418 20528
rect 16574 20516 16580 20528
rect 16535 20488 16580 20516
rect 16574 20476 16580 20488
rect 16632 20476 16638 20528
rect 10318 20448 10324 20460
rect 10279 20420 10324 20448
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 12894 20408 12900 20460
rect 12952 20448 12958 20460
rect 12989 20451 13047 20457
rect 12989 20448 13001 20451
rect 12952 20420 13001 20448
rect 12952 20408 12958 20420
rect 12989 20417 13001 20420
rect 13035 20448 13047 20451
rect 13449 20451 13507 20457
rect 13449 20448 13461 20451
rect 13035 20420 13461 20448
rect 13035 20417 13047 20420
rect 12989 20411 13047 20417
rect 13449 20417 13461 20420
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 17865 20451 17923 20457
rect 17865 20417 17877 20451
rect 17911 20448 17923 20451
rect 18046 20448 18052 20460
rect 17911 20420 18052 20448
rect 17911 20417 17923 20420
rect 17865 20411 17923 20417
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 21085 20451 21143 20457
rect 21085 20448 21097 20451
rect 20772 20420 21097 20448
rect 20772 20408 20778 20420
rect 21085 20417 21097 20420
rect 21131 20417 21143 20451
rect 21085 20411 21143 20417
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20448 24823 20451
rect 25038 20448 25044 20460
rect 24811 20420 25044 20448
rect 24811 20417 24823 20420
rect 24765 20411 24823 20417
rect 25038 20408 25044 20420
rect 25096 20448 25102 20460
rect 25516 20448 25544 20544
rect 25096 20420 25544 20448
rect 25096 20408 25102 20420
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 14642 20380 14648 20392
rect 14603 20352 14648 20380
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 20441 20383 20499 20389
rect 20441 20349 20453 20383
rect 20487 20380 20499 20383
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20487 20352 21005 20380
rect 20487 20349 20499 20352
rect 20441 20343 20499 20349
rect 20993 20349 21005 20352
rect 21039 20380 21051 20383
rect 21634 20380 21640 20392
rect 21039 20352 21640 20380
rect 21039 20349 21051 20352
rect 20993 20343 21051 20349
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20380 22615 20383
rect 24118 20380 24124 20392
rect 22603 20352 24124 20380
rect 22603 20349 22615 20352
rect 22557 20343 22615 20349
rect 24118 20340 24124 20352
rect 24176 20380 24182 20392
rect 24489 20383 24547 20389
rect 24489 20380 24501 20383
rect 24176 20352 24501 20380
rect 24176 20340 24182 20352
rect 24489 20349 24501 20352
rect 24535 20349 24547 20383
rect 24489 20343 24547 20349
rect 12526 20272 12532 20324
rect 12584 20312 12590 20324
rect 12897 20315 12955 20321
rect 12897 20312 12909 20315
rect 12584 20284 12909 20312
rect 12584 20272 12590 20284
rect 12897 20281 12909 20284
rect 12943 20312 12955 20315
rect 13817 20315 13875 20321
rect 13817 20312 13829 20315
rect 12943 20284 13829 20312
rect 12943 20281 12955 20284
rect 12897 20275 12955 20281
rect 13817 20281 13829 20284
rect 13863 20281 13875 20315
rect 13817 20275 13875 20281
rect 14826 20272 14832 20324
rect 14884 20321 14890 20324
rect 14884 20315 14948 20321
rect 14884 20281 14902 20315
rect 14936 20281 14948 20315
rect 14884 20275 14948 20281
rect 14884 20272 14890 20275
rect 17034 20272 17040 20324
rect 17092 20312 17098 20324
rect 17497 20315 17555 20321
rect 17497 20312 17509 20315
rect 17092 20284 17509 20312
rect 17092 20272 17098 20284
rect 17497 20281 17509 20284
rect 17543 20312 17555 20315
rect 18316 20315 18374 20321
rect 18316 20312 18328 20315
rect 17543 20284 18328 20312
rect 17543 20281 17555 20284
rect 17497 20275 17555 20281
rect 18316 20281 18328 20284
rect 18362 20312 18374 20315
rect 18690 20312 18696 20324
rect 18362 20284 18696 20312
rect 18362 20281 18374 20284
rect 18316 20275 18374 20281
rect 18690 20272 18696 20284
rect 18748 20272 18754 20324
rect 24581 20315 24639 20321
rect 24581 20312 24593 20315
rect 23952 20284 24593 20312
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 1946 20244 1952 20256
rect 1907 20216 1952 20244
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 11333 20247 11391 20253
rect 11333 20213 11345 20247
rect 11379 20244 11391 20247
rect 11790 20244 11796 20256
rect 11379 20216 11796 20244
rect 11379 20213 11391 20216
rect 11333 20207 11391 20213
rect 11790 20204 11796 20216
rect 11848 20204 11854 20256
rect 12253 20247 12311 20253
rect 12253 20213 12265 20247
rect 12299 20244 12311 20247
rect 12805 20247 12863 20253
rect 12805 20244 12817 20247
rect 12299 20216 12817 20244
rect 12299 20213 12311 20216
rect 12253 20207 12311 20213
rect 12805 20213 12817 20216
rect 12851 20244 12863 20247
rect 13170 20244 13176 20256
rect 12851 20216 13176 20244
rect 12851 20213 12863 20216
rect 12805 20207 12863 20213
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 14182 20204 14188 20256
rect 14240 20244 14246 20256
rect 14461 20247 14519 20253
rect 14461 20244 14473 20247
rect 14240 20216 14473 20244
rect 14240 20204 14246 20216
rect 14461 20213 14473 20216
rect 14507 20244 14519 20247
rect 15378 20244 15384 20256
rect 14507 20216 15384 20244
rect 14507 20213 14519 20216
rect 14461 20207 14519 20213
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 20530 20244 20536 20256
rect 20491 20216 20536 20244
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 20901 20247 20959 20253
rect 20901 20244 20913 20247
rect 20680 20216 20913 20244
rect 20680 20204 20686 20216
rect 20901 20213 20913 20216
rect 20947 20244 20959 20247
rect 21358 20244 21364 20256
rect 20947 20216 21364 20244
rect 20947 20213 20959 20216
rect 20901 20207 20959 20213
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 23474 20204 23480 20256
rect 23532 20244 23538 20256
rect 23952 20253 23980 20284
rect 24581 20281 24593 20284
rect 24627 20312 24639 20315
rect 24854 20312 24860 20324
rect 24627 20284 24860 20312
rect 24627 20281 24639 20284
rect 24581 20275 24639 20281
rect 24854 20272 24860 20284
rect 24912 20272 24918 20324
rect 23937 20247 23995 20253
rect 23937 20244 23949 20247
rect 23532 20216 23949 20244
rect 23532 20204 23538 20216
rect 23937 20213 23949 20216
rect 23983 20213 23995 20247
rect 24118 20244 24124 20256
rect 24079 20216 24124 20244
rect 23937 20207 23995 20213
rect 24118 20204 24124 20216
rect 24176 20204 24182 20256
rect 24946 20204 24952 20256
rect 25004 20244 25010 20256
rect 25133 20247 25191 20253
rect 25133 20244 25145 20247
rect 25004 20216 25145 20244
rect 25004 20204 25010 20216
rect 25133 20213 25145 20216
rect 25179 20213 25191 20247
rect 25133 20207 25191 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 12158 20000 12164 20052
rect 12216 20040 12222 20052
rect 13909 20043 13967 20049
rect 13909 20040 13921 20043
rect 12216 20012 13921 20040
rect 12216 20000 12222 20012
rect 13909 20009 13921 20012
rect 13955 20009 13967 20043
rect 17678 20040 17684 20052
rect 17639 20012 17684 20040
rect 13909 20003 13967 20009
rect 17678 20000 17684 20012
rect 17736 20000 17742 20052
rect 18414 20040 18420 20052
rect 18375 20012 18420 20040
rect 18414 20000 18420 20012
rect 18472 20000 18478 20052
rect 18601 20043 18659 20049
rect 18601 20009 18613 20043
rect 18647 20040 18659 20043
rect 19150 20040 19156 20052
rect 18647 20012 19156 20040
rect 18647 20009 18659 20012
rect 18601 20003 18659 20009
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22281 20043 22339 20049
rect 22281 20040 22293 20043
rect 22152 20012 22293 20040
rect 22152 20000 22158 20012
rect 22281 20009 22293 20012
rect 22327 20009 22339 20043
rect 22281 20003 22339 20009
rect 23845 20043 23903 20049
rect 23845 20009 23857 20043
rect 23891 20040 23903 20043
rect 24118 20040 24124 20052
rect 23891 20012 24124 20040
rect 23891 20009 23903 20012
rect 23845 20003 23903 20009
rect 24118 20000 24124 20012
rect 24176 20000 24182 20052
rect 12796 19975 12854 19981
rect 12796 19941 12808 19975
rect 12842 19972 12854 19975
rect 12894 19972 12900 19984
rect 12842 19944 12900 19972
rect 12842 19941 12854 19944
rect 12796 19935 12854 19941
rect 12894 19932 12900 19944
rect 12952 19932 12958 19984
rect 15648 19975 15706 19981
rect 15648 19941 15660 19975
rect 15694 19972 15706 19975
rect 15838 19972 15844 19984
rect 15694 19944 15844 19972
rect 15694 19941 15706 19944
rect 15648 19935 15706 19941
rect 15838 19932 15844 19944
rect 15896 19932 15902 19984
rect 19058 19972 19064 19984
rect 18971 19944 19064 19972
rect 19058 19932 19064 19944
rect 19116 19972 19122 19984
rect 20530 19972 20536 19984
rect 19116 19944 20536 19972
rect 19116 19932 19122 19944
rect 20530 19932 20536 19944
rect 20588 19932 20594 19984
rect 21082 19932 21088 19984
rect 21140 19981 21146 19984
rect 21140 19975 21204 19981
rect 21140 19941 21158 19975
rect 21192 19941 21204 19975
rect 21140 19935 21204 19941
rect 24204 19975 24262 19981
rect 24204 19941 24216 19975
rect 24250 19972 24262 19975
rect 25038 19972 25044 19984
rect 24250 19944 25044 19972
rect 24250 19941 24262 19944
rect 24204 19935 24262 19941
rect 21140 19932 21146 19935
rect 25038 19932 25044 19944
rect 25096 19932 25102 19984
rect 10042 19904 10048 19916
rect 10003 19876 10048 19904
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 10134 19864 10140 19916
rect 10192 19904 10198 19916
rect 10301 19907 10359 19913
rect 10301 19904 10313 19907
rect 10192 19876 10313 19904
rect 10192 19864 10198 19876
rect 10301 19873 10313 19876
rect 10347 19904 10359 19907
rect 12158 19904 12164 19916
rect 10347 19876 12164 19904
rect 10347 19873 10359 19876
rect 10301 19867 10359 19873
rect 12158 19864 12164 19876
rect 12216 19864 12222 19916
rect 12529 19907 12587 19913
rect 12529 19873 12541 19907
rect 12575 19904 12587 19907
rect 13354 19904 13360 19916
rect 12575 19876 13360 19904
rect 12575 19873 12587 19876
rect 12529 19867 12587 19873
rect 13354 19864 13360 19876
rect 13412 19904 13418 19916
rect 14182 19904 14188 19916
rect 13412 19876 14188 19904
rect 13412 19864 13418 19876
rect 14182 19864 14188 19876
rect 14240 19904 14246 19916
rect 14642 19904 14648 19916
rect 14240 19876 14648 19904
rect 14240 19864 14246 19876
rect 14642 19864 14648 19876
rect 14700 19904 14706 19916
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14700 19876 14749 19904
rect 14700 19864 14706 19876
rect 14737 19873 14749 19876
rect 14783 19904 14795 19907
rect 15381 19907 15439 19913
rect 15381 19904 15393 19907
rect 14783 19876 15393 19904
rect 14783 19873 14795 19876
rect 14737 19867 14795 19873
rect 15381 19873 15393 19876
rect 15427 19904 15439 19907
rect 16206 19904 16212 19916
rect 15427 19876 16212 19904
rect 15427 19873 15439 19876
rect 15381 19867 15439 19873
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 18966 19904 18972 19916
rect 18927 19876 18972 19904
rect 18966 19864 18972 19876
rect 19024 19864 19030 19916
rect 20898 19904 20904 19916
rect 20859 19876 20904 19904
rect 20898 19864 20904 19876
rect 20956 19864 20962 19916
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19836 17463 19839
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 17451 19808 19257 19836
rect 17451 19805 17463 19808
rect 17405 19799 17463 19805
rect 19245 19805 19257 19808
rect 19291 19836 19303 19839
rect 19518 19836 19524 19848
rect 19291 19808 19524 19836
rect 19291 19805 19303 19808
rect 19245 19799 19303 19805
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 23842 19796 23848 19848
rect 23900 19836 23906 19848
rect 23937 19839 23995 19845
rect 23937 19836 23949 19839
rect 23900 19808 23949 19836
rect 23900 19796 23906 19808
rect 23937 19805 23949 19808
rect 23983 19805 23995 19839
rect 23937 19799 23995 19805
rect 19797 19771 19855 19777
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 20254 19768 20260 19780
rect 19843 19740 20260 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 20254 19728 20260 19740
rect 20312 19728 20318 19780
rect 1394 19660 1400 19712
rect 1452 19700 1458 19712
rect 1581 19703 1639 19709
rect 1581 19700 1593 19703
rect 1452 19672 1593 19700
rect 1452 19660 1458 19672
rect 1581 19669 1593 19672
rect 1627 19669 1639 19703
rect 11422 19700 11428 19712
rect 11383 19672 11428 19700
rect 1581 19663 1639 19669
rect 11422 19660 11428 19672
rect 11480 19660 11486 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 12526 19700 12532 19712
rect 11848 19672 12532 19700
rect 11848 19660 11854 19672
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 16758 19700 16764 19712
rect 16719 19672 16764 19700
rect 16758 19660 16764 19672
rect 16816 19660 16822 19712
rect 18138 19700 18144 19712
rect 18099 19672 18144 19700
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 20162 19700 20168 19712
rect 20123 19672 20168 19700
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 20622 19700 20628 19712
rect 20583 19672 20628 19700
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 22002 19660 22008 19712
rect 22060 19700 22066 19712
rect 22833 19703 22891 19709
rect 22833 19700 22845 19703
rect 22060 19672 22845 19700
rect 22060 19660 22066 19672
rect 22833 19669 22845 19672
rect 22879 19669 22891 19703
rect 25314 19700 25320 19712
rect 25275 19672 25320 19700
rect 22833 19663 22891 19669
rect 25314 19660 25320 19672
rect 25372 19660 25378 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 9769 19499 9827 19505
rect 9769 19465 9781 19499
rect 9815 19496 9827 19499
rect 10042 19496 10048 19508
rect 9815 19468 10048 19496
rect 9815 19465 9827 19468
rect 9769 19459 9827 19465
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 11790 19496 11796 19508
rect 11751 19468 11796 19496
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 15838 19456 15844 19508
rect 15896 19496 15902 19508
rect 16485 19499 16543 19505
rect 16485 19496 16497 19499
rect 15896 19468 16497 19496
rect 15896 19456 15902 19468
rect 16485 19465 16497 19468
rect 16531 19465 16543 19499
rect 16485 19459 16543 19465
rect 19153 19499 19211 19505
rect 19153 19465 19165 19499
rect 19199 19496 19211 19499
rect 19518 19496 19524 19508
rect 19199 19468 19524 19496
rect 19199 19465 19211 19468
rect 19153 19459 19211 19465
rect 19518 19456 19524 19468
rect 19576 19456 19582 19508
rect 20898 19496 20904 19508
rect 20859 19468 20904 19496
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 22094 19456 22100 19508
rect 22152 19496 22158 19508
rect 22281 19499 22339 19505
rect 22281 19496 22293 19499
rect 22152 19468 22293 19496
rect 22152 19456 22158 19468
rect 22281 19465 22293 19468
rect 22327 19465 22339 19499
rect 25038 19496 25044 19508
rect 24999 19468 25044 19496
rect 22281 19459 22339 19465
rect 25038 19456 25044 19468
rect 25096 19456 25102 19508
rect 18049 19431 18107 19437
rect 18049 19397 18061 19431
rect 18095 19428 18107 19431
rect 18966 19428 18972 19440
rect 18095 19400 18972 19428
rect 18095 19397 18107 19400
rect 18049 19391 18107 19397
rect 18966 19388 18972 19400
rect 19024 19388 19030 19440
rect 19705 19431 19763 19437
rect 19705 19397 19717 19431
rect 19751 19397 19763 19431
rect 21174 19428 21180 19440
rect 19705 19391 19763 19397
rect 20916 19400 21180 19428
rect 10134 19360 10140 19372
rect 9600 19332 10140 19360
rect 9401 19295 9459 19301
rect 9401 19261 9413 19295
rect 9447 19292 9459 19295
rect 9600 19292 9628 19332
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 10870 19360 10876 19372
rect 10831 19332 10876 19360
rect 10870 19320 10876 19332
rect 10928 19360 10934 19372
rect 11241 19363 11299 19369
rect 11241 19360 11253 19363
rect 10928 19332 11253 19360
rect 10928 19320 10934 19332
rect 11241 19329 11253 19332
rect 11287 19360 11299 19363
rect 11422 19360 11428 19372
rect 11287 19332 11428 19360
rect 11287 19329 11299 19332
rect 11241 19323 11299 19329
rect 11422 19320 11428 19332
rect 11480 19320 11486 19372
rect 12434 19320 12440 19372
rect 12492 19320 12498 19372
rect 12894 19320 12900 19372
rect 12952 19360 12958 19372
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 12952 19332 13001 19360
rect 12952 19320 12958 19332
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 14093 19363 14151 19369
rect 14093 19329 14105 19363
rect 14139 19360 14151 19363
rect 14182 19360 14188 19372
rect 14139 19332 14188 19360
rect 14139 19329 14151 19332
rect 14093 19323 14151 19329
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 17497 19363 17555 19369
rect 17497 19329 17509 19363
rect 17543 19360 17555 19363
rect 18690 19360 18696 19372
rect 17543 19332 18696 19360
rect 17543 19329 17555 19332
rect 17497 19323 17555 19329
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 9447 19264 9628 19292
rect 9447 19261 9459 19264
rect 9401 19255 9459 19261
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 10045 19295 10103 19301
rect 10045 19292 10057 19295
rect 9732 19264 10057 19292
rect 9732 19252 9738 19264
rect 10045 19261 10057 19264
rect 10091 19292 10103 19295
rect 10597 19295 10655 19301
rect 10597 19292 10609 19295
rect 10091 19264 10609 19292
rect 10091 19261 10103 19264
rect 10045 19255 10103 19261
rect 10597 19261 10609 19264
rect 10643 19261 10655 19295
rect 12452 19292 12480 19320
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12452 19264 12817 19292
rect 10597 19255 10655 19261
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 16945 19295 17003 19301
rect 16945 19261 16957 19295
rect 16991 19292 17003 19295
rect 18138 19292 18144 19304
rect 16991 19264 18144 19292
rect 16991 19261 17003 19264
rect 16945 19255 17003 19261
rect 18138 19252 18144 19264
rect 18196 19292 18202 19304
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 18196 19264 18429 19292
rect 18196 19252 18202 19264
rect 18417 19261 18429 19264
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 19720 19292 19748 19391
rect 20916 19372 20944 19400
rect 21174 19388 21180 19400
rect 21232 19388 21238 19440
rect 20254 19360 20260 19372
rect 20215 19332 20260 19360
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 20898 19320 20904 19372
rect 20956 19320 20962 19372
rect 21913 19363 21971 19369
rect 21913 19329 21925 19363
rect 21959 19360 21971 19363
rect 22112 19360 22140 19456
rect 24578 19360 24584 19372
rect 21959 19332 22140 19360
rect 23584 19332 24584 19360
rect 21959 19329 21971 19332
rect 21913 19323 21971 19329
rect 19300 19264 19748 19292
rect 19300 19252 19306 19264
rect 21174 19252 21180 19304
rect 21232 19292 21238 19304
rect 21637 19295 21695 19301
rect 21637 19292 21649 19295
rect 21232 19264 21649 19292
rect 21232 19252 21238 19264
rect 21637 19261 21649 19264
rect 21683 19292 21695 19295
rect 22002 19292 22008 19304
rect 21683 19264 22008 19292
rect 21683 19261 21695 19264
rect 21637 19255 21695 19261
rect 22002 19252 22008 19264
rect 22060 19252 22066 19304
rect 23109 19295 23167 19301
rect 23109 19261 23121 19295
rect 23155 19292 23167 19295
rect 23584 19292 23612 19332
rect 24578 19320 24584 19332
rect 24636 19360 24642 19372
rect 25314 19360 25320 19372
rect 24636 19332 25320 19360
rect 24636 19320 24642 19332
rect 25314 19320 25320 19332
rect 25372 19320 25378 19372
rect 23155 19264 23612 19292
rect 23155 19261 23167 19264
rect 23109 19255 23167 19261
rect 23934 19252 23940 19304
rect 23992 19292 23998 19304
rect 23992 19264 24072 19292
rect 23992 19252 23998 19264
rect 12253 19227 12311 19233
rect 12253 19193 12265 19227
rect 12299 19224 12311 19227
rect 13725 19227 13783 19233
rect 12299 19196 12940 19224
rect 12299 19193 12311 19196
rect 12253 19187 12311 19193
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10229 19159 10287 19165
rect 10229 19156 10241 19159
rect 10192 19128 10241 19156
rect 10192 19116 10198 19128
rect 10229 19125 10241 19128
rect 10275 19125 10287 19159
rect 10229 19119 10287 19125
rect 10689 19159 10747 19165
rect 10689 19125 10701 19159
rect 10735 19156 10747 19159
rect 10778 19156 10784 19168
rect 10735 19128 10784 19156
rect 10735 19125 10747 19128
rect 10689 19119 10747 19125
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 12434 19156 12440 19168
rect 12395 19128 12440 19156
rect 12434 19116 12440 19128
rect 12492 19116 12498 19168
rect 12912 19165 12940 19196
rect 13725 19193 13737 19227
rect 13771 19224 13783 19227
rect 14430 19227 14488 19233
rect 14430 19224 14442 19227
rect 13771 19196 14442 19224
rect 13771 19193 13783 19196
rect 13725 19187 13783 19193
rect 14430 19193 14442 19196
rect 14476 19224 14488 19227
rect 15746 19224 15752 19236
rect 14476 19196 15752 19224
rect 14476 19193 14488 19196
rect 14430 19187 14488 19193
rect 15746 19184 15752 19196
rect 15804 19184 15810 19236
rect 17126 19184 17132 19236
rect 17184 19224 17190 19236
rect 20073 19227 20131 19233
rect 20073 19224 20085 19227
rect 17184 19196 17908 19224
rect 17184 19184 17190 19196
rect 12897 19159 12955 19165
rect 12897 19125 12909 19159
rect 12943 19156 12955 19159
rect 13170 19156 13176 19168
rect 12943 19128 13176 19156
rect 12943 19125 12955 19128
rect 12897 19119 12955 19125
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 14182 19116 14188 19168
rect 14240 19156 14246 19168
rect 14826 19156 14832 19168
rect 14240 19128 14832 19156
rect 14240 19116 14246 19128
rect 14826 19116 14832 19128
rect 14884 19156 14890 19168
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 14884 19128 15577 19156
rect 14884 19116 14890 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 16206 19156 16212 19168
rect 16119 19128 16212 19156
rect 15565 19119 15623 19125
rect 16206 19116 16212 19128
rect 16264 19156 16270 19168
rect 16942 19156 16948 19168
rect 16264 19128 16948 19156
rect 16264 19116 16270 19128
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 17880 19165 17908 19196
rect 19536 19196 20085 19224
rect 19536 19168 19564 19196
rect 20073 19193 20085 19196
rect 20119 19193 20131 19227
rect 20073 19187 20131 19193
rect 23477 19227 23535 19233
rect 23477 19193 23489 19227
rect 23523 19224 23535 19227
rect 23842 19224 23848 19236
rect 23523 19196 23848 19224
rect 23523 19193 23535 19196
rect 23477 19187 23535 19193
rect 23842 19184 23848 19196
rect 23900 19184 23906 19236
rect 17865 19159 17923 19165
rect 17865 19125 17877 19159
rect 17911 19156 17923 19159
rect 18506 19156 18512 19168
rect 17911 19128 18512 19156
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 19518 19156 19524 19168
rect 19479 19128 19524 19156
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 20162 19156 20168 19168
rect 20075 19128 20168 19156
rect 20162 19116 20168 19128
rect 20220 19156 20226 19168
rect 20622 19156 20628 19168
rect 20220 19128 20628 19156
rect 20220 19116 20226 19128
rect 20622 19116 20628 19128
rect 20680 19116 20686 19168
rect 21266 19156 21272 19168
rect 21227 19128 21272 19156
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 21726 19156 21732 19168
rect 21687 19128 21732 19156
rect 21726 19116 21732 19128
rect 21784 19116 21790 19168
rect 22278 19116 22284 19168
rect 22336 19156 22342 19168
rect 22649 19159 22707 19165
rect 22649 19156 22661 19159
rect 22336 19128 22661 19156
rect 22336 19116 22342 19128
rect 22649 19125 22661 19128
rect 22695 19125 22707 19159
rect 23934 19156 23940 19168
rect 23895 19128 23940 19156
rect 22649 19119 22707 19125
rect 23934 19116 23940 19128
rect 23992 19116 23998 19168
rect 24044 19156 24072 19264
rect 24118 19252 24124 19304
rect 24176 19292 24182 19304
rect 24305 19295 24363 19301
rect 24305 19292 24317 19295
rect 24176 19264 24317 19292
rect 24176 19252 24182 19264
rect 24305 19261 24317 19264
rect 24351 19261 24363 19295
rect 25498 19292 25504 19304
rect 25459 19264 25504 19292
rect 24305 19255 24363 19261
rect 25498 19252 25504 19264
rect 25556 19292 25562 19304
rect 26053 19295 26111 19301
rect 26053 19292 26065 19295
rect 25556 19264 26065 19292
rect 25556 19252 25562 19264
rect 26053 19261 26065 19264
rect 26099 19261 26111 19295
rect 26053 19255 26111 19261
rect 24210 19184 24216 19236
rect 24268 19224 24274 19236
rect 24397 19227 24455 19233
rect 24397 19224 24409 19227
rect 24268 19196 24409 19224
rect 24268 19184 24274 19196
rect 24397 19193 24409 19196
rect 24443 19224 24455 19227
rect 25317 19227 25375 19233
rect 25317 19224 25329 19227
rect 24443 19196 25329 19224
rect 24443 19193 24455 19196
rect 24397 19187 24455 19193
rect 25317 19193 25329 19196
rect 25363 19193 25375 19227
rect 25317 19187 25375 19193
rect 24118 19156 24124 19168
rect 24044 19128 24124 19156
rect 24118 19116 24124 19128
rect 24176 19116 24182 19168
rect 25682 19156 25688 19168
rect 25643 19128 25688 19156
rect 25682 19116 25688 19128
rect 25740 19116 25746 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 12894 18952 12900 18964
rect 12855 18924 12900 18952
rect 12894 18912 12900 18924
rect 12952 18952 12958 18964
rect 13265 18955 13323 18961
rect 13265 18952 13277 18955
rect 12952 18924 13277 18952
rect 12952 18912 12958 18924
rect 13265 18921 13277 18924
rect 13311 18921 13323 18955
rect 13265 18915 13323 18921
rect 13633 18955 13691 18961
rect 13633 18921 13645 18955
rect 13679 18952 13691 18955
rect 13722 18952 13728 18964
rect 13679 18924 13728 18952
rect 13679 18921 13691 18924
rect 13633 18915 13691 18921
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 14001 18955 14059 18961
rect 14001 18952 14013 18955
rect 13964 18924 14013 18952
rect 13964 18912 13970 18924
rect 14001 18921 14013 18924
rect 14047 18921 14059 18955
rect 14001 18915 14059 18921
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 15105 18955 15163 18961
rect 14148 18924 14193 18952
rect 14148 18912 14154 18924
rect 15105 18921 15117 18955
rect 15151 18952 15163 18955
rect 15286 18952 15292 18964
rect 15151 18924 15292 18952
rect 15151 18921 15163 18924
rect 15105 18915 15163 18921
rect 15286 18912 15292 18924
rect 15344 18952 15350 18964
rect 15749 18955 15807 18961
rect 15749 18952 15761 18955
rect 15344 18924 15761 18952
rect 15344 18912 15350 18924
rect 15749 18921 15761 18924
rect 15795 18921 15807 18955
rect 15749 18915 15807 18921
rect 18966 18912 18972 18964
rect 19024 18952 19030 18964
rect 19337 18955 19395 18961
rect 19337 18952 19349 18955
rect 19024 18924 19349 18952
rect 19024 18912 19030 18924
rect 19337 18921 19349 18924
rect 19383 18921 19395 18955
rect 21174 18952 21180 18964
rect 21135 18924 21180 18952
rect 19337 18915 19395 18921
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 21542 18952 21548 18964
rect 21503 18924 21548 18952
rect 21542 18912 21548 18924
rect 21600 18912 21606 18964
rect 21726 18912 21732 18964
rect 21784 18952 21790 18964
rect 22557 18955 22615 18961
rect 22557 18952 22569 18955
rect 21784 18924 22569 18952
rect 21784 18912 21790 18924
rect 22557 18921 22569 18924
rect 22603 18921 22615 18955
rect 23658 18952 23664 18964
rect 23619 18924 23664 18952
rect 22557 18915 22615 18921
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 14734 18844 14740 18896
rect 14792 18884 14798 18896
rect 15841 18887 15899 18893
rect 15841 18884 15853 18887
rect 14792 18856 15853 18884
rect 14792 18844 14798 18856
rect 15841 18853 15853 18856
rect 15887 18884 15899 18887
rect 16666 18884 16672 18896
rect 15887 18856 16672 18884
rect 15887 18853 15899 18856
rect 15841 18847 15899 18853
rect 16666 18844 16672 18856
rect 16724 18844 16730 18896
rect 19058 18884 19064 18896
rect 19019 18856 19064 18884
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 24112 18887 24170 18893
rect 24112 18853 24124 18887
rect 24158 18884 24170 18887
rect 24210 18884 24216 18896
rect 24158 18856 24216 18884
rect 24158 18853 24170 18856
rect 24112 18847 24170 18853
rect 24210 18844 24216 18856
rect 24268 18884 24274 18896
rect 24578 18884 24584 18896
rect 24268 18856 24584 18884
rect 24268 18844 24274 18856
rect 24578 18844 24584 18856
rect 24636 18844 24642 18896
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 10870 18825 10876 18828
rect 10853 18819 10876 18825
rect 10853 18816 10865 18819
rect 10376 18788 10865 18816
rect 10376 18776 10382 18788
rect 10853 18785 10865 18788
rect 10928 18816 10934 18828
rect 17304 18819 17362 18825
rect 10928 18788 11001 18816
rect 10853 18779 10876 18785
rect 10870 18776 10876 18779
rect 10928 18776 10934 18788
rect 17304 18785 17316 18819
rect 17350 18816 17362 18819
rect 17678 18816 17684 18828
rect 17350 18788 17684 18816
rect 17350 18785 17362 18788
rect 17304 18779 17362 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 19794 18816 19800 18828
rect 19755 18788 19800 18816
rect 19794 18776 19800 18788
rect 19852 18776 19858 18828
rect 22278 18816 22284 18828
rect 22239 18788 22284 18816
rect 22278 18776 22284 18788
rect 22336 18776 22342 18828
rect 10042 18708 10048 18760
rect 10100 18748 10106 18760
rect 10594 18748 10600 18760
rect 10100 18720 10600 18748
rect 10100 18708 10106 18720
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 14182 18708 14188 18760
rect 14240 18748 14246 18760
rect 16022 18748 16028 18760
rect 14240 18720 14285 18748
rect 15983 18720 16028 18748
rect 14240 18708 14246 18720
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17037 18751 17095 18757
rect 17037 18748 17049 18751
rect 17000 18720 17049 18748
rect 17000 18708 17006 18720
rect 17037 18717 17049 18720
rect 17083 18717 17095 18751
rect 17037 18711 17095 18717
rect 21174 18708 21180 18760
rect 21232 18748 21238 18760
rect 21634 18748 21640 18760
rect 21232 18720 21640 18748
rect 21232 18708 21238 18720
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 21729 18751 21787 18757
rect 21729 18717 21741 18751
rect 21775 18748 21787 18751
rect 22296 18748 22324 18776
rect 21775 18720 22324 18748
rect 22833 18751 22891 18757
rect 21775 18717 21787 18720
rect 21729 18711 21787 18717
rect 22833 18717 22845 18751
rect 22879 18748 22891 18751
rect 23382 18748 23388 18760
rect 22879 18720 23388 18748
rect 22879 18717 22891 18720
rect 22833 18711 22891 18717
rect 18417 18683 18475 18689
rect 18417 18649 18429 18683
rect 18463 18680 18475 18683
rect 20717 18683 20775 18689
rect 20717 18680 20729 18683
rect 18463 18652 20729 18680
rect 18463 18649 18475 18652
rect 18417 18643 18475 18649
rect 20717 18649 20729 18652
rect 20763 18680 20775 18683
rect 21082 18680 21088 18692
rect 20763 18652 21088 18680
rect 20763 18649 20775 18652
rect 20717 18643 20775 18649
rect 21082 18640 21088 18652
rect 21140 18680 21146 18692
rect 21744 18680 21772 18711
rect 23382 18708 23388 18720
rect 23440 18708 23446 18760
rect 23842 18748 23848 18760
rect 23803 18720 23848 18748
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 21140 18652 21772 18680
rect 21140 18640 21146 18652
rect 22922 18640 22928 18692
rect 22980 18680 22986 18692
rect 23474 18680 23480 18692
rect 22980 18652 23480 18680
rect 22980 18640 22986 18652
rect 23474 18640 23480 18652
rect 23532 18640 23538 18692
rect 10321 18615 10379 18621
rect 10321 18581 10333 18615
rect 10367 18612 10379 18615
rect 10778 18612 10784 18624
rect 10367 18584 10784 18612
rect 10367 18581 10379 18584
rect 10321 18575 10379 18581
rect 10778 18572 10784 18584
rect 10836 18572 10842 18624
rect 11974 18612 11980 18624
rect 11935 18584 11980 18612
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12621 18615 12679 18621
rect 12621 18581 12633 18615
rect 12667 18612 12679 18615
rect 13998 18612 14004 18624
rect 12667 18584 14004 18612
rect 12667 18581 12679 18584
rect 12621 18575 12679 18581
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 14642 18612 14648 18624
rect 14603 18584 14648 18612
rect 14642 18572 14648 18584
rect 14700 18572 14706 18624
rect 15378 18612 15384 18624
rect 15339 18584 15384 18612
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 16853 18615 16911 18621
rect 16853 18612 16865 18615
rect 16632 18584 16865 18612
rect 16632 18572 16638 18584
rect 16853 18581 16865 18584
rect 16899 18581 16911 18615
rect 19978 18612 19984 18624
rect 19939 18584 19984 18612
rect 16853 18575 16911 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 25222 18612 25228 18624
rect 25183 18584 25228 18612
rect 25222 18572 25228 18584
rect 25280 18572 25286 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 10318 18408 10324 18420
rect 10279 18380 10324 18408
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 10594 18408 10600 18420
rect 10555 18380 10600 18408
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 13906 18368 13912 18420
rect 13964 18408 13970 18420
rect 14185 18411 14243 18417
rect 14185 18408 14197 18411
rect 13964 18380 14197 18408
rect 13964 18368 13970 18380
rect 14185 18377 14197 18380
rect 14231 18377 14243 18411
rect 15746 18408 15752 18420
rect 15707 18380 15752 18408
rect 14185 18371 14243 18377
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 16022 18368 16028 18420
rect 16080 18408 16086 18420
rect 16393 18411 16451 18417
rect 16393 18408 16405 18411
rect 16080 18380 16405 18408
rect 16080 18368 16086 18380
rect 16393 18377 16405 18380
rect 16439 18408 16451 18411
rect 16758 18408 16764 18420
rect 16439 18380 16764 18408
rect 16439 18377 16451 18380
rect 16393 18371 16451 18377
rect 16758 18368 16764 18380
rect 16816 18408 16822 18420
rect 17678 18408 17684 18420
rect 16816 18380 17684 18408
rect 16816 18368 16822 18380
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 18598 18408 18604 18420
rect 18559 18380 18604 18408
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 20438 18408 20444 18420
rect 20399 18380 20444 18408
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 21545 18411 21603 18417
rect 21545 18377 21557 18411
rect 21591 18408 21603 18411
rect 21726 18408 21732 18420
rect 21591 18380 21732 18408
rect 21591 18377 21603 18380
rect 21545 18371 21603 18377
rect 21726 18368 21732 18380
rect 21784 18368 21790 18420
rect 23198 18368 23204 18420
rect 23256 18408 23262 18420
rect 23385 18411 23443 18417
rect 23385 18408 23397 18411
rect 23256 18380 23397 18408
rect 23256 18368 23262 18380
rect 23385 18377 23397 18380
rect 23431 18377 23443 18411
rect 23385 18371 23443 18377
rect 10781 18343 10839 18349
rect 10781 18309 10793 18343
rect 10827 18340 10839 18343
rect 11146 18340 11152 18352
rect 10827 18312 11152 18340
rect 10827 18309 10839 18312
rect 10781 18303 10839 18309
rect 11146 18300 11152 18312
rect 11204 18300 11210 18352
rect 11793 18343 11851 18349
rect 11793 18340 11805 18343
rect 11256 18312 11805 18340
rect 10134 18232 10140 18284
rect 10192 18272 10198 18284
rect 11256 18281 11284 18312
rect 11793 18309 11805 18312
rect 11839 18309 11851 18343
rect 11793 18303 11851 18309
rect 13817 18343 13875 18349
rect 13817 18309 13829 18343
rect 13863 18340 13875 18343
rect 14090 18340 14096 18352
rect 13863 18312 14096 18340
rect 13863 18309 13875 18312
rect 13817 18303 13875 18309
rect 14090 18300 14096 18312
rect 14148 18300 14154 18352
rect 16666 18340 16672 18352
rect 16627 18312 16672 18340
rect 16666 18300 16672 18312
rect 16724 18300 16730 18352
rect 11241 18275 11299 18281
rect 11241 18272 11253 18275
rect 10192 18244 11253 18272
rect 10192 18232 10198 18244
rect 11241 18241 11253 18244
rect 11287 18241 11299 18275
rect 11422 18272 11428 18284
rect 11335 18244 11428 18272
rect 11241 18235 11299 18241
rect 11422 18232 11428 18244
rect 11480 18272 11486 18284
rect 11974 18272 11980 18284
rect 11480 18244 11980 18272
rect 11480 18232 11486 18244
rect 11974 18232 11980 18244
rect 12032 18232 12038 18284
rect 13265 18275 13323 18281
rect 13265 18241 13277 18275
rect 13311 18272 13323 18275
rect 14182 18272 14188 18284
rect 13311 18244 14188 18272
rect 13311 18241 13323 18244
rect 13265 18235 13323 18241
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18272 22063 18275
rect 22094 18272 22100 18284
rect 22051 18244 22100 18272
rect 22051 18241 22063 18244
rect 22005 18235 22063 18241
rect 22094 18232 22100 18244
rect 22152 18232 22158 18284
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18272 22247 18275
rect 22278 18272 22284 18284
rect 22235 18244 22284 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 22278 18232 22284 18244
rect 22336 18232 22342 18284
rect 23400 18272 23428 18371
rect 23842 18368 23848 18420
rect 23900 18408 23906 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 23900 18380 24685 18408
rect 23900 18368 23906 18380
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 24673 18371 24731 18377
rect 25133 18411 25191 18417
rect 25133 18377 25145 18411
rect 25179 18408 25191 18411
rect 25222 18408 25228 18420
rect 25179 18380 25228 18408
rect 25179 18377 25191 18380
rect 25133 18371 25191 18377
rect 24121 18275 24179 18281
rect 24121 18272 24133 18275
rect 23400 18244 24133 18272
rect 24121 18241 24133 18244
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18272 24363 18275
rect 24762 18272 24768 18284
rect 24351 18244 24768 18272
rect 24351 18241 24363 18244
rect 24305 18235 24363 18241
rect 24762 18232 24768 18244
rect 24820 18272 24826 18284
rect 25148 18272 25176 18371
rect 25222 18368 25228 18380
rect 25280 18368 25286 18420
rect 24820 18244 25176 18272
rect 24820 18232 24826 18244
rect 9953 18207 10011 18213
rect 9953 18173 9965 18207
rect 9999 18204 10011 18207
rect 11440 18204 11468 18232
rect 13354 18204 13360 18216
rect 9999 18176 11468 18204
rect 13315 18176 13360 18204
rect 9999 18173 10011 18176
rect 9953 18167 10011 18173
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 13998 18164 14004 18216
rect 14056 18204 14062 18216
rect 14642 18213 14648 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 14056 18176 14381 18204
rect 14056 18164 14062 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14636 18204 14648 18213
rect 14603 18176 14648 18204
rect 14369 18167 14427 18173
rect 14636 18167 14648 18176
rect 14384 18136 14412 18167
rect 14642 18164 14648 18167
rect 14700 18164 14706 18216
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 16853 18207 16911 18213
rect 16853 18204 16865 18207
rect 16632 18176 16865 18204
rect 16632 18164 16638 18176
rect 16853 18173 16865 18176
rect 16899 18173 16911 18207
rect 16853 18167 16911 18173
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 18598 18204 18604 18216
rect 18095 18176 18604 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 19061 18207 19119 18213
rect 19061 18173 19073 18207
rect 19107 18173 19119 18207
rect 19061 18167 19119 18173
rect 14734 18136 14740 18148
rect 14384 18108 14740 18136
rect 14734 18096 14740 18108
rect 14792 18096 14798 18148
rect 16942 18096 16948 18148
rect 17000 18136 17006 18148
rect 17313 18139 17371 18145
rect 17313 18136 17325 18139
rect 17000 18108 17325 18136
rect 17000 18096 17006 18108
rect 17313 18105 17325 18108
rect 17359 18136 17371 18139
rect 18877 18139 18935 18145
rect 18877 18136 18889 18139
rect 17359 18108 18889 18136
rect 17359 18105 17371 18108
rect 17313 18099 17371 18105
rect 18064 18080 18092 18108
rect 18877 18105 18889 18108
rect 18923 18136 18935 18139
rect 19076 18136 19104 18167
rect 21542 18164 21548 18216
rect 21600 18204 21606 18216
rect 22925 18207 22983 18213
rect 22925 18204 22937 18207
rect 21600 18176 22937 18204
rect 21600 18164 21606 18176
rect 22925 18173 22937 18176
rect 22971 18173 22983 18207
rect 22925 18167 22983 18173
rect 23658 18164 23664 18216
rect 23716 18204 23722 18216
rect 24029 18207 24087 18213
rect 24029 18204 24041 18207
rect 23716 18176 24041 18204
rect 23716 18164 23722 18176
rect 24029 18173 24041 18176
rect 24075 18173 24087 18207
rect 25222 18204 25228 18216
rect 25183 18176 25228 18204
rect 24029 18167 24087 18173
rect 25222 18164 25228 18176
rect 25280 18204 25286 18216
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25280 18176 25789 18204
rect 25280 18164 25286 18176
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 19334 18145 19340 18148
rect 19328 18136 19340 18145
rect 18923 18108 19104 18136
rect 19295 18108 19340 18136
rect 18923 18105 18935 18108
rect 18877 18099 18935 18105
rect 19328 18099 19340 18108
rect 19334 18096 19340 18099
rect 19392 18096 19398 18148
rect 21358 18096 21364 18148
rect 21416 18136 21422 18148
rect 21913 18139 21971 18145
rect 21913 18136 21925 18139
rect 21416 18108 21925 18136
rect 21416 18096 21422 18108
rect 21913 18105 21925 18108
rect 21959 18136 21971 18139
rect 22554 18136 22560 18148
rect 21959 18108 22560 18136
rect 21959 18105 21971 18108
rect 21913 18099 21971 18105
rect 22554 18096 22560 18108
rect 22612 18096 22618 18148
rect 23566 18096 23572 18148
rect 23624 18136 23630 18148
rect 23842 18136 23848 18148
rect 23624 18108 23848 18136
rect 23624 18096 23630 18108
rect 23842 18096 23848 18108
rect 23900 18096 23906 18148
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11149 18071 11207 18077
rect 11149 18068 11161 18071
rect 11112 18040 11161 18068
rect 11112 18028 11118 18040
rect 11149 18037 11161 18040
rect 11195 18037 11207 18071
rect 13538 18068 13544 18080
rect 13499 18040 13544 18068
rect 11149 18031 11207 18037
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 17037 18071 17095 18077
rect 17037 18037 17049 18071
rect 17083 18068 17095 18071
rect 17218 18068 17224 18080
rect 17083 18040 17224 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 17218 18028 17224 18040
rect 17276 18028 17282 18080
rect 18046 18028 18052 18080
rect 18104 18028 18110 18080
rect 18230 18068 18236 18080
rect 18191 18040 18236 18068
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 21266 18068 21272 18080
rect 21227 18040 21272 18068
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 23658 18068 23664 18080
rect 23619 18040 23664 18068
rect 23658 18028 23664 18040
rect 23716 18028 23722 18080
rect 25406 18068 25412 18080
rect 25367 18040 25412 18068
rect 25406 18028 25412 18040
rect 25464 18028 25470 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 13354 17864 13360 17876
rect 13315 17836 13360 17864
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 13633 17867 13691 17873
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 15749 17867 15807 17873
rect 15749 17864 15761 17867
rect 13679 17836 15761 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 15749 17833 15761 17836
rect 15795 17864 15807 17867
rect 16669 17867 16727 17873
rect 16669 17864 16681 17867
rect 15795 17836 16681 17864
rect 15795 17833 15807 17836
rect 15749 17827 15807 17833
rect 16669 17833 16681 17836
rect 16715 17833 16727 17867
rect 16669 17827 16727 17833
rect 19981 17867 20039 17873
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 20070 17864 20076 17876
rect 20027 17836 20076 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 20346 17864 20352 17876
rect 20307 17836 20352 17864
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 20901 17867 20959 17873
rect 20901 17864 20913 17867
rect 20772 17836 20913 17864
rect 20772 17824 20778 17836
rect 20901 17833 20913 17836
rect 20947 17833 20959 17867
rect 20901 17827 20959 17833
rect 20990 17824 20996 17876
rect 21048 17864 21054 17876
rect 21361 17867 21419 17873
rect 21361 17864 21373 17867
rect 21048 17836 21373 17864
rect 21048 17824 21054 17836
rect 21361 17833 21373 17836
rect 21407 17833 21419 17867
rect 21361 17827 21419 17833
rect 23109 17867 23167 17873
rect 23109 17833 23121 17867
rect 23155 17864 23167 17867
rect 23658 17864 23664 17876
rect 23155 17836 23664 17864
rect 23155 17833 23167 17836
rect 23109 17827 23167 17833
rect 23658 17824 23664 17836
rect 23716 17824 23722 17876
rect 24210 17864 24216 17876
rect 24171 17836 24216 17864
rect 24210 17824 24216 17836
rect 24268 17824 24274 17876
rect 11422 17805 11428 17808
rect 11416 17796 11428 17805
rect 11383 17768 11428 17796
rect 11416 17759 11428 17768
rect 11422 17756 11428 17759
rect 11480 17756 11486 17808
rect 13998 17796 14004 17808
rect 13959 17768 14004 17796
rect 13998 17756 14004 17768
rect 14056 17756 14062 17808
rect 14093 17799 14151 17805
rect 14093 17765 14105 17799
rect 14139 17796 14151 17799
rect 14274 17796 14280 17808
rect 14139 17768 14280 17796
rect 14139 17765 14151 17768
rect 14093 17759 14151 17765
rect 14274 17756 14280 17768
rect 14332 17756 14338 17808
rect 14734 17796 14740 17808
rect 14695 17768 14740 17796
rect 14734 17756 14740 17768
rect 14792 17756 14798 17808
rect 17212 17799 17270 17805
rect 17212 17765 17224 17799
rect 17258 17796 17270 17799
rect 17402 17796 17408 17808
rect 17258 17768 17408 17796
rect 17258 17765 17270 17768
rect 17212 17759 17270 17765
rect 17402 17756 17408 17768
rect 17460 17756 17466 17808
rect 23290 17756 23296 17808
rect 23348 17796 23354 17808
rect 23348 17768 24808 17796
rect 23348 17756 23354 17768
rect 14 17688 20 17740
rect 72 17728 78 17740
rect 9582 17728 9588 17740
rect 72 17700 9588 17728
rect 72 17688 78 17700
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 10686 17688 10692 17740
rect 10744 17728 10750 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10744 17700 11161 17728
rect 10744 17688 10750 17700
rect 11149 17697 11161 17700
rect 11195 17728 11207 17731
rect 11790 17728 11796 17740
rect 11195 17700 11796 17728
rect 11195 17697 11207 17700
rect 11149 17691 11207 17697
rect 11790 17688 11796 17700
rect 11848 17688 11854 17740
rect 14642 17688 14648 17740
rect 14700 17728 14706 17740
rect 15654 17728 15660 17740
rect 14700 17700 15424 17728
rect 15615 17700 15660 17728
rect 14700 17688 14706 17700
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 14826 17660 14832 17672
rect 14323 17632 14832 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 14826 17620 14832 17632
rect 14884 17660 14890 17672
rect 15013 17663 15071 17669
rect 15013 17660 15025 17663
rect 14884 17632 15025 17660
rect 14884 17620 14890 17632
rect 15013 17629 15025 17632
rect 15059 17629 15071 17663
rect 15396 17660 15424 17700
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 19794 17728 19800 17740
rect 19755 17700 19800 17728
rect 19794 17688 19800 17700
rect 19852 17688 19858 17740
rect 20714 17688 20720 17740
rect 20772 17728 20778 17740
rect 20898 17728 20904 17740
rect 20772 17700 20904 17728
rect 20772 17688 20778 17700
rect 20898 17688 20904 17700
rect 20956 17688 20962 17740
rect 21269 17731 21327 17737
rect 21269 17697 21281 17731
rect 21315 17728 21327 17731
rect 21358 17728 21364 17740
rect 21315 17700 21364 17728
rect 21315 17697 21327 17700
rect 21269 17691 21327 17697
rect 21358 17688 21364 17700
rect 21416 17688 21422 17740
rect 23566 17728 23572 17740
rect 23527 17700 23572 17728
rect 23566 17688 23572 17700
rect 23624 17688 23630 17740
rect 24780 17737 24808 17768
rect 24765 17731 24823 17737
rect 24765 17697 24777 17731
rect 24811 17728 24823 17731
rect 25590 17728 25596 17740
rect 24811 17700 25596 17728
rect 24811 17697 24823 17700
rect 24765 17691 24823 17697
rect 25590 17688 25596 17700
rect 25648 17688 25654 17740
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15396 17632 15853 17660
rect 15013 17623 15071 17629
rect 15841 17629 15853 17632
rect 15887 17660 15899 17663
rect 16298 17660 16304 17672
rect 15887 17632 16304 17660
rect 15887 17629 15899 17632
rect 15841 17623 15899 17629
rect 16298 17620 16304 17632
rect 16356 17620 16362 17672
rect 16942 17660 16948 17672
rect 16903 17632 16948 17660
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 21453 17663 21511 17669
rect 21453 17660 21465 17663
rect 21100 17632 21465 17660
rect 21100 17536 21128 17632
rect 21453 17629 21465 17632
rect 21499 17629 21511 17663
rect 21453 17623 21511 17629
rect 23290 17620 23296 17672
rect 23348 17660 23354 17672
rect 23753 17663 23811 17669
rect 23753 17660 23765 17663
rect 23348 17632 23765 17660
rect 23348 17620 23354 17632
rect 23753 17629 23765 17632
rect 23799 17629 23811 17663
rect 23753 17623 23811 17629
rect 23198 17592 23204 17604
rect 23159 17564 23204 17592
rect 23198 17552 23204 17564
rect 23256 17552 23262 17604
rect 10870 17524 10876 17536
rect 10831 17496 10876 17524
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 15286 17524 15292 17536
rect 15247 17496 15292 17524
rect 15286 17484 15292 17496
rect 15344 17484 15350 17536
rect 18322 17524 18328 17536
rect 18283 17496 18328 17524
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 19150 17524 19156 17536
rect 19111 17496 19156 17524
rect 19150 17484 19156 17496
rect 19208 17524 19214 17536
rect 19334 17524 19340 17536
rect 19208 17496 19340 17524
rect 19208 17484 19214 17496
rect 19334 17484 19340 17496
rect 19392 17484 19398 17536
rect 20717 17527 20775 17533
rect 20717 17493 20729 17527
rect 20763 17524 20775 17527
rect 21082 17524 21088 17536
rect 20763 17496 21088 17524
rect 20763 17493 20775 17496
rect 20717 17487 20775 17493
rect 21082 17484 21088 17496
rect 21140 17484 21146 17536
rect 22005 17527 22063 17533
rect 22005 17493 22017 17527
rect 22051 17524 22063 17527
rect 22094 17524 22100 17536
rect 22051 17496 22100 17524
rect 22051 17493 22063 17496
rect 22005 17487 22063 17493
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 24946 17524 24952 17536
rect 24907 17496 24952 17524
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 11790 17320 11796 17332
rect 11751 17292 11796 17320
rect 11790 17280 11796 17292
rect 11848 17320 11854 17332
rect 12161 17323 12219 17329
rect 12161 17320 12173 17323
rect 11848 17292 12173 17320
rect 11848 17280 11854 17292
rect 12161 17289 12173 17292
rect 12207 17289 12219 17323
rect 14734 17320 14740 17332
rect 14695 17292 14740 17320
rect 12161 17283 12219 17289
rect 12176 17252 12204 17283
rect 14734 17280 14740 17292
rect 14792 17280 14798 17332
rect 16298 17320 16304 17332
rect 16259 17292 16304 17320
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 22554 17320 22560 17332
rect 22515 17292 22560 17320
rect 22554 17280 22560 17292
rect 22612 17280 22618 17332
rect 23290 17280 23296 17332
rect 23348 17320 23354 17332
rect 25041 17323 25099 17329
rect 25041 17320 25053 17323
rect 23348 17292 25053 17320
rect 23348 17280 23354 17292
rect 25041 17289 25053 17292
rect 25087 17289 25099 17323
rect 25590 17320 25596 17332
rect 25551 17292 25596 17320
rect 25041 17283 25099 17289
rect 25590 17280 25596 17292
rect 25648 17280 25654 17332
rect 12176 17224 12480 17252
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 11238 17184 11244 17196
rect 10367 17156 11244 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 11238 17144 11244 17156
rect 11296 17184 11302 17196
rect 11422 17184 11428 17196
rect 11296 17156 11428 17184
rect 11296 17144 11302 17156
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 12452 17193 12480 17224
rect 12437 17187 12495 17193
rect 12437 17153 12449 17187
rect 12483 17153 12495 17187
rect 14752 17184 14780 17280
rect 22005 17255 22063 17261
rect 22005 17221 22017 17255
rect 22051 17252 22063 17255
rect 22281 17255 22339 17261
rect 22281 17252 22293 17255
rect 22051 17224 22293 17252
rect 22051 17221 22063 17224
rect 22005 17215 22063 17221
rect 22281 17221 22293 17224
rect 22327 17252 22339 17255
rect 23658 17252 23664 17264
rect 22327 17224 23664 17252
rect 22327 17221 22339 17224
rect 22281 17215 22339 17221
rect 23658 17212 23664 17224
rect 23716 17212 23722 17264
rect 14921 17187 14979 17193
rect 14921 17184 14933 17187
rect 14752 17156 14933 17184
rect 12437 17147 12495 17153
rect 14921 17153 14933 17156
rect 14967 17153 14979 17187
rect 21818 17184 21824 17196
rect 21779 17156 21824 17184
rect 14921 17147 14979 17153
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 10962 17116 10968 17128
rect 10735 17088 10968 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 10962 17076 10968 17088
rect 11020 17116 11026 17128
rect 11020 17088 11459 17116
rect 11020 17076 11026 17088
rect 11149 17051 11207 17057
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 11330 17048 11336 17060
rect 11195 17020 11336 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 11330 17008 11336 17020
rect 11388 17008 11394 17060
rect 10781 16983 10839 16989
rect 10781 16949 10793 16983
rect 10827 16980 10839 16983
rect 11054 16980 11060 16992
rect 10827 16952 11060 16980
rect 10827 16949 10839 16952
rect 10781 16943 10839 16949
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11241 16983 11299 16989
rect 11241 16949 11253 16983
rect 11287 16980 11299 16983
rect 11431 16980 11459 17088
rect 12526 17076 12532 17128
rect 12584 17116 12590 17128
rect 12693 17119 12751 17125
rect 12693 17116 12705 17119
rect 12584 17088 12705 17116
rect 12584 17076 12590 17088
rect 12693 17085 12705 17088
rect 12739 17085 12751 17119
rect 16022 17116 16028 17128
rect 12693 17079 12751 17085
rect 13096 17088 16028 17116
rect 13096 16980 13124 17088
rect 16022 17076 16028 17088
rect 16080 17076 16086 17128
rect 17402 17116 17408 17128
rect 17363 17088 17408 17116
rect 17402 17076 17408 17088
rect 17460 17076 17466 17128
rect 18693 17119 18751 17125
rect 18693 17116 18705 17119
rect 18524 17088 18705 17116
rect 14826 17048 14832 17060
rect 13832 17020 14832 17048
rect 13832 16989 13860 17020
rect 14826 17008 14832 17020
rect 14884 17048 14890 17060
rect 15166 17051 15224 17057
rect 15166 17048 15178 17051
rect 14884 17020 15178 17048
rect 14884 17008 14890 17020
rect 15166 17017 15178 17020
rect 15212 17017 15224 17051
rect 15166 17011 15224 17017
rect 11287 16952 13124 16980
rect 13817 16983 13875 16989
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 13817 16949 13829 16983
rect 13863 16949 13875 16983
rect 13817 16943 13875 16949
rect 14274 16940 14280 16992
rect 14332 16980 14338 16992
rect 14369 16983 14427 16989
rect 14369 16980 14381 16983
rect 14332 16952 14381 16980
rect 14332 16940 14338 16952
rect 14369 16949 14381 16952
rect 14415 16949 14427 16983
rect 16942 16980 16948 16992
rect 16903 16952 16948 16980
rect 14369 16943 14427 16949
rect 16942 16940 16948 16952
rect 17000 16980 17006 16992
rect 18524 16989 18552 17088
rect 18693 17085 18705 17088
rect 18739 17085 18751 17119
rect 18693 17079 18751 17085
rect 20898 17076 20904 17128
rect 20956 17116 20962 17128
rect 23477 17119 23535 17125
rect 23477 17116 23489 17119
rect 20956 17088 23489 17116
rect 20956 17076 20962 17088
rect 23477 17085 23489 17088
rect 23523 17116 23535 17119
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 23523 17088 23673 17116
rect 23523 17085 23535 17088
rect 23477 17079 23535 17085
rect 23661 17085 23673 17088
rect 23707 17085 23719 17119
rect 23661 17079 23719 17085
rect 23928 17119 23986 17125
rect 23928 17085 23940 17119
rect 23974 17116 23986 17119
rect 24762 17116 24768 17128
rect 23974 17088 24768 17116
rect 23974 17085 23986 17088
rect 23928 17079 23986 17085
rect 24762 17076 24768 17088
rect 24820 17076 24826 17128
rect 18960 17051 19018 17057
rect 18960 17017 18972 17051
rect 19006 17048 19018 17051
rect 19058 17048 19064 17060
rect 19006 17020 19064 17048
rect 19006 17017 19018 17020
rect 18960 17011 19018 17017
rect 19058 17008 19064 17020
rect 19116 17008 19122 17060
rect 19334 17008 19340 17060
rect 19392 17048 19398 17060
rect 20993 17051 21051 17057
rect 20993 17048 21005 17051
rect 19392 17020 21005 17048
rect 19392 17008 19398 17020
rect 20993 17017 21005 17020
rect 21039 17048 21051 17051
rect 21358 17048 21364 17060
rect 21039 17020 21364 17048
rect 21039 17017 21051 17020
rect 20993 17011 21051 17017
rect 21358 17008 21364 17020
rect 21416 17008 21422 17060
rect 21545 17051 21603 17057
rect 21545 17017 21557 17051
rect 21591 17048 21603 17051
rect 22554 17048 22560 17060
rect 21591 17020 22560 17048
rect 21591 17017 21603 17020
rect 21545 17011 21603 17017
rect 22554 17008 22560 17020
rect 22612 17008 22618 17060
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 17000 16952 18521 16980
rect 17000 16940 17006 16952
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 18509 16943 18567 16949
rect 19150 16940 19156 16992
rect 19208 16980 19214 16992
rect 20073 16983 20131 16989
rect 20073 16980 20085 16983
rect 19208 16952 20085 16980
rect 19208 16940 19214 16952
rect 20073 16949 20085 16952
rect 20119 16949 20131 16983
rect 21174 16980 21180 16992
rect 21135 16952 21180 16980
rect 20073 16943 20131 16949
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 21634 16980 21640 16992
rect 21547 16952 21640 16980
rect 21634 16940 21640 16952
rect 21692 16980 21698 16992
rect 22005 16983 22063 16989
rect 22005 16980 22017 16983
rect 21692 16952 22017 16980
rect 21692 16940 21698 16952
rect 22005 16949 22017 16952
rect 22051 16949 22063 16983
rect 23014 16980 23020 16992
rect 22975 16952 23020 16980
rect 22005 16943 22063 16949
rect 23014 16940 23020 16952
rect 23072 16940 23078 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 11238 16776 11244 16788
rect 11199 16748 11244 16776
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 12526 16776 12532 16788
rect 12487 16748 12532 16776
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 13725 16779 13783 16785
rect 13725 16745 13737 16779
rect 13771 16776 13783 16779
rect 13998 16776 14004 16788
rect 13771 16748 14004 16776
rect 13771 16745 13783 16748
rect 13725 16739 13783 16745
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 14093 16779 14151 16785
rect 14093 16745 14105 16779
rect 14139 16776 14151 16779
rect 14826 16776 14832 16788
rect 14139 16748 14832 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 14826 16736 14832 16748
rect 14884 16736 14890 16788
rect 15105 16779 15163 16785
rect 15105 16745 15117 16779
rect 15151 16776 15163 16779
rect 15654 16776 15660 16788
rect 15151 16748 15660 16776
rect 15151 16745 15163 16748
rect 15105 16739 15163 16745
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 15838 16736 15844 16788
rect 15896 16776 15902 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 15896 16748 16405 16776
rect 15896 16736 15902 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 18877 16779 18935 16785
rect 18877 16745 18889 16779
rect 18923 16776 18935 16779
rect 19058 16776 19064 16788
rect 18923 16748 19064 16776
rect 18923 16745 18935 16748
rect 18877 16739 18935 16745
rect 11054 16668 11060 16720
rect 11112 16708 11118 16720
rect 11701 16711 11759 16717
rect 11701 16708 11713 16711
rect 11112 16680 11713 16708
rect 11112 16668 11118 16680
rect 11701 16677 11713 16680
rect 11747 16677 11759 16711
rect 12544 16708 12572 16736
rect 14642 16708 14648 16720
rect 11701 16671 11759 16677
rect 11992 16680 12572 16708
rect 14603 16680 14648 16708
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 11330 16640 11336 16652
rect 10919 16612 11336 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 11992 16584 12020 16680
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 15286 16668 15292 16720
rect 15344 16708 15350 16720
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 15344 16680 15761 16708
rect 15344 16668 15350 16680
rect 15749 16677 15761 16680
rect 15795 16677 15807 16711
rect 15749 16671 15807 16677
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15120 16612 15669 16640
rect 11146 16532 11152 16584
rect 11204 16572 11210 16584
rect 11790 16572 11796 16584
rect 11204 16544 11796 16572
rect 11204 16532 11210 16544
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 11974 16572 11980 16584
rect 11887 16544 11980 16572
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 14185 16575 14243 16581
rect 14185 16541 14197 16575
rect 14231 16572 14243 16575
rect 14642 16572 14648 16584
rect 14231 16544 14648 16572
rect 14231 16541 14243 16544
rect 14185 16535 14243 16541
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 14734 16532 14740 16584
rect 14792 16572 14798 16584
rect 15120 16572 15148 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 16408 16640 16436 16739
rect 19058 16736 19064 16748
rect 19116 16736 19122 16788
rect 19518 16736 19524 16788
rect 19576 16776 19582 16788
rect 19797 16779 19855 16785
rect 19797 16776 19809 16779
rect 19576 16748 19809 16776
rect 19576 16736 19582 16748
rect 19797 16745 19809 16748
rect 19843 16745 19855 16779
rect 20346 16776 20352 16788
rect 20307 16748 20352 16776
rect 19797 16739 19855 16745
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 20717 16779 20775 16785
rect 20717 16745 20729 16779
rect 20763 16776 20775 16779
rect 20990 16776 20996 16788
rect 20763 16748 20996 16776
rect 20763 16745 20775 16748
rect 20717 16739 20775 16745
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 22278 16776 22284 16788
rect 22239 16748 22284 16776
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 22925 16779 22983 16785
rect 22925 16745 22937 16779
rect 22971 16776 22983 16779
rect 23477 16779 23535 16785
rect 23477 16776 23489 16779
rect 22971 16748 23489 16776
rect 22971 16745 22983 16748
rect 22925 16739 22983 16745
rect 23477 16745 23489 16748
rect 23523 16776 23535 16779
rect 23566 16776 23572 16788
rect 23523 16748 23572 16776
rect 23523 16745 23535 16748
rect 23477 16739 23535 16745
rect 23566 16736 23572 16748
rect 23624 16736 23630 16788
rect 23658 16736 23664 16788
rect 23716 16776 23722 16788
rect 24118 16776 24124 16788
rect 23716 16748 24124 16776
rect 23716 16736 23722 16748
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 24581 16779 24639 16785
rect 24581 16745 24593 16779
rect 24627 16776 24639 16779
rect 24762 16776 24768 16788
rect 24627 16748 24768 16776
rect 24627 16745 24639 16748
rect 24581 16739 24639 16745
rect 21082 16668 21088 16720
rect 21140 16717 21146 16720
rect 21140 16711 21204 16717
rect 21140 16677 21158 16711
rect 21192 16677 21204 16711
rect 23198 16708 23204 16720
rect 23159 16680 23204 16708
rect 21140 16671 21204 16677
rect 21140 16668 21146 16671
rect 23198 16668 23204 16680
rect 23256 16668 23262 16720
rect 16853 16643 16911 16649
rect 16408 16612 16528 16640
rect 15657 16603 15715 16609
rect 14792 16544 15148 16572
rect 14792 16532 14798 16544
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15804 16544 15853 16572
rect 15804 16532 15810 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 16500 16572 16528 16612
rect 16853 16609 16865 16643
rect 16899 16640 16911 16643
rect 16942 16640 16948 16652
rect 16899 16612 16948 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17126 16649 17132 16652
rect 17120 16640 17132 16649
rect 17039 16612 17132 16640
rect 17120 16603 17132 16612
rect 17184 16640 17190 16652
rect 18322 16640 18328 16652
rect 17184 16612 18328 16640
rect 17126 16600 17132 16603
rect 17184 16600 17190 16612
rect 18322 16600 18328 16612
rect 18380 16600 18386 16652
rect 20898 16640 20904 16652
rect 20859 16612 20904 16640
rect 20898 16600 20904 16612
rect 20956 16600 20962 16652
rect 23474 16600 23480 16652
rect 23532 16640 23538 16652
rect 23845 16643 23903 16649
rect 23845 16640 23857 16643
rect 23532 16612 23857 16640
rect 23532 16600 23538 16612
rect 23845 16609 23857 16612
rect 23891 16640 23903 16643
rect 24210 16640 24216 16652
rect 23891 16612 24216 16640
rect 23891 16609 23903 16612
rect 23845 16603 23903 16609
rect 24210 16600 24216 16612
rect 24268 16600 24274 16652
rect 16758 16572 16764 16584
rect 16500 16544 16764 16572
rect 15841 16535 15899 16541
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 23658 16532 23664 16584
rect 23716 16572 23722 16584
rect 23937 16575 23995 16581
rect 23937 16572 23949 16575
rect 23716 16544 23949 16572
rect 23716 16532 23722 16544
rect 23937 16541 23949 16544
rect 23983 16541 23995 16575
rect 23937 16535 23995 16541
rect 24026 16532 24032 16584
rect 24084 16572 24090 16584
rect 24121 16575 24179 16581
rect 24121 16572 24133 16575
rect 24084 16544 24133 16572
rect 24084 16532 24090 16544
rect 24121 16541 24133 16544
rect 24167 16572 24179 16575
rect 24596 16572 24624 16739
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 25222 16776 25228 16788
rect 25183 16748 25228 16776
rect 25222 16736 25228 16748
rect 25280 16736 25286 16788
rect 25038 16640 25044 16652
rect 24999 16612 25044 16640
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 24167 16544 24624 16572
rect 24167 16541 24179 16544
rect 24121 16535 24179 16541
rect 14274 16464 14280 16516
rect 14332 16504 14338 16516
rect 15289 16507 15347 16513
rect 15289 16504 15301 16507
rect 14332 16476 15301 16504
rect 14332 16464 14338 16476
rect 15289 16473 15301 16476
rect 15335 16473 15347 16507
rect 15289 16467 15347 16473
rect 11333 16439 11391 16445
rect 11333 16405 11345 16439
rect 11379 16436 11391 16439
rect 12434 16436 12440 16448
rect 11379 16408 12440 16436
rect 11379 16405 11391 16408
rect 11333 16399 11391 16405
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 18230 16436 18236 16448
rect 18191 16408 18236 16436
rect 18230 16396 18236 16408
rect 18288 16396 18294 16448
rect 21082 16396 21088 16448
rect 21140 16436 21146 16448
rect 21818 16436 21824 16448
rect 21140 16408 21824 16436
rect 21140 16396 21146 16408
rect 21818 16396 21824 16408
rect 21876 16436 21882 16448
rect 23014 16436 23020 16448
rect 21876 16408 23020 16436
rect 21876 16396 21882 16408
rect 23014 16396 23020 16408
rect 23072 16396 23078 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11149 16235 11207 16241
rect 11149 16232 11161 16235
rect 11112 16204 11161 16232
rect 11112 16192 11118 16204
rect 11149 16201 11161 16204
rect 11195 16201 11207 16235
rect 11149 16195 11207 16201
rect 11885 16235 11943 16241
rect 11885 16201 11897 16235
rect 11931 16232 11943 16235
rect 11974 16232 11980 16244
rect 11931 16204 11980 16232
rect 11931 16201 11943 16204
rect 11885 16195 11943 16201
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 14185 16235 14243 16241
rect 14185 16201 14197 16235
rect 14231 16232 14243 16235
rect 14645 16235 14703 16241
rect 14645 16232 14657 16235
rect 14231 16204 14657 16232
rect 14231 16201 14243 16204
rect 14185 16195 14243 16201
rect 14645 16201 14657 16204
rect 14691 16232 14703 16235
rect 14734 16232 14740 16244
rect 14691 16204 14740 16232
rect 14691 16201 14703 16204
rect 14645 16195 14703 16201
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 15746 16232 15752 16244
rect 15707 16204 15752 16232
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 18509 16235 18567 16241
rect 18509 16201 18521 16235
rect 18555 16232 18567 16235
rect 19150 16232 19156 16244
rect 18555 16204 19156 16232
rect 18555 16201 18567 16204
rect 18509 16195 18567 16201
rect 19150 16192 19156 16204
rect 19208 16192 19214 16244
rect 20898 16192 20904 16244
rect 20956 16232 20962 16244
rect 21177 16235 21235 16241
rect 21177 16232 21189 16235
rect 20956 16204 21189 16232
rect 20956 16192 20962 16204
rect 21177 16201 21189 16204
rect 21223 16232 21235 16235
rect 21910 16232 21916 16244
rect 21223 16204 21916 16232
rect 21223 16201 21235 16204
rect 21177 16195 21235 16201
rect 21910 16192 21916 16204
rect 21968 16192 21974 16244
rect 23477 16235 23535 16241
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 24026 16232 24032 16244
rect 23523 16204 24032 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 24026 16192 24032 16204
rect 24084 16192 24090 16244
rect 24210 16232 24216 16244
rect 24171 16204 24216 16232
rect 24210 16192 24216 16204
rect 24268 16192 24274 16244
rect 25038 16192 25044 16244
rect 25096 16232 25102 16244
rect 25501 16235 25559 16241
rect 25501 16232 25513 16235
rect 25096 16204 25513 16232
rect 25096 16192 25102 16204
rect 25501 16201 25513 16204
rect 25547 16201 25559 16235
rect 25501 16195 25559 16201
rect 11790 16124 11796 16176
rect 11848 16164 11854 16176
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 11848 16136 12173 16164
rect 11848 16124 11854 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 17126 16164 17132 16176
rect 12161 16127 12219 16133
rect 17052 16136 17132 16164
rect 11330 16096 11336 16108
rect 11291 16068 11336 16096
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 14826 16056 14832 16108
rect 14884 16096 14890 16108
rect 17052 16105 17080 16136
rect 17126 16124 17132 16136
rect 17184 16124 17190 16176
rect 21729 16167 21787 16173
rect 21729 16164 21741 16167
rect 19076 16136 21741 16164
rect 19076 16105 19104 16136
rect 21729 16133 21741 16136
rect 21775 16133 21787 16167
rect 21729 16127 21787 16133
rect 15197 16099 15255 16105
rect 15197 16096 15209 16099
rect 14884 16068 15209 16096
rect 14884 16056 14890 16068
rect 15197 16065 15209 16068
rect 15243 16065 15255 16099
rect 15197 16059 15255 16065
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16096 17923 16099
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 17911 16068 19073 16096
rect 17911 16065 17923 16068
rect 17865 16059 17923 16065
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 19150 16056 19156 16108
rect 19208 16096 19214 16108
rect 19705 16099 19763 16105
rect 19208 16068 19253 16096
rect 19208 16056 19214 16068
rect 19705 16065 19717 16099
rect 19751 16096 19763 16099
rect 20717 16099 20775 16105
rect 20717 16096 20729 16099
rect 19751 16068 20729 16096
rect 19751 16065 19763 16068
rect 19705 16059 19763 16065
rect 20717 16065 20729 16068
rect 20763 16096 20775 16099
rect 21082 16096 21088 16108
rect 20763 16068 21088 16096
rect 20763 16065 20775 16068
rect 20717 16059 20775 16065
rect 21082 16056 21088 16068
rect 21140 16096 21146 16108
rect 21545 16099 21603 16105
rect 21545 16096 21557 16099
rect 21140 16068 21557 16096
rect 21140 16056 21146 16068
rect 21545 16065 21557 16068
rect 21591 16065 21603 16099
rect 21545 16059 21603 16065
rect 21818 16056 21824 16108
rect 21876 16096 21882 16108
rect 22278 16096 22284 16108
rect 21876 16068 22284 16096
rect 21876 16056 21882 16068
rect 22278 16056 22284 16068
rect 22336 16056 22342 16108
rect 12434 16028 12440 16040
rect 12395 16000 12440 16028
rect 12434 15988 12440 16000
rect 12492 16028 12498 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12492 16000 12909 16028
rect 12492 15988 12498 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 14642 15988 14648 16040
rect 14700 16028 14706 16040
rect 15013 16031 15071 16037
rect 15013 16028 15025 16031
rect 14700 16000 15025 16028
rect 14700 15988 14706 16000
rect 15013 15997 15025 16000
rect 15059 15997 15071 16031
rect 16758 16028 16764 16040
rect 16719 16000 16764 16028
rect 15013 15991 15071 15997
rect 16758 15988 16764 16000
rect 16816 15988 16822 16040
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 16028 19027 16031
rect 19242 16028 19248 16040
rect 19015 16000 19248 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 19242 15988 19248 16000
rect 19300 15988 19306 16040
rect 20625 16031 20683 16037
rect 20625 16028 20637 16031
rect 20088 16000 20637 16028
rect 16114 15920 16120 15972
rect 16172 15960 16178 15972
rect 16301 15963 16359 15969
rect 16301 15960 16313 15963
rect 16172 15932 16313 15960
rect 16172 15920 16178 15932
rect 16301 15929 16313 15932
rect 16347 15960 16359 15963
rect 16853 15963 16911 15969
rect 16853 15960 16865 15963
rect 16347 15932 16865 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 16853 15929 16865 15932
rect 16899 15960 16911 15963
rect 18690 15960 18696 15972
rect 16899 15932 18696 15960
rect 16899 15929 16911 15932
rect 16853 15923 16911 15929
rect 18690 15920 18696 15932
rect 18748 15920 18754 15972
rect 20088 15904 20116 16000
rect 20625 15997 20637 16000
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 21174 15988 21180 16040
rect 21232 16028 21238 16040
rect 22097 16031 22155 16037
rect 22097 16028 22109 16031
rect 21232 16000 22109 16028
rect 21232 15988 21238 16000
rect 22097 15997 22109 16000
rect 22143 15997 22155 16031
rect 24578 16028 24584 16040
rect 24539 16000 24584 16028
rect 22097 15991 22155 15997
rect 24578 15988 24584 16000
rect 24636 16028 24642 16040
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24636 16000 25145 16028
rect 24636 15988 24642 16000
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 22189 15963 22247 15969
rect 22189 15960 22201 15963
rect 20180 15932 22201 15960
rect 12621 15895 12679 15901
rect 12621 15861 12633 15895
rect 12667 15892 12679 15895
rect 13722 15892 13728 15904
rect 12667 15864 13728 15892
rect 12667 15861 12679 15864
rect 12621 15855 12679 15861
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14461 15895 14519 15901
rect 14461 15892 14473 15895
rect 14240 15864 14473 15892
rect 14240 15852 14246 15864
rect 14461 15861 14473 15864
rect 14507 15892 14519 15895
rect 15105 15895 15163 15901
rect 15105 15892 15117 15895
rect 14507 15864 15117 15892
rect 14507 15861 14519 15864
rect 14461 15855 14519 15861
rect 15105 15861 15117 15864
rect 15151 15892 15163 15895
rect 15194 15892 15200 15904
rect 15151 15864 15200 15892
rect 15151 15861 15163 15864
rect 15105 15855 15163 15861
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 16390 15892 16396 15904
rect 16351 15864 16396 15892
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 16942 15852 16948 15904
rect 17000 15892 17006 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 17000 15864 17417 15892
rect 17000 15852 17006 15864
rect 17405 15861 17417 15864
rect 17451 15861 17463 15895
rect 17405 15855 17463 15861
rect 18601 15895 18659 15901
rect 18601 15861 18613 15895
rect 18647 15892 18659 15895
rect 19150 15892 19156 15904
rect 18647 15864 19156 15892
rect 18647 15861 18659 15864
rect 18601 15855 18659 15861
rect 19150 15852 19156 15864
rect 19208 15852 19214 15904
rect 20070 15892 20076 15904
rect 20031 15864 20076 15892
rect 20070 15852 20076 15864
rect 20128 15852 20134 15904
rect 20180 15901 20208 15932
rect 22189 15929 22201 15932
rect 22235 15960 22247 15963
rect 22741 15963 22799 15969
rect 22741 15960 22753 15963
rect 22235 15932 22753 15960
rect 22235 15929 22247 15932
rect 22189 15923 22247 15929
rect 22741 15929 22753 15932
rect 22787 15929 22799 15963
rect 22741 15923 22799 15929
rect 20165 15895 20223 15901
rect 20165 15861 20177 15895
rect 20211 15861 20223 15895
rect 20530 15892 20536 15904
rect 20491 15864 20536 15892
rect 20165 15855 20223 15861
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 23658 15852 23664 15904
rect 23716 15892 23722 15904
rect 23845 15895 23903 15901
rect 23845 15892 23857 15895
rect 23716 15864 23857 15892
rect 23716 15852 23722 15864
rect 23845 15861 23857 15864
rect 23891 15861 23903 15895
rect 24762 15892 24768 15904
rect 24723 15864 24768 15892
rect 23845 15855 23903 15861
rect 24762 15852 24768 15864
rect 24820 15852 24826 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 14642 15688 14648 15700
rect 14603 15660 14648 15688
rect 14642 15648 14648 15660
rect 14700 15648 14706 15700
rect 15102 15688 15108 15700
rect 15063 15660 15108 15688
rect 15102 15648 15108 15660
rect 15160 15648 15166 15700
rect 16669 15691 16727 15697
rect 16669 15657 16681 15691
rect 16715 15688 16727 15691
rect 17034 15688 17040 15700
rect 16715 15660 17040 15688
rect 16715 15657 16727 15660
rect 16669 15651 16727 15657
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 19153 15691 19211 15697
rect 19153 15657 19165 15691
rect 19199 15688 19211 15691
rect 19242 15688 19248 15700
rect 19199 15660 19248 15688
rect 19199 15657 19211 15660
rect 19153 15651 19211 15657
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 20257 15691 20315 15697
rect 20257 15657 20269 15691
rect 20303 15688 20315 15691
rect 20530 15688 20536 15700
rect 20303 15660 20536 15688
rect 20303 15657 20315 15660
rect 20257 15651 20315 15657
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 21174 15648 21180 15700
rect 21232 15688 21238 15700
rect 21361 15691 21419 15697
rect 21361 15688 21373 15691
rect 21232 15660 21373 15688
rect 21232 15648 21238 15660
rect 21361 15657 21373 15660
rect 21407 15657 21419 15691
rect 21818 15688 21824 15700
rect 21779 15660 21824 15688
rect 21361 15651 21419 15657
rect 21818 15648 21824 15660
rect 21876 15648 21882 15700
rect 23014 15648 23020 15700
rect 23072 15688 23078 15700
rect 23293 15691 23351 15697
rect 23293 15688 23305 15691
rect 23072 15660 23305 15688
rect 23072 15648 23078 15660
rect 23293 15657 23305 15660
rect 23339 15657 23351 15691
rect 23293 15651 23351 15657
rect 14185 15555 14243 15561
rect 14185 15521 14197 15555
rect 14231 15552 14243 15555
rect 14274 15552 14280 15564
rect 14231 15524 14280 15552
rect 14231 15521 14243 15524
rect 14185 15515 14243 15521
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 15746 15512 15752 15564
rect 15804 15552 15810 15564
rect 15933 15555 15991 15561
rect 15933 15552 15945 15555
rect 15804 15524 15945 15552
rect 15804 15512 15810 15524
rect 15933 15521 15945 15524
rect 15979 15521 15991 15555
rect 16390 15552 16396 15564
rect 15933 15515 15991 15521
rect 16040 15524 16396 15552
rect 14826 15444 14832 15496
rect 14884 15484 14890 15496
rect 16040 15493 16068 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 17402 15561 17408 15564
rect 17396 15552 17408 15561
rect 17363 15524 17408 15552
rect 17396 15515 17408 15524
rect 17402 15512 17408 15515
rect 17460 15512 17466 15564
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15552 20959 15555
rect 21358 15552 21364 15564
rect 20947 15524 21364 15552
rect 20947 15521 20959 15524
rect 20901 15515 20959 15521
rect 21358 15512 21364 15524
rect 21416 15512 21422 15564
rect 21910 15552 21916 15564
rect 21871 15524 21916 15552
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 22186 15561 22192 15564
rect 22180 15515 22192 15561
rect 22244 15552 22250 15564
rect 24578 15552 24584 15564
rect 22244 15524 22280 15552
rect 24539 15524 24584 15552
rect 22186 15512 22192 15515
rect 22244 15512 22250 15524
rect 24578 15512 24584 15524
rect 24636 15512 24642 15564
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 14884 15456 16037 15484
rect 14884 15444 14890 15456
rect 16025 15453 16037 15456
rect 16071 15453 16083 15487
rect 16206 15484 16212 15496
rect 16167 15456 16212 15484
rect 16025 15447 16083 15453
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 16942 15444 16948 15496
rect 17000 15484 17006 15496
rect 17129 15487 17187 15493
rect 17129 15484 17141 15487
rect 17000 15456 17141 15484
rect 17000 15444 17006 15456
rect 17129 15453 17141 15456
rect 17175 15453 17187 15487
rect 17129 15447 17187 15453
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19613 15487 19671 15493
rect 19613 15484 19625 15487
rect 19484 15456 19625 15484
rect 19484 15444 19490 15456
rect 19613 15453 19625 15456
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 14369 15419 14427 15425
rect 14369 15385 14381 15419
rect 14415 15416 14427 15419
rect 15102 15416 15108 15428
rect 14415 15388 15108 15416
rect 14415 15385 14427 15388
rect 14369 15379 14427 15385
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 24762 15416 24768 15428
rect 24723 15388 24768 15416
rect 24762 15376 24768 15388
rect 24820 15376 24826 15428
rect 15286 15308 15292 15360
rect 15344 15348 15350 15360
rect 15565 15351 15623 15357
rect 15565 15348 15577 15351
rect 15344 15320 15577 15348
rect 15344 15308 15350 15320
rect 15565 15317 15577 15320
rect 15611 15348 15623 15351
rect 16482 15348 16488 15360
rect 15611 15320 16488 15348
rect 15611 15317 15623 15320
rect 15565 15311 15623 15317
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 18509 15351 18567 15357
rect 18509 15317 18521 15351
rect 18555 15348 18567 15351
rect 18598 15348 18604 15360
rect 18555 15320 18604 15348
rect 18555 15317 18567 15320
rect 18509 15311 18567 15317
rect 18598 15308 18604 15320
rect 18656 15308 18662 15360
rect 21085 15351 21143 15357
rect 21085 15317 21097 15351
rect 21131 15348 21143 15351
rect 21542 15348 21548 15360
rect 21131 15320 21548 15348
rect 21131 15317 21143 15320
rect 21085 15311 21143 15317
rect 21542 15308 21548 15320
rect 21600 15308 21606 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 14274 15144 14280 15156
rect 14235 15116 14280 15144
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 14737 15147 14795 15153
rect 14737 15113 14749 15147
rect 14783 15144 14795 15147
rect 14826 15144 14832 15156
rect 14783 15116 14832 15144
rect 14783 15113 14795 15116
rect 14737 15107 14795 15113
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 15746 15144 15752 15156
rect 15707 15116 15752 15144
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 16209 15147 16267 15153
rect 16209 15113 16221 15147
rect 16255 15144 16267 15147
rect 16390 15144 16396 15156
rect 16255 15116 16396 15144
rect 16255 15113 16267 15116
rect 16209 15107 16267 15113
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 20806 15144 20812 15156
rect 20767 15116 20812 15144
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 21910 15144 21916 15156
rect 21871 15116 21916 15144
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 22186 15104 22192 15156
rect 22244 15144 22250 15156
rect 22281 15147 22339 15153
rect 22281 15144 22293 15147
rect 22244 15116 22293 15144
rect 22244 15104 22250 15116
rect 22281 15113 22293 15116
rect 22327 15113 22339 15147
rect 22738 15144 22744 15156
rect 22699 15116 22744 15144
rect 22281 15107 22339 15113
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 24489 15147 24547 15153
rect 24489 15113 24501 15147
rect 24535 15144 24547 15147
rect 24670 15144 24676 15156
rect 24535 15116 24676 15144
rect 24535 15113 24547 15116
rect 24489 15107 24547 15113
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16632 14980 16681 15008
rect 16632 14968 16638 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16761 15011 16819 15017
rect 16761 14977 16773 15011
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 12989 14943 13047 14949
rect 12989 14940 13001 14943
rect 12676 14912 13001 14940
rect 12676 14900 12682 14912
rect 12989 14909 13001 14912
rect 13035 14940 13047 14943
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 13035 14912 13461 14940
rect 13035 14909 13047 14912
rect 12989 14903 13047 14909
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14940 16175 14943
rect 16776 14940 16804 14971
rect 17402 14940 17408 14952
rect 16163 14912 17408 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 17402 14900 17408 14912
rect 17460 14940 17466 14952
rect 17589 14943 17647 14949
rect 17589 14940 17601 14943
rect 17460 14912 17601 14940
rect 17460 14900 17466 14912
rect 17589 14909 17601 14912
rect 17635 14909 17647 14943
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 17589 14903 17647 14909
rect 18340 14912 18521 14940
rect 15105 14875 15163 14881
rect 15105 14841 15117 14875
rect 15151 14872 15163 14875
rect 16206 14872 16212 14884
rect 15151 14844 16212 14872
rect 15151 14841 15163 14844
rect 15105 14835 15163 14841
rect 16206 14832 16212 14844
rect 16264 14832 16270 14884
rect 13170 14804 13176 14816
rect 13131 14776 13176 14804
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 15194 14804 15200 14816
rect 15155 14776 15200 14804
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 16574 14804 16580 14816
rect 16535 14776 16580 14804
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 18340 14813 18368 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 18598 14900 18604 14952
rect 18656 14940 18662 14952
rect 18765 14943 18823 14949
rect 18765 14940 18777 14943
rect 18656 14912 18777 14940
rect 18656 14900 18662 14912
rect 18765 14909 18777 14912
rect 18811 14909 18823 14943
rect 18765 14903 18823 14909
rect 20806 14900 20812 14952
rect 20864 14940 20870 14952
rect 20993 14943 21051 14949
rect 20993 14940 21005 14943
rect 20864 14912 21005 14940
rect 20864 14900 20870 14912
rect 20993 14909 21005 14912
rect 21039 14909 21051 14943
rect 20993 14903 21051 14909
rect 22557 14943 22615 14949
rect 22557 14909 22569 14943
rect 22603 14940 22615 14943
rect 24578 14940 24584 14952
rect 22603 14912 23152 14940
rect 24539 14912 24584 14940
rect 22603 14909 22615 14912
rect 22557 14903 22615 14909
rect 21358 14832 21364 14884
rect 21416 14872 21422 14884
rect 21453 14875 21511 14881
rect 21453 14872 21465 14875
rect 21416 14844 21465 14872
rect 21416 14832 21422 14844
rect 21453 14841 21465 14844
rect 21499 14841 21511 14875
rect 21453 14835 21511 14841
rect 23124 14816 23152 14912
rect 24578 14900 24584 14912
rect 24636 14940 24642 14952
rect 25133 14943 25191 14949
rect 25133 14940 25145 14943
rect 24636 14912 25145 14940
rect 24636 14900 24642 14912
rect 25133 14909 25145 14912
rect 25179 14909 25191 14943
rect 25133 14903 25191 14909
rect 17221 14807 17279 14813
rect 17221 14804 17233 14807
rect 17000 14776 17233 14804
rect 17000 14764 17006 14776
rect 17221 14773 17233 14776
rect 17267 14804 17279 14807
rect 18325 14807 18383 14813
rect 18325 14804 18337 14807
rect 17267 14776 18337 14804
rect 17267 14773 17279 14776
rect 17221 14767 17279 14773
rect 18325 14773 18337 14776
rect 18371 14773 18383 14807
rect 18325 14767 18383 14773
rect 19889 14807 19947 14813
rect 19889 14773 19901 14807
rect 19935 14804 19947 14807
rect 19978 14804 19984 14816
rect 19935 14776 19984 14804
rect 19935 14773 19947 14776
rect 19889 14767 19947 14773
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 20898 14764 20904 14816
rect 20956 14804 20962 14816
rect 21177 14807 21235 14813
rect 21177 14804 21189 14807
rect 20956 14776 21189 14804
rect 20956 14764 20962 14776
rect 21177 14773 21189 14776
rect 21223 14773 21235 14807
rect 21177 14767 21235 14773
rect 21910 14764 21916 14816
rect 21968 14804 21974 14816
rect 22738 14804 22744 14816
rect 21968 14776 22744 14804
rect 21968 14764 21974 14776
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 23106 14804 23112 14816
rect 23067 14776 23112 14804
rect 23106 14764 23112 14776
rect 23164 14764 23170 14816
rect 24762 14804 24768 14816
rect 24723 14776 24768 14804
rect 24762 14764 24768 14776
rect 24820 14764 24826 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 15749 14603 15807 14609
rect 15749 14600 15761 14603
rect 15252 14572 15761 14600
rect 15252 14560 15258 14572
rect 15749 14569 15761 14572
rect 15795 14600 15807 14603
rect 16114 14600 16120 14612
rect 15795 14572 16120 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 17402 14600 17408 14612
rect 17363 14572 17408 14600
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 18141 14603 18199 14609
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18598 14600 18604 14612
rect 18187 14572 18604 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 19058 14600 19064 14612
rect 19019 14572 19064 14600
rect 19058 14560 19064 14572
rect 19116 14560 19122 14612
rect 19426 14600 19432 14612
rect 19387 14572 19432 14600
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 25409 14603 25467 14609
rect 25409 14600 25421 14603
rect 24912 14572 25421 14600
rect 24912 14560 24918 14572
rect 25409 14569 25421 14572
rect 25455 14569 25467 14603
rect 25409 14563 25467 14569
rect 15105 14535 15163 14541
rect 15105 14501 15117 14535
rect 15151 14532 15163 14535
rect 15286 14532 15292 14544
rect 15151 14504 15292 14532
rect 15151 14501 15163 14504
rect 15105 14495 15163 14501
rect 15286 14492 15292 14504
rect 15344 14492 15350 14544
rect 16206 14492 16212 14544
rect 16264 14541 16270 14544
rect 16264 14535 16328 14541
rect 16264 14501 16282 14535
rect 16316 14532 16328 14535
rect 16390 14532 16396 14544
rect 16316 14504 16396 14532
rect 16316 14501 16328 14504
rect 16264 14495 16328 14501
rect 16264 14492 16270 14495
rect 16390 14492 16396 14504
rect 16448 14492 16454 14544
rect 20990 14492 20996 14544
rect 21048 14532 21054 14544
rect 21048 14504 25268 14532
rect 21048 14492 21054 14504
rect 13078 14464 13084 14476
rect 13039 14436 13084 14464
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 13228 14436 14105 14464
rect 13228 14424 13234 14436
rect 14093 14433 14105 14436
rect 14139 14464 14151 14467
rect 14642 14464 14648 14476
rect 14139 14436 14648 14464
rect 14139 14433 14151 14436
rect 14093 14427 14151 14433
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 16850 14464 16856 14476
rect 16071 14436 16856 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 20898 14464 20904 14476
rect 20859 14436 20904 14464
rect 20898 14424 20904 14436
rect 20956 14424 20962 14476
rect 23008 14467 23066 14473
rect 23008 14433 23020 14467
rect 23054 14464 23066 14467
rect 23290 14464 23296 14476
rect 23054 14436 23296 14464
rect 23054 14433 23066 14436
rect 23008 14427 23066 14433
rect 23290 14424 23296 14436
rect 23348 14424 23354 14476
rect 25240 14473 25268 14504
rect 25225 14467 25283 14473
rect 25225 14433 25237 14467
rect 25271 14464 25283 14467
rect 25774 14464 25780 14476
rect 25271 14436 25780 14464
rect 25271 14433 25283 14436
rect 25225 14427 25283 14433
rect 25774 14424 25780 14436
rect 25832 14424 25838 14476
rect 18046 14356 18052 14408
rect 18104 14396 18110 14408
rect 18969 14399 19027 14405
rect 18969 14396 18981 14399
rect 18104 14368 18981 14396
rect 18104 14356 18110 14368
rect 18969 14365 18981 14368
rect 19015 14396 19027 14399
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 19015 14368 19533 14396
rect 19015 14365 19027 14368
rect 18969 14359 19027 14365
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14365 19671 14399
rect 22738 14396 22744 14408
rect 22699 14368 22744 14396
rect 19613 14359 19671 14365
rect 14274 14328 14280 14340
rect 14235 14300 14280 14328
rect 14274 14288 14280 14300
rect 14332 14288 14338 14340
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 19628 14328 19656 14359
rect 22738 14356 22744 14368
rect 22796 14356 22802 14408
rect 19978 14328 19984 14340
rect 19392 14300 19984 14328
rect 19392 14288 19398 14300
rect 19978 14288 19984 14300
rect 20036 14328 20042 14340
rect 20073 14331 20131 14337
rect 20073 14328 20085 14331
rect 20036 14300 20085 14328
rect 20036 14288 20042 14300
rect 20073 14297 20085 14300
rect 20119 14297 20131 14331
rect 20073 14291 20131 14297
rect 13262 14260 13268 14272
rect 13223 14232 13268 14260
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 21082 14260 21088 14272
rect 21043 14232 21088 14260
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 24118 14260 24124 14272
rect 24079 14232 24124 14260
rect 24118 14220 24124 14232
rect 24176 14220 24182 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 13078 14056 13084 14068
rect 13039 14028 13084 14056
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 14642 14056 14648 14068
rect 14603 14028 14648 14056
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 15749 14059 15807 14065
rect 15749 14025 15761 14059
rect 15795 14056 15807 14059
rect 16574 14056 16580 14068
rect 15795 14028 16580 14056
rect 15795 14025 15807 14028
rect 15749 14019 15807 14025
rect 16574 14016 16580 14028
rect 16632 14056 16638 14068
rect 17129 14059 17187 14065
rect 17129 14056 17141 14059
rect 16632 14028 17141 14056
rect 16632 14016 16638 14028
rect 17129 14025 17141 14028
rect 17175 14025 17187 14059
rect 18046 14056 18052 14068
rect 18007 14028 18052 14056
rect 17129 14019 17187 14025
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 19153 14059 19211 14065
rect 19153 14025 19165 14059
rect 19199 14056 19211 14059
rect 19426 14056 19432 14068
rect 19199 14028 19432 14056
rect 19199 14025 19211 14028
rect 19153 14019 19211 14025
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 20898 14016 20904 14068
rect 20956 14056 20962 14068
rect 21545 14059 21603 14065
rect 21545 14056 21557 14059
rect 20956 14028 21557 14056
rect 20956 14016 20962 14028
rect 21545 14025 21557 14028
rect 21591 14025 21603 14059
rect 21545 14019 21603 14025
rect 22738 14016 22744 14068
rect 22796 14056 22802 14068
rect 23017 14059 23075 14065
rect 23017 14056 23029 14059
rect 22796 14028 23029 14056
rect 22796 14016 22802 14028
rect 23017 14025 23029 14028
rect 23063 14025 23075 14059
rect 23017 14019 23075 14025
rect 23106 14016 23112 14068
rect 23164 14056 23170 14068
rect 23661 14059 23719 14065
rect 23661 14056 23673 14059
rect 23164 14028 23673 14056
rect 23164 14016 23170 14028
rect 23661 14025 23673 14028
rect 23707 14025 23719 14059
rect 25774 14056 25780 14068
rect 25735 14028 25780 14056
rect 23661 14019 23719 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 14369 13991 14427 13997
rect 14369 13957 14381 13991
rect 14415 13988 14427 13991
rect 14550 13988 14556 14000
rect 14415 13960 14556 13988
rect 14415 13957 14427 13960
rect 14369 13951 14427 13957
rect 14550 13948 14556 13960
rect 14608 13948 14614 14000
rect 15289 13991 15347 13997
rect 15289 13957 15301 13991
rect 15335 13988 15347 13991
rect 15335 13960 16436 13988
rect 15335 13957 15347 13960
rect 15289 13951 15347 13957
rect 16408 13932 16436 13960
rect 22278 13948 22284 14000
rect 22336 13988 22342 14000
rect 23385 13991 23443 13997
rect 23385 13988 23397 13991
rect 22336 13960 23397 13988
rect 22336 13948 22342 13960
rect 23385 13957 23397 13960
rect 23431 13988 23443 13991
rect 24118 13988 24124 14000
rect 23431 13960 24124 13988
rect 23431 13957 23443 13960
rect 23385 13951 23443 13957
rect 24118 13948 24124 13960
rect 24176 13988 24182 14000
rect 25406 13988 25412 14000
rect 24176 13960 24256 13988
rect 25367 13960 25412 13988
rect 24176 13948 24182 13960
rect 16209 13923 16267 13929
rect 16209 13920 16221 13923
rect 15580 13892 16221 13920
rect 15580 13864 15608 13892
rect 16209 13889 16221 13892
rect 16255 13889 16267 13923
rect 16390 13920 16396 13932
rect 16351 13892 16396 13920
rect 16209 13883 16267 13889
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 18598 13920 18604 13932
rect 18559 13892 18604 13920
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 19334 13880 19340 13932
rect 19392 13920 19398 13932
rect 24228 13929 24256 13960
rect 25406 13948 25412 13960
rect 25464 13948 25470 14000
rect 24213 13923 24271 13929
rect 19392 13892 19748 13920
rect 19392 13880 19398 13892
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13872 13824 14013 13852
rect 13872 13812 13878 13824
rect 14001 13821 14013 13824
rect 14047 13852 14059 13855
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 14047 13824 14197 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 15562 13852 15568 13864
rect 15523 13824 15568 13852
rect 14185 13815 14243 13821
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 16114 13852 16120 13864
rect 16075 13824 16120 13852
rect 16114 13812 16120 13824
rect 16172 13812 16178 13864
rect 16853 13855 16911 13861
rect 16853 13821 16865 13855
rect 16899 13852 16911 13855
rect 16942 13852 16948 13864
rect 16899 13824 16948 13852
rect 16899 13821 16911 13824
rect 16853 13815 16911 13821
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 18012 13824 18521 13852
rect 18012 13812 18018 13824
rect 18509 13821 18521 13824
rect 18555 13821 18567 13855
rect 18509 13815 18567 13821
rect 19058 13812 19064 13864
rect 19116 13852 19122 13864
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19116 13824 19533 13852
rect 19116 13812 19122 13824
rect 19521 13821 19533 13824
rect 19567 13852 19579 13855
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19567 13824 19625 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 19613 13821 19625 13824
rect 19659 13821 19671 13855
rect 19720 13852 19748 13892
rect 24213 13889 24225 13923
rect 24259 13889 24271 13923
rect 25038 13920 25044 13932
rect 24999 13892 25044 13920
rect 24213 13883 24271 13889
rect 25038 13880 25044 13892
rect 25096 13920 25102 13932
rect 25096 13892 25268 13920
rect 25096 13880 25102 13892
rect 19869 13855 19927 13861
rect 19869 13852 19881 13855
rect 19720 13824 19881 13852
rect 19613 13815 19671 13821
rect 19869 13821 19881 13824
rect 19915 13821 19927 13855
rect 22738 13852 22744 13864
rect 19869 13815 19927 13821
rect 19996 13824 22744 13852
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 17773 13787 17831 13793
rect 17773 13784 17785 13787
rect 11296 13756 17785 13784
rect 11296 13744 11302 13756
rect 17773 13753 17785 13756
rect 17819 13784 17831 13787
rect 18417 13787 18475 13793
rect 18417 13784 18429 13787
rect 17819 13756 18429 13784
rect 17819 13753 17831 13756
rect 17773 13747 17831 13753
rect 18417 13753 18429 13756
rect 18463 13753 18475 13787
rect 19628 13784 19656 13815
rect 19996 13784 20024 13824
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 25240 13861 25268 13892
rect 25225 13855 25283 13861
rect 25225 13821 25237 13855
rect 25271 13821 25283 13855
rect 25225 13815 25283 13821
rect 19628 13756 20024 13784
rect 22465 13787 22523 13793
rect 18417 13747 18475 13753
rect 22465 13753 22477 13787
rect 22511 13784 22523 13787
rect 23290 13784 23296 13796
rect 22511 13756 23296 13784
rect 22511 13753 22523 13756
rect 22465 13747 22523 13753
rect 23290 13744 23296 13756
rect 23348 13744 23354 13796
rect 15930 13676 15936 13728
rect 15988 13716 15994 13728
rect 16390 13716 16396 13728
rect 15988 13688 16396 13716
rect 15988 13676 15994 13688
rect 16390 13676 16396 13688
rect 16448 13676 16454 13728
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 20990 13716 20996 13728
rect 20036 13688 20996 13716
rect 20036 13676 20042 13688
rect 20990 13676 20996 13688
rect 21048 13676 21054 13728
rect 22554 13716 22560 13728
rect 22515 13688 22560 13716
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 24026 13716 24032 13728
rect 23987 13688 24032 13716
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 24118 13676 24124 13728
rect 24176 13716 24182 13728
rect 24176 13688 24221 13716
rect 24176 13676 24182 13688
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13964 13484 14105 13512
rect 13964 13472 13970 13484
rect 14093 13481 14105 13484
rect 14139 13512 14151 13515
rect 14826 13512 14832 13524
rect 14139 13484 14832 13512
rect 14139 13481 14151 13484
rect 14093 13475 14151 13481
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 15473 13515 15531 13521
rect 15473 13481 15485 13515
rect 15519 13512 15531 13515
rect 16853 13515 16911 13521
rect 16853 13512 16865 13515
rect 15519 13484 16865 13512
rect 15519 13481 15531 13484
rect 15473 13475 15531 13481
rect 16853 13481 16865 13484
rect 16899 13512 16911 13515
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 16899 13484 17417 13512
rect 16899 13481 16911 13484
rect 16853 13475 16911 13481
rect 17405 13481 17417 13484
rect 17451 13481 17463 13515
rect 17405 13475 17463 13481
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18049 13515 18107 13521
rect 18049 13512 18061 13515
rect 18012 13484 18061 13512
rect 18012 13472 18018 13484
rect 18049 13481 18061 13484
rect 18095 13481 18107 13515
rect 18049 13475 18107 13481
rect 19153 13515 19211 13521
rect 19153 13481 19165 13515
rect 19199 13512 19211 13515
rect 19334 13512 19340 13524
rect 19199 13484 19340 13512
rect 19199 13481 19211 13484
rect 19153 13475 19211 13481
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 19518 13472 19524 13524
rect 19576 13512 19582 13524
rect 19613 13515 19671 13521
rect 19613 13512 19625 13515
rect 19576 13484 19625 13512
rect 19576 13472 19582 13484
rect 19613 13481 19625 13484
rect 19659 13512 19671 13515
rect 20162 13512 20168 13524
rect 19659 13484 20168 13512
rect 19659 13481 19671 13484
rect 19613 13475 19671 13481
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 22186 13512 22192 13524
rect 22147 13484 22192 13512
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22554 13472 22560 13524
rect 22612 13512 22618 13524
rect 23014 13512 23020 13524
rect 22612 13484 23020 13512
rect 22612 13472 22618 13484
rect 23014 13472 23020 13484
rect 23072 13472 23078 13524
rect 23106 13472 23112 13524
rect 23164 13512 23170 13524
rect 23753 13515 23811 13521
rect 23164 13484 23209 13512
rect 23164 13472 23170 13484
rect 23753 13481 23765 13515
rect 23799 13512 23811 13515
rect 23842 13512 23848 13524
rect 23799 13484 23848 13512
rect 23799 13481 23811 13484
rect 23753 13475 23811 13481
rect 23842 13472 23848 13484
rect 23900 13512 23906 13524
rect 24118 13512 24124 13524
rect 23900 13484 24124 13512
rect 23900 13472 23906 13484
rect 24118 13472 24124 13484
rect 24176 13472 24182 13524
rect 24210 13472 24216 13524
rect 24268 13512 24274 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 24268 13484 24777 13512
rect 24268 13472 24274 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 24765 13475 24823 13481
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 14458 13444 14464 13456
rect 13596 13416 14464 13444
rect 13596 13404 13602 13416
rect 14458 13404 14464 13416
rect 14516 13404 14522 13456
rect 16574 13444 16580 13456
rect 16535 13416 16580 13444
rect 16574 13404 16580 13416
rect 16632 13404 16638 13456
rect 17497 13447 17555 13453
rect 17497 13413 17509 13447
rect 17543 13444 17555 13447
rect 17586 13444 17592 13456
rect 17543 13416 17592 13444
rect 17543 13413 17555 13416
rect 17497 13407 17555 13413
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14001 13379 14059 13385
rect 14001 13376 14013 13379
rect 13964 13348 14013 13376
rect 13964 13336 13970 13348
rect 14001 13345 14013 13348
rect 14047 13376 14059 13379
rect 14182 13376 14188 13388
rect 14047 13348 14188 13376
rect 14047 13345 14059 13348
rect 14001 13339 14059 13345
rect 14182 13336 14188 13348
rect 14240 13336 14246 13388
rect 15838 13376 15844 13388
rect 15799 13348 15844 13376
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 20070 13376 20076 13388
rect 19720 13348 20076 13376
rect 14274 13308 14280 13320
rect 14235 13280 14280 13308
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 14844 13280 15945 13308
rect 14844 13240 14872 13280
rect 15933 13277 15945 13280
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 16022 13268 16028 13320
rect 16080 13308 16086 13320
rect 17681 13311 17739 13317
rect 16080 13280 16125 13308
rect 16080 13268 16086 13280
rect 17681 13277 17693 13311
rect 17727 13308 17739 13311
rect 17770 13308 17776 13320
rect 17727 13280 17776 13308
rect 17727 13277 17739 13280
rect 17681 13271 17739 13277
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 18874 13268 18880 13320
rect 18932 13308 18938 13320
rect 19720 13317 19748 13348
rect 20070 13336 20076 13348
rect 20128 13336 20134 13388
rect 21082 13336 21088 13388
rect 21140 13376 21146 13388
rect 21269 13379 21327 13385
rect 21269 13376 21281 13379
rect 21140 13348 21281 13376
rect 21140 13336 21146 13348
rect 21269 13345 21281 13348
rect 21315 13345 21327 13379
rect 24578 13376 24584 13388
rect 24539 13348 24584 13376
rect 21269 13339 21327 13345
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 18932 13280 19717 13308
rect 18932 13268 18938 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 21358 13308 21364 13320
rect 19852 13280 19897 13308
rect 21319 13280 21364 13308
rect 19852 13268 19858 13280
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21453 13311 21511 13317
rect 21453 13277 21465 13311
rect 21499 13277 21511 13311
rect 23290 13308 23296 13320
rect 23251 13280 23296 13308
rect 21453 13271 21511 13277
rect 14292 13212 14872 13240
rect 15105 13243 15163 13249
rect 14292 13184 14320 13212
rect 15105 13209 15117 13243
rect 15151 13240 15163 13243
rect 16666 13240 16672 13252
rect 15151 13212 16672 13240
rect 15151 13209 15163 13212
rect 15105 13203 15163 13209
rect 16666 13200 16672 13212
rect 16724 13240 16730 13252
rect 17037 13243 17095 13249
rect 17037 13240 17049 13243
rect 16724 13212 17049 13240
rect 16724 13200 16730 13212
rect 17037 13209 17049 13212
rect 17083 13209 17095 13243
rect 17037 13203 17095 13209
rect 18785 13243 18843 13249
rect 18785 13209 18797 13243
rect 18831 13240 18843 13243
rect 19245 13243 19303 13249
rect 19245 13240 19257 13243
rect 18831 13212 19257 13240
rect 18831 13209 18843 13212
rect 18785 13203 18843 13209
rect 19245 13209 19257 13212
rect 19291 13240 19303 13243
rect 19518 13240 19524 13252
rect 19291 13212 19524 13240
rect 19291 13209 19303 13212
rect 19245 13203 19303 13209
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 20990 13200 20996 13252
rect 21048 13240 21054 13252
rect 21468 13240 21496 13271
rect 23290 13268 23296 13280
rect 23348 13268 23354 13320
rect 21542 13240 21548 13252
rect 21048 13212 21548 13240
rect 21048 13200 21054 13212
rect 21542 13200 21548 13212
rect 21600 13200 21606 13252
rect 22649 13243 22707 13249
rect 22649 13209 22661 13243
rect 22695 13240 22707 13243
rect 24026 13240 24032 13252
rect 22695 13212 24032 13240
rect 22695 13209 22707 13212
rect 22649 13203 22707 13209
rect 24026 13200 24032 13212
rect 24084 13200 24090 13252
rect 13633 13175 13691 13181
rect 13633 13141 13645 13175
rect 13679 13172 13691 13175
rect 14274 13172 14280 13184
rect 13679 13144 14280 13172
rect 13679 13141 13691 13144
rect 13633 13135 13691 13141
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 14642 13172 14648 13184
rect 14516 13144 14648 13172
rect 14516 13132 14522 13144
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 20714 13172 20720 13184
rect 20675 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 20898 13172 20904 13184
rect 20859 13144 20904 13172
rect 20898 13132 20904 13144
rect 20956 13132 20962 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 14182 12968 14188 12980
rect 13127 12940 14188 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16117 12971 16175 12977
rect 16117 12968 16129 12971
rect 15896 12940 16129 12968
rect 15896 12928 15902 12940
rect 16117 12937 16129 12940
rect 16163 12968 16175 12971
rect 16206 12968 16212 12980
rect 16163 12940 16212 12968
rect 16163 12937 16175 12940
rect 16117 12931 16175 12937
rect 16206 12928 16212 12940
rect 16264 12928 16270 12980
rect 16298 12928 16304 12980
rect 16356 12968 16362 12980
rect 16853 12971 16911 12977
rect 16853 12968 16865 12971
rect 16356 12940 16865 12968
rect 16356 12928 16362 12940
rect 16853 12937 16865 12940
rect 16899 12937 16911 12971
rect 16853 12931 16911 12937
rect 18601 12971 18659 12977
rect 18601 12937 18613 12971
rect 18647 12968 18659 12971
rect 19794 12968 19800 12980
rect 18647 12940 19800 12968
rect 18647 12937 18659 12940
rect 18601 12931 18659 12937
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 20162 12968 20168 12980
rect 20123 12940 20168 12968
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20533 12971 20591 12977
rect 20533 12937 20545 12971
rect 20579 12968 20591 12971
rect 21174 12968 21180 12980
rect 20579 12940 21180 12968
rect 20579 12937 20591 12940
rect 20533 12931 20591 12937
rect 21174 12928 21180 12940
rect 21232 12968 21238 12980
rect 21358 12968 21364 12980
rect 21232 12940 21364 12968
rect 21232 12928 21238 12940
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 23014 12968 23020 12980
rect 22975 12940 23020 12968
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 24489 12971 24547 12977
rect 24489 12937 24501 12971
rect 24535 12968 24547 12971
rect 24670 12968 24676 12980
rect 24535 12940 24676 12968
rect 24535 12937 24547 12940
rect 24489 12931 24547 12937
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 11974 12860 11980 12912
rect 12032 12900 12038 12912
rect 13725 12903 13783 12909
rect 13725 12900 13737 12903
rect 12032 12872 13737 12900
rect 12032 12860 12038 12872
rect 13725 12869 13737 12872
rect 13771 12900 13783 12903
rect 13906 12900 13912 12912
rect 13771 12872 13912 12900
rect 13771 12869 13783 12872
rect 13725 12863 13783 12869
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 18233 12903 18291 12909
rect 18233 12869 18245 12903
rect 18279 12900 18291 12903
rect 18966 12900 18972 12912
rect 18279 12872 18972 12900
rect 18279 12869 18291 12872
rect 18233 12863 18291 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 20180 12900 20208 12928
rect 22373 12903 22431 12909
rect 20180 12872 22324 12900
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18874 12832 18880 12844
rect 17911 12804 18644 12832
rect 18835 12804 18880 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 14182 12764 14188 12776
rect 14143 12736 14188 12764
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 14458 12773 14464 12776
rect 14452 12764 14464 12773
rect 14419 12736 14464 12764
rect 14452 12727 14464 12736
rect 14458 12724 14464 12727
rect 14516 12724 14522 12776
rect 16666 12764 16672 12776
rect 16627 12736 16672 12764
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 17770 12764 17776 12776
rect 17267 12736 17776 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 18046 12764 18052 12776
rect 18007 12736 18052 12764
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18616 12764 18644 12804
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 19392 12804 19625 12832
rect 19392 12792 19398 12804
rect 19613 12801 19625 12804
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 21269 12835 21327 12841
rect 21269 12801 21281 12835
rect 21315 12832 21327 12835
rect 21726 12832 21732 12844
rect 21315 12804 21732 12832
rect 21315 12801 21327 12804
rect 21269 12795 21327 12801
rect 21726 12792 21732 12804
rect 21784 12792 21790 12844
rect 22296 12832 22324 12872
rect 22373 12869 22385 12903
rect 22419 12900 22431 12903
rect 23474 12900 23480 12912
rect 22419 12872 23480 12900
rect 22419 12869 22431 12872
rect 22373 12863 22431 12869
rect 23474 12860 23480 12872
rect 23532 12860 23538 12912
rect 22462 12832 22468 12844
rect 22296 12804 22468 12832
rect 22462 12792 22468 12804
rect 22520 12792 22526 12844
rect 22741 12835 22799 12841
rect 22741 12801 22753 12835
rect 22787 12832 22799 12835
rect 23106 12832 23112 12844
rect 22787 12804 23112 12832
rect 22787 12801 22799 12804
rect 22741 12795 22799 12801
rect 23106 12792 23112 12804
rect 23164 12792 23170 12844
rect 19518 12764 19524 12776
rect 18616 12736 19380 12764
rect 19479 12736 19524 12764
rect 13906 12656 13912 12708
rect 13964 12696 13970 12708
rect 14093 12699 14151 12705
rect 14093 12696 14105 12699
rect 13964 12668 14105 12696
rect 13964 12656 13970 12668
rect 14093 12665 14105 12668
rect 14139 12696 14151 12699
rect 14826 12696 14832 12708
rect 14139 12668 14832 12696
rect 14139 12665 14151 12668
rect 14093 12659 14151 12665
rect 14826 12656 14832 12668
rect 14884 12656 14890 12708
rect 18322 12696 18328 12708
rect 16592 12668 18328 12696
rect 16592 12640 16620 12668
rect 18322 12656 18328 12668
rect 18380 12656 18386 12708
rect 19352 12696 19380 12736
rect 19518 12724 19524 12736
rect 19576 12724 19582 12776
rect 20714 12724 20720 12776
rect 20772 12764 20778 12776
rect 20772 12736 21036 12764
rect 20772 12724 20778 12736
rect 19429 12699 19487 12705
rect 19429 12696 19441 12699
rect 19352 12668 19441 12696
rect 19429 12665 19441 12668
rect 19475 12696 19487 12699
rect 20898 12696 20904 12708
rect 19475 12668 20904 12696
rect 19475 12665 19487 12668
rect 19429 12659 19487 12665
rect 20898 12656 20904 12668
rect 20956 12656 20962 12708
rect 21008 12640 21036 12736
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 21637 12767 21695 12773
rect 21637 12764 21649 12767
rect 21140 12736 21649 12764
rect 21140 12724 21146 12736
rect 21637 12733 21649 12736
rect 21683 12733 21695 12767
rect 22186 12764 22192 12776
rect 22147 12736 22192 12764
rect 21637 12727 21695 12733
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 23750 12724 23756 12776
rect 23808 12764 23814 12776
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 23808 12736 24593 12764
rect 23808 12724 23814 12736
rect 24581 12733 24593 12736
rect 24627 12764 24639 12767
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 24627 12736 25145 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 13170 12628 13176 12640
rect 13131 12600 13176 12628
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 15565 12631 15623 12637
rect 15565 12628 15577 12631
rect 15528 12600 15577 12628
rect 15528 12588 15534 12600
rect 15565 12597 15577 12600
rect 15611 12597 15623 12631
rect 16574 12628 16580 12640
rect 16535 12600 16580 12628
rect 15565 12591 15623 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 19061 12631 19119 12637
rect 19061 12597 19073 12631
rect 19107 12628 19119 12631
rect 19150 12628 19156 12640
rect 19107 12600 19156 12628
rect 19107 12597 19119 12600
rect 19061 12591 19119 12597
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 20625 12631 20683 12637
rect 20625 12628 20637 12631
rect 20588 12600 20637 12628
rect 20588 12588 20594 12600
rect 20625 12597 20637 12600
rect 20671 12597 20683 12631
rect 20990 12628 20996 12640
rect 20951 12600 20996 12628
rect 20625 12591 20683 12597
rect 20990 12588 20996 12600
rect 21048 12588 21054 12640
rect 21085 12631 21143 12637
rect 21085 12597 21097 12631
rect 21131 12628 21143 12631
rect 21266 12628 21272 12640
rect 21131 12600 21272 12628
rect 21131 12597 21143 12600
rect 21085 12591 21143 12597
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 21542 12588 21548 12640
rect 21600 12628 21606 12640
rect 22097 12631 22155 12637
rect 22097 12628 22109 12631
rect 21600 12600 22109 12628
rect 21600 12588 21606 12600
rect 22097 12597 22109 12600
rect 22143 12628 22155 12631
rect 23198 12628 23204 12640
rect 22143 12600 23204 12628
rect 22143 12597 22155 12600
rect 22097 12591 22155 12597
rect 23198 12588 23204 12600
rect 23256 12588 23262 12640
rect 23290 12588 23296 12640
rect 23348 12628 23354 12640
rect 23477 12631 23535 12637
rect 23477 12628 23489 12631
rect 23348 12600 23489 12628
rect 23348 12588 23354 12600
rect 23477 12597 23489 12600
rect 23523 12628 23535 12631
rect 24026 12628 24032 12640
rect 23523 12600 24032 12628
rect 23523 12597 23535 12600
rect 23477 12591 23535 12597
rect 24026 12588 24032 12600
rect 24084 12588 24090 12640
rect 24762 12628 24768 12640
rect 24723 12600 24768 12628
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 12437 12427 12495 12433
rect 12437 12424 12449 12427
rect 12216 12396 12449 12424
rect 12216 12384 12222 12396
rect 12437 12393 12449 12396
rect 12483 12424 12495 12427
rect 13170 12424 13176 12436
rect 12483 12396 13176 12424
rect 12483 12393 12495 12396
rect 12437 12387 12495 12393
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 13633 12427 13691 12433
rect 13633 12393 13645 12427
rect 13679 12424 13691 12427
rect 13722 12424 13728 12436
rect 13679 12396 13728 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 15013 12427 15071 12433
rect 15013 12424 15025 12427
rect 14332 12396 15025 12424
rect 14332 12384 14338 12396
rect 15013 12393 15025 12396
rect 15059 12393 15071 12427
rect 17034 12424 17040 12436
rect 16995 12396 17040 12424
rect 15013 12387 15071 12393
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 19153 12427 19211 12433
rect 19153 12393 19165 12427
rect 19199 12424 19211 12427
rect 19242 12424 19248 12436
rect 19199 12396 19248 12424
rect 19199 12393 19211 12396
rect 19153 12387 19211 12393
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 20806 12424 20812 12436
rect 20763 12396 20812 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 20806 12384 20812 12396
rect 20864 12424 20870 12436
rect 21266 12424 21272 12436
rect 20864 12396 21272 12424
rect 20864 12384 20870 12396
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 23750 12424 23756 12436
rect 23711 12396 23756 12424
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 24210 12384 24216 12436
rect 24268 12424 24274 12436
rect 24946 12424 24952 12436
rect 24268 12396 24952 12424
rect 24268 12384 24274 12396
rect 24946 12384 24952 12396
rect 25004 12384 25010 12436
rect 11422 12316 11428 12368
rect 11480 12356 11486 12368
rect 12529 12359 12587 12365
rect 12529 12356 12541 12359
rect 11480 12328 12541 12356
rect 11480 12316 11486 12328
rect 12529 12325 12541 12328
rect 12575 12356 12587 12359
rect 13906 12356 13912 12368
rect 12575 12328 13912 12356
rect 12575 12325 12587 12328
rect 12529 12319 12587 12325
rect 13906 12316 13912 12328
rect 13964 12316 13970 12368
rect 18138 12356 18144 12368
rect 18099 12328 18144 12356
rect 18138 12316 18144 12328
rect 18196 12316 18202 12368
rect 20349 12359 20407 12365
rect 20349 12325 20361 12359
rect 20395 12356 20407 12359
rect 21352 12359 21410 12365
rect 21352 12356 21364 12359
rect 20395 12328 21364 12356
rect 20395 12325 20407 12328
rect 20349 12319 20407 12325
rect 21352 12325 21364 12328
rect 21398 12356 21410 12359
rect 21726 12356 21732 12368
rect 21398 12328 21732 12356
rect 21398 12325 21410 12328
rect 21352 12319 21410 12325
rect 21726 12316 21732 12328
rect 21784 12316 21790 12368
rect 23474 12316 23480 12368
rect 23532 12356 23538 12368
rect 23532 12328 24624 12356
rect 23532 12316 23538 12328
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 12066 12288 12072 12300
rect 11756 12260 12072 12288
rect 11756 12248 11762 12260
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 13173 12291 13231 12297
rect 13173 12257 13185 12291
rect 13219 12288 13231 12291
rect 14001 12291 14059 12297
rect 14001 12288 14013 12291
rect 13219 12260 14013 12288
rect 13219 12257 13231 12260
rect 13173 12251 13231 12257
rect 14001 12257 14013 12260
rect 14047 12257 14059 12291
rect 15913 12291 15971 12297
rect 15913 12288 15925 12291
rect 14001 12251 14059 12257
rect 15488 12260 15925 12288
rect 12713 12223 12771 12229
rect 12713 12189 12725 12223
rect 12759 12220 12771 12223
rect 12802 12220 12808 12232
rect 12759 12192 12808 12220
rect 12759 12189 12771 12192
rect 12713 12183 12771 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 12069 12155 12127 12161
rect 12069 12121 12081 12155
rect 12115 12152 12127 12155
rect 13188 12152 13216 12251
rect 15488 12232 15516 12260
rect 15913 12257 15925 12260
rect 15959 12288 15971 12291
rect 17126 12288 17132 12300
rect 15959 12260 17132 12288
rect 15959 12257 15971 12260
rect 15913 12251 15971 12257
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 19518 12248 19524 12300
rect 19576 12288 19582 12300
rect 19613 12291 19671 12297
rect 19613 12288 19625 12291
rect 19576 12260 19625 12288
rect 19576 12248 19582 12260
rect 19613 12257 19625 12260
rect 19659 12288 19671 12291
rect 20530 12288 20536 12300
rect 19659 12260 20536 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 20530 12248 20536 12260
rect 20588 12248 20594 12300
rect 23566 12288 23572 12300
rect 23527 12260 23572 12288
rect 23566 12248 23572 12260
rect 23624 12288 23630 12300
rect 24596 12297 24624 12328
rect 24397 12291 24455 12297
rect 24397 12288 24409 12291
rect 23624 12260 24409 12288
rect 23624 12248 23630 12260
rect 24397 12257 24409 12260
rect 24443 12257 24455 12291
rect 24397 12251 24455 12257
rect 24581 12291 24639 12297
rect 24581 12257 24593 12291
rect 24627 12288 24639 12291
rect 24670 12288 24676 12300
rect 24627 12260 24676 12288
rect 24627 12257 24639 12260
rect 24581 12251 24639 12257
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 13630 12220 13636 12232
rect 13587 12192 13636 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13630 12180 13636 12192
rect 13688 12220 13694 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13688 12192 14105 12220
rect 13688 12180 13694 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14274 12220 14280 12232
rect 14235 12192 14280 12220
rect 14093 12183 14151 12189
rect 14274 12180 14280 12192
rect 14332 12220 14338 12232
rect 15470 12220 15476 12232
rect 14332 12192 15476 12220
rect 14332 12180 14338 12192
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 15654 12180 15660 12232
rect 15712 12229 15718 12232
rect 15712 12220 15722 12229
rect 15712 12192 15757 12220
rect 15712 12183 15722 12192
rect 15712 12180 15718 12183
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 19484 12192 19717 12220
rect 19484 12180 19490 12192
rect 19705 12189 19717 12192
rect 19751 12189 19763 12223
rect 19705 12183 19763 12189
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12220 19947 12223
rect 20070 12220 20076 12232
rect 19935 12192 20076 12220
rect 19935 12189 19947 12192
rect 19889 12183 19947 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 21085 12223 21143 12229
rect 21085 12220 21097 12223
rect 20772 12192 21097 12220
rect 20772 12180 20778 12192
rect 21085 12189 21097 12192
rect 21131 12189 21143 12223
rect 21085 12183 21143 12189
rect 18046 12152 18052 12164
rect 12115 12124 13216 12152
rect 17959 12124 18052 12152
rect 12115 12121 12127 12124
rect 12069 12115 12127 12121
rect 18046 12112 18052 12124
rect 18104 12152 18110 12164
rect 19245 12155 19303 12161
rect 19245 12152 19257 12155
rect 18104 12124 19257 12152
rect 18104 12112 18110 12124
rect 19245 12121 19257 12124
rect 19291 12121 19303 12155
rect 19245 12115 19303 12121
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 14182 12084 14188 12096
rect 13596 12056 14188 12084
rect 13596 12044 13602 12056
rect 14182 12044 14188 12056
rect 14240 12084 14246 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14240 12056 14657 12084
rect 14240 12044 14246 12056
rect 14645 12053 14657 12056
rect 14691 12084 14703 12087
rect 15286 12084 15292 12096
rect 14691 12056 15292 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15470 12084 15476 12096
rect 15431 12056 15476 12084
rect 15470 12044 15476 12056
rect 15528 12084 15534 12096
rect 16022 12084 16028 12096
rect 15528 12056 16028 12084
rect 15528 12044 15534 12056
rect 16022 12044 16028 12056
rect 16080 12044 16086 12096
rect 17586 12084 17592 12096
rect 17547 12056 17592 12084
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 17678 12044 17684 12096
rect 17736 12084 17742 12096
rect 17862 12084 17868 12096
rect 17736 12056 17868 12084
rect 17736 12044 17742 12056
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 18288 12056 18613 12084
rect 18288 12044 18294 12056
rect 18601 12053 18613 12056
rect 18647 12053 18659 12087
rect 18601 12047 18659 12053
rect 21358 12044 21364 12096
rect 21416 12084 21422 12096
rect 22094 12084 22100 12096
rect 21416 12056 22100 12084
rect 21416 12044 21422 12056
rect 22094 12044 22100 12056
rect 22152 12044 22158 12096
rect 22465 12087 22523 12093
rect 22465 12053 22477 12087
rect 22511 12084 22523 12087
rect 22830 12084 22836 12096
rect 22511 12056 22836 12084
rect 22511 12053 22523 12056
rect 22465 12047 22523 12053
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 24118 12084 24124 12096
rect 24079 12056 24124 12084
rect 24118 12044 24124 12056
rect 24176 12044 24182 12096
rect 24762 12084 24768 12096
rect 24723 12056 24768 12084
rect 24762 12044 24768 12056
rect 24820 12044 24826 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 11422 11880 11428 11892
rect 11383 11852 11428 11880
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 13173 11883 13231 11889
rect 13173 11849 13185 11883
rect 13219 11880 13231 11883
rect 14274 11880 14280 11892
rect 13219 11852 14280 11880
rect 13219 11849 13231 11852
rect 13173 11843 13231 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 14642 11840 14648 11892
rect 14700 11880 14706 11892
rect 15013 11883 15071 11889
rect 15013 11880 15025 11883
rect 14700 11852 15025 11880
rect 14700 11840 14706 11852
rect 15013 11849 15025 11852
rect 15059 11849 15071 11883
rect 15013 11843 15071 11849
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 15654 11880 15660 11892
rect 15344 11852 15660 11880
rect 15344 11840 15350 11852
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 17126 11880 17132 11892
rect 17087 11852 17132 11880
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18966 11880 18972 11892
rect 18012 11852 18972 11880
rect 18012 11840 18018 11852
rect 18966 11840 18972 11852
rect 19024 11880 19030 11892
rect 19429 11883 19487 11889
rect 19429 11880 19441 11883
rect 19024 11852 19441 11880
rect 19024 11840 19030 11852
rect 19429 11849 19441 11852
rect 19475 11849 19487 11883
rect 19429 11843 19487 11849
rect 21726 11840 21732 11892
rect 21784 11880 21790 11892
rect 21913 11883 21971 11889
rect 21913 11880 21925 11883
rect 21784 11852 21925 11880
rect 21784 11840 21790 11852
rect 21913 11849 21925 11852
rect 21959 11849 21971 11883
rect 21913 11843 21971 11849
rect 23477 11883 23535 11889
rect 23477 11849 23489 11883
rect 23523 11880 23535 11883
rect 23658 11880 23664 11892
rect 23523 11852 23664 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 23658 11840 23664 11852
rect 23716 11840 23722 11892
rect 24670 11880 24676 11892
rect 24631 11852 24676 11880
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11744 11851 11747
rect 12802 11744 12808 11756
rect 11839 11716 12808 11744
rect 11839 11713 11851 11716
rect 11793 11707 11851 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 13538 11744 13544 11756
rect 13451 11716 13544 11744
rect 13538 11704 13544 11716
rect 13596 11744 13602 11756
rect 13633 11747 13691 11753
rect 13633 11744 13645 11747
rect 13596 11716 13645 11744
rect 13596 11704 13602 11716
rect 13633 11713 13645 11716
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 16298 11704 16304 11756
rect 16356 11744 16362 11756
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 16356 11716 16681 11744
rect 16356 11704 16362 11716
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 23676 11744 23704 11840
rect 24121 11747 24179 11753
rect 24121 11744 24133 11747
rect 23676 11716 24133 11744
rect 16669 11707 16727 11713
rect 24121 11713 24133 11716
rect 24167 11713 24179 11747
rect 24121 11707 24179 11713
rect 24213 11747 24271 11753
rect 24213 11713 24225 11747
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 16482 11676 16488 11688
rect 16443 11648 16488 11676
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 17788 11648 18061 11676
rect 12805 11611 12863 11617
rect 12805 11577 12817 11611
rect 12851 11608 12863 11611
rect 13878 11611 13936 11617
rect 13878 11608 13890 11611
rect 12851 11580 13890 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 13878 11577 13890 11580
rect 13924 11608 13936 11611
rect 14642 11608 14648 11620
rect 13924 11580 14648 11608
rect 13924 11577 13936 11580
rect 13878 11571 13936 11577
rect 14642 11568 14648 11580
rect 14700 11568 14706 11620
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 16117 11543 16175 11549
rect 16117 11540 16129 11543
rect 15804 11512 16129 11540
rect 15804 11500 15810 11512
rect 16117 11509 16129 11512
rect 16163 11509 16175 11543
rect 16117 11503 16175 11509
rect 16577 11543 16635 11549
rect 16577 11509 16589 11543
rect 16623 11540 16635 11543
rect 16666 11540 16672 11552
rect 16623 11512 16672 11540
rect 16623 11509 16635 11512
rect 16577 11503 16635 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 16942 11500 16948 11552
rect 17000 11540 17006 11552
rect 17788 11549 17816 11648
rect 18049 11645 18061 11648
rect 18095 11676 18107 11679
rect 19058 11676 19064 11688
rect 18095 11648 19064 11676
rect 18095 11645 18107 11648
rect 18049 11639 18107 11645
rect 19058 11636 19064 11648
rect 19116 11676 19122 11688
rect 20533 11679 20591 11685
rect 20533 11676 20545 11679
rect 19116 11648 20545 11676
rect 19116 11636 19122 11648
rect 20533 11645 20545 11648
rect 20579 11645 20591 11679
rect 24228 11676 24256 11707
rect 20533 11639 20591 11645
rect 24136 11648 24256 11676
rect 18230 11568 18236 11620
rect 18288 11617 18294 11620
rect 18288 11611 18352 11617
rect 18288 11577 18306 11611
rect 18340 11577 18352 11611
rect 18288 11571 18352 11577
rect 18288 11568 18294 11571
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 17000 11512 17785 11540
rect 17000 11500 17006 11512
rect 17773 11509 17785 11512
rect 17819 11509 17831 11543
rect 20070 11540 20076 11552
rect 20031 11512 20076 11540
rect 17773 11503 17831 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20441 11543 20499 11549
rect 20441 11509 20453 11543
rect 20487 11540 20499 11543
rect 20548 11540 20576 11639
rect 24136 11620 24164 11648
rect 20622 11568 20628 11620
rect 20680 11608 20686 11620
rect 20800 11611 20858 11617
rect 20800 11608 20812 11611
rect 20680 11580 20812 11608
rect 20680 11568 20686 11580
rect 20800 11577 20812 11580
rect 20846 11577 20858 11611
rect 24029 11611 24087 11617
rect 24029 11608 24041 11611
rect 20800 11571 20858 11577
rect 23032 11580 24041 11608
rect 20714 11540 20720 11552
rect 20487 11512 20720 11540
rect 20487 11509 20499 11512
rect 20441 11503 20499 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 21726 11500 21732 11552
rect 21784 11540 21790 11552
rect 22465 11543 22523 11549
rect 22465 11540 22477 11543
rect 21784 11512 22477 11540
rect 21784 11500 21790 11512
rect 22465 11509 22477 11512
rect 22511 11509 22523 11543
rect 22465 11503 22523 11509
rect 22738 11500 22744 11552
rect 22796 11540 22802 11552
rect 23032 11549 23060 11580
rect 24029 11577 24041 11580
rect 24075 11577 24087 11611
rect 24029 11571 24087 11577
rect 24118 11568 24124 11620
rect 24176 11568 24182 11620
rect 23017 11543 23075 11549
rect 23017 11540 23029 11543
rect 22796 11512 23029 11540
rect 22796 11500 22802 11512
rect 23017 11509 23029 11512
rect 23063 11509 23075 11543
rect 23017 11503 23075 11509
rect 23474 11500 23480 11552
rect 23532 11540 23538 11552
rect 23661 11543 23719 11549
rect 23661 11540 23673 11543
rect 23532 11512 23673 11540
rect 23532 11500 23538 11512
rect 23661 11509 23673 11512
rect 23707 11509 23719 11543
rect 23661 11503 23719 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 12066 11336 12072 11348
rect 12027 11308 12072 11336
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 13630 11336 13636 11348
rect 13591 11308 13636 11336
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14642 11336 14648 11348
rect 14603 11308 14648 11336
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 15105 11339 15163 11345
rect 15105 11305 15117 11339
rect 15151 11336 15163 11339
rect 15746 11336 15752 11348
rect 15151 11308 15752 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 18230 11296 18236 11348
rect 18288 11336 18294 11348
rect 18325 11339 18383 11345
rect 18325 11336 18337 11339
rect 18288 11308 18337 11336
rect 18288 11296 18294 11308
rect 18325 11305 18337 11308
rect 18371 11305 18383 11339
rect 18966 11336 18972 11348
rect 18927 11308 18972 11336
rect 18325 11299 18383 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 19797 11339 19855 11345
rect 19797 11305 19809 11339
rect 19843 11336 19855 11339
rect 20990 11336 20996 11348
rect 19843 11308 20996 11336
rect 19843 11305 19855 11308
rect 19797 11299 19855 11305
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 21450 11336 21456 11348
rect 21411 11308 21456 11336
rect 21450 11296 21456 11308
rect 21508 11296 21514 11348
rect 25222 11336 25228 11348
rect 25183 11308 25228 11336
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 14458 11228 14464 11280
rect 14516 11268 14522 11280
rect 14734 11268 14740 11280
rect 14516 11240 14740 11268
rect 14516 11228 14522 11240
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 17034 11228 17040 11280
rect 17092 11268 17098 11280
rect 17190 11271 17248 11277
rect 17190 11268 17202 11271
rect 17092 11240 17202 11268
rect 17092 11228 17098 11240
rect 17190 11237 17202 11240
rect 17236 11237 17248 11271
rect 17190 11231 17248 11237
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 13541 11203 13599 11209
rect 12492 11172 12537 11200
rect 12492 11160 12498 11172
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 14001 11203 14059 11209
rect 14001 11200 14013 11203
rect 13587 11172 14013 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 14001 11169 14013 11172
rect 14047 11200 14059 11203
rect 15286 11200 15292 11212
rect 14047 11172 15292 11200
rect 14047 11169 14059 11172
rect 14001 11163 14059 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15657 11203 15715 11209
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 16574 11200 16580 11212
rect 15703 11172 16580 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 21266 11200 21272 11212
rect 21227 11172 21272 11200
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 22548 11203 22606 11209
rect 22548 11169 22560 11203
rect 22594 11200 22606 11203
rect 22830 11200 22836 11212
rect 22594 11172 22836 11200
rect 22594 11169 22606 11172
rect 22548 11163 22606 11169
rect 22830 11160 22836 11172
rect 22888 11160 22894 11212
rect 25133 11203 25191 11209
rect 25133 11169 25145 11203
rect 25179 11200 25191 11203
rect 25590 11200 25596 11212
rect 25179 11172 25596 11200
rect 25179 11169 25191 11172
rect 25133 11163 25191 11169
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 11609 11135 11667 11141
rect 11609 11101 11621 11135
rect 11655 11132 11667 11135
rect 12526 11132 12532 11144
rect 11655 11104 12532 11132
rect 11655 11101 11667 11104
rect 11609 11095 11667 11101
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11101 12679 11135
rect 14090 11132 14096 11144
rect 14051 11104 14096 11132
rect 12621 11095 12679 11101
rect 12636 11008 12664 11095
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 14550 11132 14556 11144
rect 14323 11104 14556 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 12802 11024 12808 11076
rect 12860 11064 12866 11076
rect 13722 11064 13728 11076
rect 12860 11036 13728 11064
rect 12860 11024 12866 11036
rect 13722 11024 13728 11036
rect 13780 11064 13786 11076
rect 14292 11064 14320 11095
rect 14550 11092 14556 11104
rect 14608 11092 14614 11144
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 15436 11104 15853 11132
rect 15436 11092 15442 11104
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 16942 11132 16948 11144
rect 15841 11095 15899 11101
rect 16132 11104 16948 11132
rect 15289 11067 15347 11073
rect 15289 11064 15301 11067
rect 13780 11036 14320 11064
rect 15120 11036 15301 11064
rect 13780 11024 13786 11036
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 1581 10999 1639 11005
rect 1581 10996 1593 10999
rect 1544 10968 1593 10996
rect 1544 10956 1550 10968
rect 1581 10965 1593 10968
rect 1627 10965 1639 10999
rect 11882 10996 11888 11008
rect 11843 10968 11888 10996
rect 1581 10959 1639 10965
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 12618 10956 12624 11008
rect 12676 10956 12682 11008
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13081 10999 13139 11005
rect 13081 10996 13093 10999
rect 12952 10968 13093 10996
rect 12952 10956 12958 10968
rect 13081 10965 13093 10968
rect 13127 10965 13139 10999
rect 13081 10959 13139 10965
rect 14734 10956 14740 11008
rect 14792 10996 14798 11008
rect 15120 10996 15148 11036
rect 15289 11033 15301 11036
rect 15335 11033 15347 11067
rect 15289 11027 15347 11033
rect 15654 11024 15660 11076
rect 15712 11064 15718 11076
rect 16132 11064 16160 11104
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 20530 11092 20536 11144
rect 20588 11132 20594 11144
rect 21729 11135 21787 11141
rect 21729 11132 21741 11135
rect 20588 11104 21741 11132
rect 20588 11092 20594 11104
rect 21729 11101 21741 11104
rect 21775 11132 21787 11135
rect 22002 11132 22008 11144
rect 21775 11104 22008 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 22281 11135 22339 11141
rect 22281 11101 22293 11135
rect 22327 11101 22339 11135
rect 25406 11132 25412 11144
rect 25367 11104 25412 11132
rect 22281 11095 22339 11101
rect 16298 11064 16304 11076
rect 15712 11036 16160 11064
rect 16259 11036 16304 11064
rect 15712 11024 15718 11036
rect 16298 11024 16304 11036
rect 16356 11024 16362 11076
rect 16666 11064 16672 11076
rect 16627 11036 16672 11064
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 19426 11064 19432 11076
rect 19339 11036 19432 11064
rect 19426 11024 19432 11036
rect 19484 11064 19490 11076
rect 19484 11036 20668 11064
rect 19484 11024 19490 11036
rect 14792 10968 15148 10996
rect 14792 10956 14798 10968
rect 20162 10956 20168 11008
rect 20220 10996 20226 11008
rect 20530 10996 20536 11008
rect 20220 10968 20536 10996
rect 20220 10956 20226 10968
rect 20530 10956 20536 10968
rect 20588 10956 20594 11008
rect 20640 10996 20668 11036
rect 20714 11024 20720 11076
rect 20772 11064 20778 11076
rect 21177 11067 21235 11073
rect 21177 11064 21189 11067
rect 20772 11036 21189 11064
rect 20772 11024 20778 11036
rect 21177 11033 21189 11036
rect 21223 11064 21235 11067
rect 22186 11064 22192 11076
rect 21223 11036 22192 11064
rect 21223 11033 21235 11036
rect 21177 11027 21235 11033
rect 22186 11024 22192 11036
rect 22244 11064 22250 11076
rect 22296 11064 22324 11095
rect 25406 11092 25412 11104
rect 25464 11092 25470 11144
rect 22244 11036 22324 11064
rect 22244 11024 22250 11036
rect 23566 11024 23572 11076
rect 23624 11064 23630 11076
rect 24765 11067 24823 11073
rect 24765 11064 24777 11067
rect 23624 11036 24777 11064
rect 23624 11024 23630 11036
rect 24765 11033 24777 11036
rect 24811 11033 24823 11067
rect 24765 11027 24823 11033
rect 20898 10996 20904 11008
rect 20640 10968 20904 10996
rect 20898 10956 20904 10968
rect 20956 10956 20962 11008
rect 23661 10999 23719 11005
rect 23661 10965 23673 10999
rect 23707 10996 23719 10999
rect 23842 10996 23848 11008
rect 23707 10968 23848 10996
rect 23707 10965 23719 10968
rect 23661 10959 23719 10965
rect 23842 10956 23848 10968
rect 23900 10996 23906 11008
rect 24213 10999 24271 11005
rect 24213 10996 24225 10999
rect 23900 10968 24225 10996
rect 23900 10956 23906 10968
rect 24213 10965 24225 10968
rect 24259 10965 24271 10999
rect 24213 10959 24271 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 11517 10795 11575 10801
rect 11517 10761 11529 10795
rect 11563 10792 11575 10795
rect 11606 10792 11612 10804
rect 11563 10764 11612 10792
rect 11563 10761 11575 10764
rect 11517 10755 11575 10761
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 12618 10792 12624 10804
rect 11931 10764 12624 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 12618 10752 12624 10764
rect 12676 10792 12682 10804
rect 13630 10792 13636 10804
rect 12676 10764 13636 10792
rect 12676 10752 12682 10764
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14093 10795 14151 10801
rect 14093 10792 14105 10795
rect 13964 10764 14105 10792
rect 13964 10752 13970 10764
rect 14093 10761 14105 10764
rect 14139 10761 14151 10795
rect 14093 10755 14151 10761
rect 14458 10752 14464 10804
rect 14516 10792 14522 10804
rect 15197 10795 15255 10801
rect 15197 10792 15209 10795
rect 14516 10764 15209 10792
rect 14516 10752 14522 10764
rect 15197 10761 15209 10764
rect 15243 10792 15255 10795
rect 15381 10795 15439 10801
rect 15381 10792 15393 10795
rect 15243 10764 15393 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15381 10761 15393 10764
rect 15427 10761 15439 10795
rect 16942 10792 16948 10804
rect 16903 10764 16948 10792
rect 15381 10755 15439 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 17034 10752 17040 10804
rect 17092 10792 17098 10804
rect 17313 10795 17371 10801
rect 17313 10792 17325 10795
rect 17092 10764 17325 10792
rect 17092 10752 17098 10764
rect 17313 10761 17325 10764
rect 17359 10792 17371 10795
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 17359 10764 18245 10792
rect 17359 10761 17371 10764
rect 17313 10755 17371 10761
rect 18233 10761 18245 10764
rect 18279 10792 18291 10795
rect 18874 10792 18880 10804
rect 18279 10764 18880 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 22830 10792 22836 10804
rect 22791 10764 22836 10792
rect 22830 10752 22836 10764
rect 22888 10752 22894 10804
rect 25406 10752 25412 10804
rect 25464 10792 25470 10804
rect 25961 10795 26019 10801
rect 25961 10792 25973 10795
rect 25464 10764 25973 10792
rect 25464 10752 25470 10764
rect 25961 10761 25973 10764
rect 26007 10761 26019 10795
rect 25961 10755 26019 10761
rect 10870 10724 10876 10736
rect 10831 10696 10876 10724
rect 10870 10684 10876 10696
rect 10928 10684 10934 10736
rect 11241 10727 11299 10733
rect 11241 10693 11253 10727
rect 11287 10724 11299 10727
rect 12437 10727 12495 10733
rect 12437 10724 12449 10727
rect 11287 10696 12449 10724
rect 11287 10693 11299 10696
rect 11241 10687 11299 10693
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 9398 10656 9404 10668
rect 8260 10628 9404 10656
rect 8260 10616 8266 10628
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1486 10588 1492 10600
rect 1443 10560 1492 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1486 10548 1492 10560
rect 1544 10548 1550 10600
rect 1670 10597 1676 10600
rect 1664 10588 1676 10597
rect 1631 10560 1676 10588
rect 1664 10551 1676 10560
rect 1670 10548 1676 10551
rect 1728 10548 1734 10600
rect 11348 10597 11376 10696
rect 12437 10693 12449 10696
rect 12483 10693 12495 10727
rect 12437 10687 12495 10693
rect 14921 10727 14979 10733
rect 14921 10693 14933 10727
rect 14967 10724 14979 10727
rect 16758 10724 16764 10736
rect 14967 10696 16764 10724
rect 14967 10693 14979 10696
rect 14921 10687 14979 10693
rect 16758 10684 16764 10696
rect 16816 10684 16822 10736
rect 16960 10724 16988 10752
rect 18785 10727 18843 10733
rect 18785 10724 18797 10727
rect 16960 10696 18797 10724
rect 18785 10693 18797 10696
rect 18831 10724 18843 10727
rect 18831 10696 19012 10724
rect 18831 10693 18843 10696
rect 18785 10687 18843 10693
rect 12894 10656 12900 10668
rect 12855 10628 12900 10656
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 14642 10656 14648 10668
rect 14603 10628 14648 10656
rect 12989 10619 13047 10625
rect 11333 10591 11391 10597
rect 11333 10557 11345 10591
rect 11379 10557 11391 10591
rect 11333 10551 11391 10557
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 12618 10588 12624 10600
rect 12299 10560 12624 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 12618 10548 12624 10560
rect 12676 10588 12682 10600
rect 13004 10588 13032 10619
rect 14642 10616 14648 10628
rect 14700 10656 14706 10668
rect 16206 10656 16212 10668
rect 14700 10628 16212 10656
rect 14700 10616 14706 10628
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 18984 10665 19012 10696
rect 18969 10659 19027 10665
rect 18969 10625 18981 10659
rect 19015 10625 19027 10659
rect 22002 10656 22008 10668
rect 21963 10628 22008 10656
rect 18969 10619 19027 10625
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 12676 10560 13032 10588
rect 12676 10548 12682 10560
rect 13538 10548 13544 10600
rect 13596 10588 13602 10600
rect 13633 10591 13691 10597
rect 13633 10588 13645 10591
rect 13596 10560 13645 10588
rect 13596 10548 13602 10560
rect 13633 10557 13645 10560
rect 13679 10588 13691 10591
rect 14550 10588 14556 10600
rect 13679 10560 14556 10588
rect 13679 10557 13691 10560
rect 13633 10551 13691 10557
rect 14550 10548 14556 10560
rect 14608 10548 14614 10600
rect 15565 10591 15623 10597
rect 15565 10557 15577 10591
rect 15611 10588 15623 10591
rect 15746 10588 15752 10600
rect 15611 10560 15752 10588
rect 15611 10557 15623 10560
rect 15565 10551 15623 10557
rect 15746 10548 15752 10560
rect 15804 10588 15810 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15804 10560 16037 10588
rect 15804 10548 15810 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 19058 10548 19064 10600
rect 19116 10588 19122 10600
rect 19225 10591 19283 10597
rect 19225 10588 19237 10591
rect 19116 10560 19237 10588
rect 19116 10548 19122 10560
rect 19225 10557 19237 10560
rect 19271 10557 19283 10591
rect 19225 10551 19283 10557
rect 21361 10591 21419 10597
rect 21361 10557 21373 10591
rect 21407 10588 21419 10591
rect 21910 10588 21916 10600
rect 21407 10560 21916 10588
rect 21407 10557 21419 10560
rect 21361 10551 21419 10557
rect 21910 10548 21916 10560
rect 21968 10548 21974 10600
rect 23661 10591 23719 10597
rect 23661 10557 23673 10591
rect 23707 10557 23719 10591
rect 23661 10551 23719 10557
rect 11882 10480 11888 10532
rect 11940 10520 11946 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 11940 10492 12817 10520
rect 11940 10480 11946 10492
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 14001 10523 14059 10529
rect 14001 10520 14013 10523
rect 13964 10492 14013 10520
rect 13964 10480 13970 10492
rect 14001 10489 14013 10492
rect 14047 10520 14059 10523
rect 14461 10523 14519 10529
rect 14461 10520 14473 10523
rect 14047 10492 14473 10520
rect 14047 10489 14059 10492
rect 14001 10483 14059 10489
rect 14461 10489 14473 10492
rect 14507 10520 14519 10523
rect 14921 10523 14979 10529
rect 14921 10520 14933 10523
rect 14507 10492 14933 10520
rect 14507 10489 14519 10492
rect 14461 10483 14519 10489
rect 14921 10489 14933 10492
rect 14967 10489 14979 10523
rect 14921 10483 14979 10489
rect 15381 10523 15439 10529
rect 15381 10489 15393 10523
rect 15427 10520 15439 10523
rect 16117 10523 16175 10529
rect 16117 10520 16129 10523
rect 15427 10492 16129 10520
rect 15427 10489 15439 10492
rect 15381 10483 15439 10489
rect 16117 10489 16129 10492
rect 16163 10520 16175 10523
rect 16482 10520 16488 10532
rect 16163 10492 16488 10520
rect 16163 10489 16175 10492
rect 16117 10483 16175 10489
rect 16482 10480 16488 10492
rect 16540 10480 16546 10532
rect 20806 10480 20812 10532
rect 20864 10520 20870 10532
rect 20901 10523 20959 10529
rect 20901 10520 20913 10523
rect 20864 10492 20913 10520
rect 20864 10480 20870 10492
rect 20901 10489 20913 10492
rect 20947 10520 20959 10523
rect 21821 10523 21879 10529
rect 21821 10520 21833 10523
rect 20947 10492 21833 10520
rect 20947 10489 20959 10492
rect 20901 10483 20959 10489
rect 21821 10489 21833 10492
rect 21867 10489 21879 10523
rect 21821 10483 21879 10489
rect 23676 10464 23704 10551
rect 23842 10480 23848 10532
rect 23900 10529 23906 10532
rect 23900 10523 23964 10529
rect 23900 10489 23918 10523
rect 23952 10489 23964 10523
rect 23900 10483 23964 10489
rect 23900 10480 23906 10483
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 2832 10424 2877 10452
rect 2832 10412 2838 10424
rect 14550 10412 14556 10464
rect 14608 10452 14614 10464
rect 14608 10424 14653 10452
rect 14608 10412 14614 10424
rect 15562 10412 15568 10464
rect 15620 10452 15626 10464
rect 15657 10455 15715 10461
rect 15657 10452 15669 10455
rect 15620 10424 15669 10452
rect 15620 10412 15626 10424
rect 15657 10421 15669 10424
rect 15703 10421 15715 10455
rect 15657 10415 15715 10421
rect 20162 10412 20168 10464
rect 20220 10452 20226 10464
rect 20349 10455 20407 10461
rect 20349 10452 20361 10455
rect 20220 10424 20361 10452
rect 20220 10412 20226 10424
rect 20349 10421 20361 10424
rect 20395 10421 20407 10455
rect 20349 10415 20407 10421
rect 21453 10455 21511 10461
rect 21453 10421 21465 10455
rect 21499 10452 21511 10455
rect 21542 10452 21548 10464
rect 21499 10424 21548 10452
rect 21499 10421 21511 10424
rect 21453 10415 21511 10421
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 22186 10412 22192 10464
rect 22244 10452 22250 10464
rect 22557 10455 22615 10461
rect 22557 10452 22569 10455
rect 22244 10424 22569 10452
rect 22244 10412 22250 10424
rect 22557 10421 22569 10424
rect 22603 10452 22615 10455
rect 23385 10455 23443 10461
rect 23385 10452 23397 10455
rect 22603 10424 23397 10452
rect 22603 10421 22615 10424
rect 22557 10415 22615 10421
rect 23385 10421 23397 10424
rect 23431 10452 23443 10455
rect 23658 10452 23664 10464
rect 23431 10424 23664 10452
rect 23431 10421 23443 10424
rect 23385 10415 23443 10421
rect 23658 10412 23664 10424
rect 23716 10412 23722 10464
rect 25038 10452 25044 10464
rect 24999 10424 25044 10452
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 25590 10452 25596 10464
rect 25551 10424 25596 10452
rect 25590 10412 25596 10424
rect 25648 10412 25654 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1670 10248 1676 10260
rect 1631 10220 1676 10248
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 11057 10251 11115 10257
rect 11057 10217 11069 10251
rect 11103 10248 11115 10251
rect 11882 10248 11888 10260
rect 11103 10220 11888 10248
rect 11103 10217 11115 10220
rect 11057 10211 11115 10217
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 12621 10251 12679 10257
rect 12621 10217 12633 10251
rect 12667 10248 12679 10251
rect 12894 10248 12900 10260
rect 12667 10220 12900 10248
rect 12667 10217 12679 10220
rect 12621 10211 12679 10217
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 13722 10248 13728 10260
rect 13683 10220 13728 10248
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 14274 10208 14280 10260
rect 14332 10248 14338 10260
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 14332 10220 14381 10248
rect 14332 10208 14338 10220
rect 14369 10217 14381 10220
rect 14415 10217 14427 10251
rect 15286 10248 15292 10260
rect 15247 10220 15292 10248
rect 14369 10211 14427 10217
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 16206 10208 16212 10260
rect 16264 10248 16270 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 16264 10220 16313 10248
rect 16264 10208 16270 10220
rect 16301 10217 16313 10220
rect 16347 10217 16359 10251
rect 16301 10211 16359 10217
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 16632 10220 16681 10248
rect 16632 10208 16638 10220
rect 16669 10217 16681 10220
rect 16715 10248 16727 10251
rect 16853 10251 16911 10257
rect 16853 10248 16865 10251
rect 16715 10220 16865 10248
rect 16715 10217 16727 10220
rect 16669 10211 16727 10217
rect 16853 10217 16865 10220
rect 16899 10217 16911 10251
rect 18414 10248 18420 10260
rect 18375 10220 18420 10248
rect 16853 10211 16911 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18785 10251 18843 10257
rect 18785 10217 18797 10251
rect 18831 10248 18843 10251
rect 19242 10248 19248 10260
rect 18831 10220 19248 10248
rect 18831 10217 18843 10220
rect 18785 10211 18843 10217
rect 12161 10183 12219 10189
rect 12161 10149 12173 10183
rect 12207 10180 12219 10183
rect 12989 10183 13047 10189
rect 12989 10180 13001 10183
rect 12207 10152 13001 10180
rect 12207 10149 12219 10152
rect 12161 10143 12219 10149
rect 12989 10149 13001 10152
rect 13035 10180 13047 10183
rect 13630 10180 13636 10192
rect 13035 10152 13636 10180
rect 13035 10149 13047 10152
rect 12989 10143 13047 10149
rect 13630 10140 13636 10152
rect 13688 10140 13694 10192
rect 14090 10180 14096 10192
rect 14003 10152 14096 10180
rect 14090 10140 14096 10152
rect 14148 10180 14154 10192
rect 15562 10180 15568 10192
rect 14148 10152 15568 10180
rect 14148 10140 14154 10152
rect 15562 10140 15568 10152
rect 15620 10140 15626 10192
rect 15749 10183 15807 10189
rect 15749 10149 15761 10183
rect 15795 10180 15807 10183
rect 16114 10180 16120 10192
rect 15795 10152 16120 10180
rect 15795 10149 15807 10152
rect 15749 10143 15807 10149
rect 16114 10140 16120 10152
rect 16172 10140 16178 10192
rect 17862 10140 17868 10192
rect 17920 10180 17926 10192
rect 18800 10180 18828 10211
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 19518 10248 19524 10260
rect 19479 10220 19524 10248
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 20898 10248 20904 10260
rect 20859 10220 20904 10248
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 21266 10208 21272 10260
rect 21324 10248 21330 10260
rect 21913 10251 21971 10257
rect 21913 10248 21925 10251
rect 21324 10220 21925 10248
rect 21324 10208 21330 10220
rect 21913 10217 21925 10220
rect 21959 10248 21971 10251
rect 22278 10248 22284 10260
rect 21959 10220 22284 10248
rect 21959 10217 21971 10220
rect 21913 10211 21971 10217
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 22465 10251 22523 10257
rect 22465 10217 22477 10251
rect 22511 10248 22523 10251
rect 22738 10248 22744 10260
rect 22511 10220 22744 10248
rect 22511 10217 22523 10220
rect 22465 10211 22523 10217
rect 22738 10208 22744 10220
rect 22796 10208 22802 10260
rect 23014 10248 23020 10260
rect 22927 10220 23020 10248
rect 23014 10208 23020 10220
rect 23072 10248 23078 10260
rect 23382 10248 23388 10260
rect 23072 10220 23388 10248
rect 23072 10208 23078 10220
rect 23382 10208 23388 10220
rect 23440 10208 23446 10260
rect 25222 10208 25228 10260
rect 25280 10248 25286 10260
rect 25409 10251 25467 10257
rect 25409 10248 25421 10251
rect 25280 10220 25421 10248
rect 25280 10208 25286 10220
rect 25409 10217 25421 10220
rect 25455 10217 25467 10251
rect 25409 10211 25467 10217
rect 17920 10152 18828 10180
rect 17920 10140 17926 10152
rect 23474 10140 23480 10192
rect 23532 10180 23538 10192
rect 23722 10183 23780 10189
rect 23722 10180 23734 10183
rect 23532 10152 23734 10180
rect 23532 10140 23538 10152
rect 23722 10149 23734 10152
rect 23768 10180 23780 10183
rect 24118 10180 24124 10192
rect 23768 10152 24124 10180
rect 23768 10149 23780 10152
rect 23722 10143 23780 10149
rect 24118 10140 24124 10152
rect 24176 10180 24182 10192
rect 25038 10180 25044 10192
rect 24176 10152 25044 10180
rect 24176 10140 24182 10152
rect 25038 10140 25044 10152
rect 25096 10140 25102 10192
rect 11330 10072 11336 10124
rect 11388 10112 11394 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 11388 10084 11437 10112
rect 11388 10072 11394 10084
rect 11425 10081 11437 10084
rect 11471 10081 11483 10115
rect 11425 10075 11483 10081
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10112 13139 10115
rect 13722 10112 13728 10124
rect 13127 10084 13728 10112
rect 13127 10081 13139 10084
rect 13081 10075 13139 10081
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 14185 10115 14243 10121
rect 14185 10081 14197 10115
rect 14231 10112 14243 10115
rect 14274 10112 14280 10124
rect 14231 10084 14280 10112
rect 14231 10081 14243 10084
rect 14185 10075 14243 10081
rect 14274 10072 14280 10084
rect 14332 10112 14338 10124
rect 14734 10112 14740 10124
rect 14332 10084 14740 10112
rect 14332 10072 14338 10084
rect 14734 10072 14740 10084
rect 14792 10072 14798 10124
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 15344 10084 15669 10112
rect 15344 10072 15350 10084
rect 15657 10081 15669 10084
rect 15703 10112 15715 10115
rect 16758 10112 16764 10124
rect 15703 10084 16764 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 16758 10072 16764 10084
rect 16816 10072 16822 10124
rect 17218 10112 17224 10124
rect 17179 10084 17224 10112
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 17770 10112 17776 10124
rect 17328 10084 17776 10112
rect 10965 10047 11023 10053
rect 10965 10013 10977 10047
rect 11011 10044 11023 10047
rect 11514 10044 11520 10056
rect 11011 10016 11520 10044
rect 11011 10013 11023 10016
rect 10965 10007 11023 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11606 10004 11612 10056
rect 11664 10044 11670 10056
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11664 10016 11713 10044
rect 11664 10004 11670 10016
rect 11701 10013 11713 10016
rect 11747 10044 11759 10047
rect 13170 10044 13176 10056
rect 11747 10016 13176 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16206 10044 16212 10056
rect 15979 10016 16212 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 16942 10004 16948 10056
rect 17000 10044 17006 10056
rect 17328 10053 17356 10084
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 18877 10115 18935 10121
rect 18877 10081 18889 10115
rect 18923 10112 18935 10115
rect 19058 10112 19064 10124
rect 18923 10084 19064 10112
rect 18923 10081 18935 10084
rect 18877 10075 18935 10081
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 21269 10115 21327 10121
rect 21269 10081 21281 10115
rect 21315 10112 21327 10115
rect 21542 10112 21548 10124
rect 21315 10084 21548 10112
rect 21315 10081 21327 10084
rect 21269 10075 21327 10081
rect 21542 10072 21548 10084
rect 21600 10112 21606 10124
rect 22094 10112 22100 10124
rect 21600 10084 22100 10112
rect 21600 10072 21606 10084
rect 22094 10072 22100 10084
rect 22152 10072 22158 10124
rect 17313 10047 17371 10053
rect 17313 10044 17325 10047
rect 17000 10016 17325 10044
rect 17000 10004 17006 10016
rect 17313 10013 17325 10016
rect 17359 10013 17371 10047
rect 17313 10007 17371 10013
rect 17402 10004 17408 10056
rect 17460 10044 17466 10056
rect 18966 10044 18972 10056
rect 17460 10016 17505 10044
rect 18927 10016 18972 10044
rect 17460 10004 17466 10016
rect 18966 10004 18972 10016
rect 19024 10004 19030 10056
rect 21358 10044 21364 10056
rect 21319 10016 21364 10044
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 21453 10047 21511 10053
rect 21453 10013 21465 10047
rect 21499 10044 21511 10047
rect 21726 10044 21732 10056
rect 21499 10016 21732 10044
rect 21499 10013 21511 10016
rect 21453 10007 21511 10013
rect 21726 10004 21732 10016
rect 21784 10004 21790 10056
rect 23477 10047 23535 10053
rect 23477 10013 23489 10047
rect 23523 10013 23535 10047
rect 23477 10007 23535 10013
rect 12434 9936 12440 9988
rect 12492 9976 12498 9988
rect 15838 9976 15844 9988
rect 12492 9948 15844 9976
rect 12492 9936 12498 9948
rect 15838 9936 15844 9948
rect 15896 9936 15902 9988
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12894 9908 12900 9920
rect 12575 9880 12900 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12894 9868 12900 9880
rect 12952 9908 12958 9920
rect 13262 9908 13268 9920
rect 12952 9880 13268 9908
rect 12952 9868 12958 9880
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 14737 9911 14795 9917
rect 14737 9877 14749 9911
rect 14783 9908 14795 9911
rect 14826 9908 14832 9920
rect 14783 9880 14832 9908
rect 14783 9877 14795 9880
rect 14737 9871 14795 9877
rect 14826 9868 14832 9880
rect 14884 9908 14890 9920
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14884 9880 15025 9908
rect 14884 9868 14890 9880
rect 15013 9877 15025 9880
rect 15059 9908 15071 9911
rect 15378 9908 15384 9920
rect 15059 9880 15384 9908
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 18138 9908 18144 9920
rect 18099 9880 18144 9908
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 23492 9908 23520 10007
rect 23658 9908 23664 9920
rect 23492 9880 23664 9908
rect 23658 9868 23664 9880
rect 23716 9868 23722 9920
rect 24854 9908 24860 9920
rect 24815 9880 24860 9908
rect 24854 9868 24860 9880
rect 24912 9868 24918 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 15930 9704 15936 9716
rect 11572 9676 12296 9704
rect 11572 9664 11578 9676
rect 11241 9639 11299 9645
rect 11241 9605 11253 9639
rect 11287 9636 11299 9639
rect 11606 9636 11612 9648
rect 11287 9608 11612 9636
rect 11287 9605 11299 9608
rect 11241 9599 11299 9605
rect 11606 9596 11612 9608
rect 11664 9596 11670 9648
rect 12268 9636 12296 9676
rect 14660 9676 15936 9704
rect 12437 9639 12495 9645
rect 12437 9636 12449 9639
rect 12268 9608 12449 9636
rect 12437 9605 12449 9608
rect 12483 9605 12495 9639
rect 12437 9599 12495 9605
rect 14553 9639 14611 9645
rect 14553 9605 14565 9639
rect 14599 9636 14611 9639
rect 14660 9636 14688 9676
rect 15930 9664 15936 9676
rect 15988 9664 15994 9716
rect 16025 9707 16083 9713
rect 16025 9673 16037 9707
rect 16071 9704 16083 9707
rect 16206 9704 16212 9716
rect 16071 9676 16212 9704
rect 16071 9673 16083 9676
rect 16025 9667 16083 9673
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 16390 9704 16396 9716
rect 16316 9676 16396 9704
rect 14599 9608 14688 9636
rect 14599 9605 14611 9608
rect 14553 9599 14611 9605
rect 15746 9596 15752 9648
rect 15804 9596 15810 9648
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 10888 9540 13001 9568
rect 10134 9509 10140 9512
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9692 9472 9873 9500
rect 9692 9376 9720 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 10128 9463 10140 9509
rect 10192 9500 10198 9512
rect 10888 9500 10916 9540
rect 12989 9537 13001 9540
rect 13035 9568 13047 9571
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 13035 9540 13461 9568
rect 13035 9537 13047 9540
rect 12989 9531 13047 9537
rect 13449 9537 13461 9540
rect 13495 9568 13507 9571
rect 13630 9568 13636 9580
rect 13495 9540 13636 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 15764 9512 15792 9596
rect 16022 9528 16028 9580
rect 16080 9568 16086 9580
rect 16316 9568 16344 9676
rect 16390 9664 16396 9676
rect 16448 9664 16454 9716
rect 19889 9707 19947 9713
rect 19889 9673 19901 9707
rect 19935 9704 19947 9707
rect 20162 9704 20168 9716
rect 19935 9676 20168 9704
rect 19935 9673 19947 9676
rect 19889 9667 19947 9673
rect 20162 9664 20168 9676
rect 20220 9704 20226 9716
rect 20717 9707 20775 9713
rect 20220 9676 20392 9704
rect 20220 9664 20226 9676
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 17405 9639 17463 9645
rect 17405 9636 17417 9639
rect 16632 9608 17417 9636
rect 16632 9596 16638 9608
rect 17405 9605 17417 9608
rect 17451 9605 17463 9639
rect 17405 9599 17463 9605
rect 16080 9540 16344 9568
rect 16669 9571 16727 9577
rect 16080 9528 16086 9540
rect 16669 9537 16681 9571
rect 16715 9568 16727 9571
rect 16758 9568 16764 9580
rect 16715 9540 16764 9568
rect 16715 9537 16727 9540
rect 16669 9531 16727 9537
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 17420 9568 17448 9599
rect 17494 9596 17500 9648
rect 17552 9636 17558 9648
rect 17862 9636 17868 9648
rect 17552 9608 17868 9636
rect 17552 9596 17558 9608
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 18046 9636 18052 9648
rect 18007 9608 18052 9636
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 17678 9568 17684 9580
rect 17420 9540 17684 9568
rect 17678 9528 17684 9540
rect 17736 9568 17742 9580
rect 18230 9568 18236 9580
rect 17736 9540 18236 9568
rect 17736 9528 17742 9540
rect 18230 9528 18236 9540
rect 18288 9568 18294 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18288 9540 18521 9568
rect 18288 9528 18294 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9568 18751 9571
rect 18874 9568 18880 9580
rect 18739 9540 18880 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 18874 9528 18880 9540
rect 18932 9568 18938 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 18932 9540 19441 9568
rect 18932 9528 18938 9540
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 20364 9568 20392 9676
rect 20717 9673 20729 9707
rect 20763 9704 20775 9707
rect 21358 9704 21364 9716
rect 20763 9676 21364 9704
rect 20763 9673 20775 9676
rect 20717 9667 20775 9673
rect 21358 9664 21364 9676
rect 21416 9704 21422 9716
rect 22097 9707 22155 9713
rect 22097 9704 22109 9707
rect 21416 9676 22109 9704
rect 21416 9664 21422 9676
rect 22097 9673 22109 9676
rect 22143 9673 22155 9707
rect 22097 9667 22155 9673
rect 21726 9636 21732 9648
rect 21687 9608 21732 9636
rect 21726 9596 21732 9608
rect 21784 9596 21790 9648
rect 23658 9596 23664 9648
rect 23716 9636 23722 9648
rect 24118 9636 24124 9648
rect 23716 9608 24124 9636
rect 23716 9596 23722 9608
rect 24118 9596 24124 9608
rect 24176 9596 24182 9648
rect 21269 9571 21327 9577
rect 21269 9568 21281 9571
rect 20364 9540 21281 9568
rect 19429 9531 19487 9537
rect 21269 9537 21281 9540
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 22094 9528 22100 9580
rect 22152 9568 22158 9580
rect 22465 9571 22523 9577
rect 22465 9568 22477 9571
rect 22152 9540 22477 9568
rect 22152 9528 22158 9540
rect 22465 9537 22477 9540
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 10192 9472 10916 9500
rect 10134 9460 10140 9463
rect 10192 9460 10198 9472
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12768 9472 12817 9500
rect 12768 9460 12774 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 14645 9503 14703 9509
rect 14645 9469 14657 9503
rect 14691 9500 14703 9503
rect 14734 9500 14740 9512
rect 14691 9472 14740 9500
rect 14691 9469 14703 9472
rect 14645 9463 14703 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 15746 9460 15752 9512
rect 15804 9460 15810 9512
rect 20625 9503 20683 9509
rect 20625 9469 20637 9503
rect 20671 9500 20683 9503
rect 21082 9500 21088 9512
rect 20671 9472 21088 9500
rect 20671 9469 20683 9472
rect 20625 9463 20683 9469
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 21174 9460 21180 9512
rect 21232 9500 21238 9512
rect 24121 9503 24179 9509
rect 24121 9500 24133 9503
rect 21232 9472 21277 9500
rect 23952 9472 24133 9500
rect 21232 9460 21238 9472
rect 12728 9432 12756 9460
rect 14918 9441 14924 9444
rect 14912 9432 14924 9441
rect 12268 9404 12756 9432
rect 14879 9404 14924 9432
rect 12268 9376 12296 9404
rect 14912 9395 14924 9404
rect 14918 9392 14924 9395
rect 14976 9392 14982 9444
rect 18138 9392 18144 9444
rect 18196 9432 18202 9444
rect 18417 9435 18475 9441
rect 18417 9432 18429 9435
rect 18196 9404 18429 9432
rect 18196 9392 18202 9404
rect 18417 9401 18429 9404
rect 18463 9432 18475 9435
rect 18782 9432 18788 9444
rect 18463 9404 18788 9432
rect 18463 9401 18475 9404
rect 18417 9395 18475 9401
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 20257 9435 20315 9441
rect 20257 9401 20269 9435
rect 20303 9432 20315 9435
rect 21192 9432 21220 9460
rect 23474 9432 23480 9444
rect 20303 9404 21220 9432
rect 23032 9404 23480 9432
rect 20303 9401 20315 9404
rect 20257 9395 20315 9401
rect 9674 9364 9680 9376
rect 9635 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11388 9336 11805 9364
rect 11388 9324 11394 9336
rect 11793 9333 11805 9336
rect 11839 9333 11851 9367
rect 12250 9364 12256 9376
rect 12211 9336 12256 9364
rect 11793 9327 11851 9333
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 12894 9364 12900 9376
rect 12855 9336 12900 9364
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 13906 9364 13912 9376
rect 13780 9336 13912 9364
rect 13780 9324 13786 9336
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 16942 9364 16948 9376
rect 16816 9336 16948 9364
rect 16816 9324 16822 9336
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 18874 9324 18880 9376
rect 18932 9364 18938 9376
rect 19058 9364 19064 9376
rect 18932 9336 19064 9364
rect 18932 9324 18938 9336
rect 19058 9324 19064 9336
rect 19116 9324 19122 9376
rect 22002 9324 22008 9376
rect 22060 9364 22066 9376
rect 23032 9373 23060 9404
rect 23474 9392 23480 9404
rect 23532 9392 23538 9444
rect 23017 9367 23075 9373
rect 23017 9364 23029 9367
rect 22060 9336 23029 9364
rect 22060 9324 22066 9336
rect 23017 9333 23029 9336
rect 23063 9333 23075 9367
rect 23382 9364 23388 9376
rect 23343 9336 23388 9364
rect 23017 9327 23075 9333
rect 23382 9324 23388 9336
rect 23440 9364 23446 9376
rect 23566 9364 23572 9376
rect 23440 9336 23572 9364
rect 23440 9324 23446 9336
rect 23566 9324 23572 9336
rect 23624 9364 23630 9376
rect 23952 9373 23980 9472
rect 24121 9469 24133 9472
rect 24167 9469 24179 9503
rect 24121 9463 24179 9469
rect 24388 9503 24446 9509
rect 24388 9469 24400 9503
rect 24434 9500 24446 9503
rect 24762 9500 24768 9512
rect 24434 9472 24768 9500
rect 24434 9469 24446 9472
rect 24388 9463 24446 9469
rect 24762 9460 24768 9472
rect 24820 9460 24826 9512
rect 23937 9367 23995 9373
rect 23937 9364 23949 9367
rect 23624 9336 23949 9364
rect 23624 9324 23630 9336
rect 23937 9333 23949 9336
rect 23983 9333 23995 9367
rect 23937 9327 23995 9333
rect 24854 9324 24860 9376
rect 24912 9364 24918 9376
rect 25501 9367 25559 9373
rect 25501 9364 25513 9367
rect 24912 9336 25513 9364
rect 24912 9324 24918 9336
rect 25501 9333 25513 9336
rect 25547 9333 25559 9367
rect 25501 9327 25559 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 9953 9163 10011 9169
rect 9953 9129 9965 9163
rect 9999 9160 10011 9163
rect 10134 9160 10140 9172
rect 9999 9132 10140 9160
rect 9999 9129 10011 9132
rect 9953 9123 10011 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 12618 9160 12624 9172
rect 12579 9132 12624 9160
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 13170 9160 13176 9172
rect 13131 9132 13176 9160
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 14274 9160 14280 9172
rect 14235 9132 14280 9160
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 14918 9120 14924 9172
rect 14976 9160 14982 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 14976 9132 16681 9160
rect 14976 9120 14982 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 17770 9160 17776 9172
rect 17731 9132 17776 9160
rect 16669 9123 16727 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 18230 9160 18236 9172
rect 18191 9132 18236 9160
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 19978 9160 19984 9172
rect 19939 9132 19984 9160
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 21085 9163 21143 9169
rect 21085 9129 21097 9163
rect 21131 9160 21143 9163
rect 23109 9163 23167 9169
rect 23109 9160 23121 9163
rect 21131 9132 23121 9160
rect 21131 9129 21143 9132
rect 21085 9123 21143 9129
rect 23109 9129 23121 9132
rect 23155 9160 23167 9163
rect 23661 9163 23719 9169
rect 23661 9160 23673 9163
rect 23155 9132 23673 9160
rect 23155 9129 23167 9132
rect 23109 9123 23167 9129
rect 23661 9129 23673 9132
rect 23707 9129 23719 9163
rect 23661 9123 23719 9129
rect 23934 9120 23940 9172
rect 23992 9160 23998 9172
rect 24213 9163 24271 9169
rect 24213 9160 24225 9163
rect 23992 9132 24225 9160
rect 23992 9120 23998 9132
rect 24213 9129 24225 9132
rect 24259 9129 24271 9163
rect 24213 9123 24271 9129
rect 11146 9092 11152 9104
rect 11059 9064 11152 9092
rect 11146 9052 11152 9064
rect 11204 9092 11210 9104
rect 11508 9095 11566 9101
rect 11508 9092 11520 9095
rect 11204 9064 11520 9092
rect 11204 9052 11210 9064
rect 11508 9061 11520 9064
rect 11554 9092 11566 9095
rect 11606 9092 11612 9104
rect 11554 9064 11612 9092
rect 11554 9061 11566 9064
rect 11508 9055 11566 9061
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 15105 9095 15163 9101
rect 15105 9061 15117 9095
rect 15151 9092 15163 9095
rect 16206 9092 16212 9104
rect 15151 9064 16212 9092
rect 15151 9061 15163 9064
rect 15105 9055 15163 9061
rect 16206 9052 16212 9064
rect 16264 9052 16270 9104
rect 21453 9095 21511 9101
rect 21453 9061 21465 9095
rect 21499 9092 21511 9095
rect 21726 9092 21732 9104
rect 21499 9064 21732 9092
rect 21499 9061 21511 9064
rect 21453 9055 21511 9061
rect 21726 9052 21732 9064
rect 21784 9052 21790 9104
rect 23014 9092 23020 9104
rect 22975 9064 23020 9092
rect 23014 9052 23020 9064
rect 23072 9052 23078 9104
rect 24121 9095 24179 9101
rect 24121 9061 24133 9095
rect 24167 9092 24179 9095
rect 24762 9092 24768 9104
rect 24167 9064 24768 9092
rect 24167 9061 24179 9064
rect 24121 9055 24179 9061
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 11241 9027 11299 9033
rect 11241 9024 11253 9027
rect 9732 8996 11253 9024
rect 9732 8984 9738 8996
rect 11241 8993 11253 8996
rect 11287 9024 11299 9027
rect 11790 9024 11796 9036
rect 11287 8996 11796 9024
rect 11287 8993 11299 8996
rect 11241 8987 11299 8993
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 15556 9027 15614 9033
rect 15556 8993 15568 9027
rect 15602 9024 15614 9027
rect 16298 9024 16304 9036
rect 15602 8996 16304 9024
rect 15602 8993 15614 8996
rect 15556 8987 15614 8993
rect 16298 8984 16304 8996
rect 16356 9024 16362 9036
rect 17402 9024 17408 9036
rect 16356 8996 17408 9024
rect 16356 8984 16362 8996
rect 17402 8984 17408 8996
rect 17460 9024 17466 9036
rect 17589 9027 17647 9033
rect 17589 9024 17601 9027
rect 17460 8996 17601 9024
rect 17460 8984 17466 8996
rect 17589 8993 17601 8996
rect 17635 8993 17647 9027
rect 17589 8987 17647 8993
rect 17862 8984 17868 9036
rect 17920 9024 17926 9036
rect 18141 9027 18199 9033
rect 18141 9024 18153 9027
rect 17920 8996 18153 9024
rect 17920 8984 17926 8996
rect 18141 8993 18153 8996
rect 18187 9024 18199 9027
rect 19426 9024 19432 9036
rect 18187 8996 19432 9024
rect 18187 8993 18199 8996
rect 18141 8987 18199 8993
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14752 8928 15301 8956
rect 14752 8832 14780 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17770 8956 17776 8968
rect 17092 8928 17776 8956
rect 17092 8916 17098 8928
rect 17770 8916 17776 8928
rect 17828 8956 17834 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 17828 8928 18337 8956
rect 17828 8916 17834 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 19518 8956 19524 8968
rect 19479 8928 19524 8956
rect 18325 8919 18383 8925
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 20717 8959 20775 8965
rect 20717 8925 20729 8959
rect 20763 8956 20775 8959
rect 21082 8956 21088 8968
rect 20763 8928 21088 8956
rect 20763 8925 20775 8928
rect 20717 8919 20775 8925
rect 21082 8916 21088 8928
rect 21140 8956 21146 8968
rect 21545 8959 21603 8965
rect 21545 8956 21557 8959
rect 21140 8928 21557 8956
rect 21140 8916 21146 8928
rect 21545 8925 21557 8928
rect 21591 8925 21603 8959
rect 21545 8919 21603 8925
rect 21729 8959 21787 8965
rect 21729 8925 21741 8959
rect 21775 8956 21787 8959
rect 22002 8956 22008 8968
rect 21775 8928 22008 8956
rect 21775 8925 21787 8928
rect 21729 8919 21787 8925
rect 22002 8916 22008 8928
rect 22060 8916 22066 8968
rect 22922 8916 22928 8968
rect 22980 8956 22986 8968
rect 23293 8959 23351 8965
rect 23293 8956 23305 8959
rect 22980 8928 23305 8956
rect 22980 8916 22986 8928
rect 23293 8925 23305 8928
rect 23339 8956 23351 8959
rect 24136 8956 24164 9055
rect 24762 9052 24768 9064
rect 24820 9052 24826 9104
rect 24578 9024 24584 9036
rect 24539 8996 24584 9024
rect 24578 8984 24584 8996
rect 24636 8984 24642 9036
rect 24670 8984 24676 9036
rect 24728 9024 24734 9036
rect 25225 9027 25283 9033
rect 25225 9024 25237 9027
rect 24728 8996 25237 9024
rect 24728 8984 24734 8996
rect 25225 8993 25237 8996
rect 25271 8993 25283 9027
rect 25225 8987 25283 8993
rect 23339 8928 24164 8956
rect 24765 8959 24823 8965
rect 23339 8925 23351 8928
rect 23293 8919 23351 8925
rect 24765 8925 24777 8959
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 16574 8848 16580 8900
rect 16632 8888 16638 8900
rect 17218 8888 17224 8900
rect 16632 8860 17224 8888
rect 16632 8848 16638 8860
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 22278 8848 22284 8900
rect 22336 8888 22342 8900
rect 22649 8891 22707 8897
rect 22649 8888 22661 8891
rect 22336 8860 22661 8888
rect 22336 8848 22342 8860
rect 22649 8857 22661 8860
rect 22695 8857 22707 8891
rect 22649 8851 22707 8857
rect 24026 8848 24032 8900
rect 24084 8888 24090 8900
rect 24780 8888 24808 8919
rect 24946 8888 24952 8900
rect 24084 8860 24952 8888
rect 24084 8848 24090 8860
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 14734 8820 14740 8832
rect 14695 8792 14740 8820
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 18690 8780 18696 8832
rect 18748 8820 18754 8832
rect 18785 8823 18843 8829
rect 18785 8820 18797 8823
rect 18748 8792 18797 8820
rect 18748 8780 18754 8792
rect 18785 8789 18797 8792
rect 18831 8789 18843 8823
rect 22186 8820 22192 8832
rect 22147 8792 22192 8820
rect 18785 8783 18843 8789
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 22370 8780 22376 8832
rect 22428 8820 22434 8832
rect 22465 8823 22523 8829
rect 22465 8820 22477 8823
rect 22428 8792 22477 8820
rect 22428 8780 22434 8792
rect 22465 8789 22477 8792
rect 22511 8789 22523 8823
rect 22465 8783 22523 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 11790 8576 11796 8588
rect 11848 8616 11854 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11848 8588 12173 8616
rect 11848 8576 11854 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 17034 8616 17040 8628
rect 16995 8588 17040 8616
rect 12161 8579 12219 8585
rect 12176 8548 12204 8579
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 17497 8619 17555 8625
rect 17497 8585 17509 8619
rect 17543 8616 17555 8619
rect 17862 8616 17868 8628
rect 17543 8588 17868 8616
rect 17543 8585 17555 8588
rect 17497 8579 17555 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 18322 8616 18328 8628
rect 18095 8588 18328 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 20990 8576 20996 8628
rect 21048 8616 21054 8628
rect 21269 8619 21327 8625
rect 21269 8616 21281 8619
rect 21048 8588 21281 8616
rect 21048 8576 21054 8588
rect 21269 8585 21281 8588
rect 21315 8585 21327 8619
rect 21269 8579 21327 8585
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 22189 8619 22247 8625
rect 22189 8616 22201 8619
rect 22060 8588 22201 8616
rect 22060 8576 22066 8588
rect 22189 8585 22201 8588
rect 22235 8585 22247 8619
rect 22922 8616 22928 8628
rect 22883 8588 22928 8616
rect 22189 8579 22247 8585
rect 22922 8576 22928 8588
rect 22980 8576 22986 8628
rect 12176 8520 12480 8548
rect 11330 8480 11336 8492
rect 11291 8452 11336 8480
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 12452 8489 12480 8520
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 21821 8551 21879 8557
rect 21821 8548 21833 8551
rect 21784 8520 21833 8548
rect 21784 8508 21790 8520
rect 21821 8517 21833 8520
rect 21867 8517 21879 8551
rect 22554 8548 22560 8560
rect 22515 8520 22560 8548
rect 21821 8511 21879 8517
rect 22554 8508 22560 8520
rect 22612 8508 22618 8560
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12452 8412 12480 8443
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18690 8480 18696 8492
rect 17920 8452 18696 8480
rect 17920 8440 17926 8452
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 14734 8412 14740 8424
rect 12452 8384 14740 8412
rect 14734 8372 14740 8384
rect 14792 8412 14798 8424
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14792 8384 14933 8412
rect 14792 8372 14798 8384
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 17773 8415 17831 8421
rect 17773 8381 17785 8415
rect 17819 8412 17831 8415
rect 18138 8412 18144 8424
rect 17819 8384 18144 8412
rect 17819 8381 17831 8384
rect 17773 8375 17831 8381
rect 18138 8372 18144 8384
rect 18196 8412 18202 8424
rect 18506 8412 18512 8424
rect 18196 8384 18512 8412
rect 18196 8372 18202 8384
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 19889 8415 19947 8421
rect 19889 8381 19901 8415
rect 19935 8381 19947 8415
rect 19889 8375 19947 8381
rect 12618 8304 12624 8356
rect 12676 8353 12682 8356
rect 12676 8347 12740 8353
rect 12676 8313 12694 8347
rect 12728 8313 12740 8347
rect 14461 8347 14519 8353
rect 14461 8344 14473 8347
rect 12676 8307 12740 8313
rect 13832 8316 14473 8344
rect 12676 8304 12682 8307
rect 13832 8285 13860 8316
rect 14461 8313 14473 8316
rect 14507 8344 14519 8347
rect 15188 8347 15246 8353
rect 15188 8344 15200 8347
rect 14507 8316 15200 8344
rect 14507 8313 14519 8316
rect 14461 8307 14519 8313
rect 15188 8313 15200 8316
rect 15234 8344 15246 8347
rect 18414 8344 18420 8356
rect 15234 8316 17172 8344
rect 18375 8316 18420 8344
rect 15234 8313 15246 8316
rect 15188 8307 15246 8313
rect 13817 8279 13875 8285
rect 13817 8245 13829 8279
rect 13863 8245 13875 8279
rect 16298 8276 16304 8288
rect 16259 8248 16304 8276
rect 13817 8239 13875 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 17144 8276 17172 8316
rect 18414 8304 18420 8316
rect 18472 8344 18478 8356
rect 19061 8347 19119 8353
rect 19061 8344 19073 8347
rect 18472 8316 19073 8344
rect 18472 8304 18478 8316
rect 19061 8313 19073 8316
rect 19107 8313 19119 8347
rect 19061 8307 19119 8313
rect 17218 8276 17224 8288
rect 17144 8248 17224 8276
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 19797 8279 19855 8285
rect 19797 8245 19809 8279
rect 19843 8276 19855 8279
rect 19904 8276 19932 8375
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20145 8415 20203 8421
rect 20145 8412 20157 8415
rect 20036 8384 20157 8412
rect 20036 8372 20042 8384
rect 20145 8381 20157 8384
rect 20191 8381 20203 8415
rect 20145 8375 20203 8381
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 22373 8415 22431 8421
rect 22373 8412 22385 8415
rect 22152 8384 22385 8412
rect 22152 8372 22158 8384
rect 22373 8381 22385 8384
rect 22419 8381 22431 8415
rect 23382 8412 23388 8424
rect 23295 8384 23388 8412
rect 22373 8375 22431 8381
rect 23382 8372 23388 8384
rect 23440 8412 23446 8424
rect 24121 8415 24179 8421
rect 24121 8412 24133 8415
rect 23440 8384 24133 8412
rect 23440 8372 23446 8384
rect 24121 8381 24133 8384
rect 24167 8381 24179 8415
rect 24670 8412 24676 8424
rect 24121 8375 24179 8381
rect 24320 8384 24676 8412
rect 19978 8276 19984 8288
rect 19843 8248 19984 8276
rect 19843 8245 19855 8248
rect 19797 8239 19855 8245
rect 19978 8236 19984 8248
rect 20036 8236 20042 8288
rect 22554 8236 22560 8288
rect 22612 8276 22618 8288
rect 23400 8285 23428 8372
rect 24026 8344 24032 8356
rect 23939 8316 24032 8344
rect 24026 8304 24032 8316
rect 24084 8344 24090 8356
rect 24320 8344 24348 8384
rect 24670 8372 24676 8384
rect 24728 8372 24734 8424
rect 24394 8353 24400 8356
rect 24084 8316 24348 8344
rect 24084 8304 24090 8316
rect 24388 8307 24400 8353
rect 24452 8344 24458 8356
rect 24854 8344 24860 8356
rect 24452 8316 24860 8344
rect 24394 8304 24400 8307
rect 24452 8304 24458 8316
rect 24854 8304 24860 8316
rect 24912 8304 24918 8356
rect 23385 8279 23443 8285
rect 23385 8276 23397 8279
rect 22612 8248 23397 8276
rect 22612 8236 22618 8248
rect 23385 8245 23397 8248
rect 23431 8245 23443 8279
rect 23385 8239 23443 8245
rect 24946 8236 24952 8288
rect 25004 8276 25010 8288
rect 25501 8279 25559 8285
rect 25501 8276 25513 8279
rect 25004 8248 25513 8276
rect 25004 8236 25010 8248
rect 25501 8245 25513 8248
rect 25547 8245 25559 8279
rect 25501 8239 25559 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12676 8044 12909 8072
rect 12676 8032 12682 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 12897 8035 12955 8041
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 13909 8075 13967 8081
rect 13909 8072 13921 8075
rect 13872 8044 13921 8072
rect 13872 8032 13878 8044
rect 13909 8041 13921 8044
rect 13955 8041 13967 8075
rect 13909 8035 13967 8041
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 14921 8075 14979 8081
rect 14921 8072 14933 8075
rect 14792 8044 14933 8072
rect 14792 8032 14798 8044
rect 14921 8041 14933 8044
rect 14967 8041 14979 8075
rect 14921 8035 14979 8041
rect 15289 8075 15347 8081
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 16482 8072 16488 8084
rect 15335 8044 16488 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 16666 8072 16672 8084
rect 16623 8044 16672 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 16945 8075 17003 8081
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17034 8072 17040 8084
rect 16991 8044 17040 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 17865 8075 17923 8081
rect 17865 8072 17877 8075
rect 17736 8044 17877 8072
rect 17736 8032 17742 8044
rect 17865 8041 17877 8044
rect 17911 8041 17923 8075
rect 17865 8035 17923 8041
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18141 8075 18199 8081
rect 18141 8072 18153 8075
rect 18012 8044 18153 8072
rect 18012 8032 18018 8044
rect 18141 8041 18153 8044
rect 18187 8041 18199 8075
rect 18141 8035 18199 8041
rect 19334 8032 19340 8084
rect 19392 8072 19398 8084
rect 19429 8075 19487 8081
rect 19429 8072 19441 8075
rect 19392 8044 19441 8072
rect 19392 8032 19398 8044
rect 19429 8041 19441 8044
rect 19475 8041 19487 8075
rect 21082 8072 21088 8084
rect 21043 8044 21088 8072
rect 19429 8035 19487 8041
rect 21082 8032 21088 8044
rect 21140 8032 21146 8084
rect 24946 8072 24952 8084
rect 24907 8044 24952 8072
rect 24946 8032 24952 8044
rect 25004 8032 25010 8084
rect 15841 8007 15899 8013
rect 15841 7973 15853 8007
rect 15887 8004 15899 8007
rect 16298 8004 16304 8016
rect 15887 7976 16304 8004
rect 15887 7973 15899 7976
rect 15841 7967 15899 7973
rect 16298 7964 16304 7976
rect 16356 7964 16362 8016
rect 21545 8007 21603 8013
rect 21545 7973 21557 8007
rect 21591 8004 21603 8007
rect 21634 8004 21640 8016
rect 21591 7976 21640 8004
rect 21591 7973 21603 7976
rect 21545 7967 21603 7973
rect 21634 7964 21640 7976
rect 21692 7964 21698 8016
rect 22278 7964 22284 8016
rect 22336 8004 22342 8016
rect 24394 8004 24400 8016
rect 22336 7976 24400 8004
rect 22336 7964 22342 7976
rect 24394 7964 24400 7976
rect 24452 8004 24458 8016
rect 24581 8007 24639 8013
rect 24581 8004 24593 8007
rect 24452 7976 24593 8004
rect 24452 7964 24458 7976
rect 24581 7973 24593 7976
rect 24627 7973 24639 8007
rect 24581 7967 24639 7973
rect 12250 7936 12256 7948
rect 12211 7908 12256 7936
rect 12250 7896 12256 7908
rect 12308 7896 12314 7948
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 13906 7936 13912 7948
rect 13863 7908 13912 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 17037 7939 17095 7945
rect 17037 7905 17049 7939
rect 17083 7936 17095 7939
rect 17678 7936 17684 7948
rect 17083 7908 17684 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 18506 7936 18512 7948
rect 18467 7908 18512 7936
rect 18506 7896 18512 7908
rect 18564 7896 18570 7948
rect 21450 7936 21456 7948
rect 21411 7908 21456 7936
rect 21450 7896 21456 7908
rect 21508 7896 21514 7948
rect 22922 7945 22928 7948
rect 22916 7936 22928 7945
rect 22883 7908 22928 7936
rect 22916 7899 22928 7908
rect 22922 7896 22928 7899
rect 22980 7896 22986 7948
rect 12342 7868 12348 7880
rect 12303 7840 12348 7868
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 12710 7868 12716 7880
rect 12483 7840 12716 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 13446 7868 13452 7880
rect 12860 7840 13452 7868
rect 12860 7828 12866 7840
rect 13446 7828 13452 7840
rect 13504 7828 13510 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7868 14151 7871
rect 14182 7868 14188 7880
rect 14139 7840 14188 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 17218 7868 17224 7880
rect 17131 7840 17224 7868
rect 17218 7828 17224 7840
rect 17276 7868 17282 7880
rect 17862 7868 17868 7880
rect 17276 7840 17868 7868
rect 17276 7828 17282 7840
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 18598 7868 18604 7880
rect 18559 7840 18604 7868
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7868 19855 7871
rect 19978 7868 19984 7880
rect 19843 7840 19984 7868
rect 19843 7837 19855 7840
rect 19797 7831 19855 7837
rect 12360 7800 12388 7828
rect 12526 7800 12532 7812
rect 12360 7772 12532 7800
rect 12526 7760 12532 7772
rect 12584 7760 12590 7812
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 18708 7800 18736 7831
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 21729 7871 21787 7877
rect 21729 7868 21741 7871
rect 20763 7840 21741 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 21729 7837 21741 7840
rect 21775 7868 21787 7871
rect 21910 7868 21916 7880
rect 21775 7840 21916 7868
rect 21775 7837 21787 7840
rect 21729 7831 21787 7837
rect 21910 7828 21916 7840
rect 21968 7828 21974 7880
rect 22649 7871 22707 7877
rect 22649 7837 22661 7871
rect 22695 7837 22707 7871
rect 22649 7831 22707 7837
rect 17828 7772 18736 7800
rect 17828 7760 17834 7772
rect 19886 7760 19892 7812
rect 19944 7800 19950 7812
rect 22554 7800 22560 7812
rect 19944 7772 22560 7800
rect 19944 7760 19950 7772
rect 22554 7760 22560 7772
rect 22612 7800 22618 7812
rect 22664 7800 22692 7831
rect 22612 7772 22692 7800
rect 22612 7760 22618 7772
rect 11882 7732 11888 7744
rect 11843 7704 11888 7732
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 16482 7732 16488 7744
rect 16443 7704 16488 7732
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 22094 7692 22100 7744
rect 22152 7732 22158 7744
rect 22373 7735 22431 7741
rect 22373 7732 22385 7735
rect 22152 7704 22385 7732
rect 22152 7692 22158 7704
rect 22373 7701 22385 7704
rect 22419 7701 22431 7735
rect 22373 7695 22431 7701
rect 22646 7692 22652 7744
rect 22704 7732 22710 7744
rect 24029 7735 24087 7741
rect 24029 7732 24041 7735
rect 22704 7704 24041 7732
rect 22704 7692 22710 7704
rect 24029 7701 24041 7704
rect 24075 7701 24087 7735
rect 24029 7695 24087 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 11977 7531 12035 7537
rect 11977 7497 11989 7531
rect 12023 7528 12035 7531
rect 12250 7528 12256 7540
rect 12023 7500 12256 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 13814 7528 13820 7540
rect 12759 7500 13820 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 13814 7488 13820 7500
rect 13872 7528 13878 7540
rect 15470 7528 15476 7540
rect 13872 7500 15476 7528
rect 13872 7488 13878 7500
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 16850 7528 16856 7540
rect 15571 7500 16856 7528
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 13081 7463 13139 7469
rect 13081 7460 13093 7463
rect 13044 7432 13093 7460
rect 13044 7420 13050 7432
rect 13081 7429 13093 7432
rect 13127 7460 13139 7463
rect 13906 7460 13912 7472
rect 13127 7432 13912 7460
rect 13127 7429 13139 7432
rect 13081 7423 13139 7429
rect 13906 7420 13912 7432
rect 13964 7460 13970 7472
rect 15571 7460 15599 7500
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 17770 7528 17776 7540
rect 17731 7500 17776 7528
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 18325 7531 18383 7537
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 18506 7528 18512 7540
rect 18371 7500 18512 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 18877 7531 18935 7537
rect 18877 7528 18889 7531
rect 18656 7500 18889 7528
rect 18656 7488 18662 7500
rect 18877 7497 18889 7500
rect 18923 7497 18935 7531
rect 21450 7528 21456 7540
rect 21411 7500 21456 7528
rect 18877 7491 18935 7497
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 21726 7488 21732 7540
rect 21784 7528 21790 7540
rect 21821 7531 21879 7537
rect 21821 7528 21833 7531
rect 21784 7500 21833 7528
rect 21784 7488 21790 7500
rect 21821 7497 21833 7500
rect 21867 7528 21879 7531
rect 22646 7528 22652 7540
rect 21867 7500 22652 7528
rect 21867 7497 21879 7500
rect 21821 7491 21879 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 13964 7432 15599 7460
rect 13964 7420 13970 7432
rect 15838 7420 15844 7472
rect 15896 7460 15902 7472
rect 16393 7463 16451 7469
rect 16393 7460 16405 7463
rect 15896 7432 16405 7460
rect 15896 7420 15902 7432
rect 16393 7429 16405 7432
rect 16439 7429 16451 7463
rect 22278 7460 22284 7472
rect 16393 7423 16451 7429
rect 21744 7432 22284 7460
rect 21744 7404 21772 7432
rect 22278 7420 22284 7432
rect 22336 7420 22342 7472
rect 22370 7420 22376 7472
rect 22428 7460 22434 7472
rect 23661 7463 23719 7469
rect 23661 7460 23673 7463
rect 22428 7432 23673 7460
rect 22428 7420 22434 7432
rect 23661 7429 23673 7432
rect 23707 7429 23719 7463
rect 23661 7423 23719 7429
rect 11609 7395 11667 7401
rect 11609 7361 11621 7395
rect 11655 7392 11667 7395
rect 12710 7392 12716 7404
rect 11655 7364 12716 7392
rect 11655 7361 11667 7364
rect 11609 7355 11667 7361
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 14240 7364 14473 7392
rect 14240 7352 14246 7364
rect 14461 7361 14473 7364
rect 14507 7392 14519 7395
rect 14921 7395 14979 7401
rect 14921 7392 14933 7395
rect 14507 7364 14933 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14921 7361 14933 7364
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 16482 7352 16488 7404
rect 16540 7392 16546 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16540 7364 16865 7392
rect 16540 7352 16546 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 19337 7395 19395 7401
rect 17000 7364 17045 7392
rect 17000 7352 17006 7364
rect 19337 7361 19349 7395
rect 19383 7392 19395 7395
rect 19383 7364 19472 7392
rect 19383 7361 19395 7364
rect 19337 7355 19395 7361
rect 13449 7327 13507 7333
rect 13449 7293 13461 7327
rect 13495 7324 13507 7327
rect 14369 7327 14427 7333
rect 14369 7324 14381 7327
rect 13495 7296 14381 7324
rect 13495 7293 13507 7296
rect 13449 7287 13507 7293
rect 14369 7293 14381 7296
rect 14415 7324 14427 7327
rect 15102 7324 15108 7336
rect 14415 7296 15108 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7324 16359 7327
rect 17034 7324 17040 7336
rect 16347 7296 17040 7324
rect 16347 7293 16359 7296
rect 16301 7287 16359 7293
rect 17034 7284 17040 7296
rect 17092 7324 17098 7336
rect 18230 7324 18236 7336
rect 17092 7296 18236 7324
rect 17092 7284 17098 7296
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18598 7324 18604 7336
rect 18463 7296 18604 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 19444 7333 19472 7364
rect 21726 7352 21732 7404
rect 21784 7352 21790 7404
rect 22186 7352 22192 7404
rect 22244 7392 22250 7404
rect 22465 7395 22523 7401
rect 22465 7392 22477 7395
rect 22244 7364 22477 7392
rect 22244 7352 22250 7364
rect 22465 7361 22477 7364
rect 22511 7361 22523 7395
rect 22646 7392 22652 7404
rect 22607 7364 22652 7392
rect 22465 7355 22523 7361
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 24118 7392 24124 7404
rect 23523 7364 24124 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 19429 7327 19487 7333
rect 19429 7293 19441 7327
rect 19475 7324 19487 7327
rect 19518 7324 19524 7336
rect 19475 7296 19524 7324
rect 19475 7293 19487 7296
rect 19429 7287 19487 7293
rect 19518 7284 19524 7296
rect 19576 7324 19582 7336
rect 22370 7324 22376 7336
rect 19576 7296 19923 7324
rect 22331 7296 22376 7324
rect 19576 7284 19582 7296
rect 19895 7268 19923 7296
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 22554 7284 22560 7336
rect 22612 7324 22618 7336
rect 23017 7327 23075 7333
rect 23017 7324 23029 7327
rect 22612 7296 23029 7324
rect 22612 7284 22618 7296
rect 23017 7293 23029 7296
rect 23063 7293 23075 7327
rect 23017 7287 23075 7293
rect 14277 7259 14335 7265
rect 14277 7256 14289 7259
rect 13740 7228 14289 7256
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 13740 7197 13768 7228
rect 14277 7225 14289 7228
rect 14323 7225 14335 7259
rect 14277 7219 14335 7225
rect 15933 7259 15991 7265
rect 15933 7225 15945 7259
rect 15979 7256 15991 7259
rect 16761 7259 16819 7265
rect 16761 7256 16773 7259
rect 15979 7228 16773 7256
rect 15979 7225 15991 7228
rect 15933 7219 15991 7225
rect 16761 7225 16773 7228
rect 16807 7256 16819 7259
rect 17862 7256 17868 7268
rect 16807 7228 17868 7256
rect 16807 7225 16819 7228
rect 16761 7219 16819 7225
rect 17862 7216 17868 7228
rect 17920 7216 17926 7268
rect 19334 7216 19340 7268
rect 19392 7256 19398 7268
rect 19674 7259 19732 7265
rect 19674 7256 19686 7259
rect 19392 7228 19686 7256
rect 19392 7216 19398 7228
rect 19674 7225 19686 7228
rect 19720 7225 19732 7259
rect 19674 7219 19732 7225
rect 19886 7216 19892 7268
rect 19944 7216 19950 7268
rect 21450 7216 21456 7268
rect 21508 7256 21514 7268
rect 23492 7256 23520 7355
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 24302 7392 24308 7404
rect 24215 7364 24308 7392
rect 24302 7352 24308 7364
rect 24360 7392 24366 7404
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 24360 7364 25053 7392
rect 24360 7352 24366 7364
rect 25041 7361 25053 7364
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 21508 7228 23520 7256
rect 24029 7259 24087 7265
rect 21508 7216 21514 7228
rect 24029 7225 24041 7259
rect 24075 7256 24087 7259
rect 24765 7259 24823 7265
rect 24765 7256 24777 7259
rect 24075 7228 24777 7256
rect 24075 7225 24087 7228
rect 24029 7219 24087 7225
rect 24765 7225 24777 7228
rect 24811 7256 24823 7259
rect 25225 7259 25283 7265
rect 25225 7256 25237 7259
rect 24811 7228 25237 7256
rect 24811 7225 24823 7228
rect 24765 7219 24823 7225
rect 25225 7225 25237 7228
rect 25271 7225 25283 7259
rect 25225 7219 25283 7225
rect 13725 7191 13783 7197
rect 13725 7188 13737 7191
rect 12676 7160 13737 7188
rect 12676 7148 12682 7160
rect 13725 7157 13737 7160
rect 13771 7157 13783 7191
rect 13725 7151 13783 7157
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 13909 7191 13967 7197
rect 13909 7188 13921 7191
rect 13872 7160 13921 7188
rect 13872 7148 13878 7160
rect 13909 7157 13921 7160
rect 13955 7157 13967 7191
rect 13909 7151 13967 7157
rect 17497 7191 17555 7197
rect 17497 7157 17509 7191
rect 17543 7188 17555 7191
rect 17678 7188 17684 7200
rect 17543 7160 17684 7188
rect 17543 7157 17555 7160
rect 17497 7151 17555 7157
rect 17678 7148 17684 7160
rect 17736 7148 17742 7200
rect 18414 7148 18420 7200
rect 18472 7188 18478 7200
rect 18601 7191 18659 7197
rect 18601 7188 18613 7191
rect 18472 7160 18613 7188
rect 18472 7148 18478 7160
rect 18601 7157 18613 7160
rect 18647 7157 18659 7191
rect 20806 7188 20812 7200
rect 20767 7160 20812 7188
rect 18601 7151 18659 7157
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 22002 7188 22008 7200
rect 21963 7160 22008 7188
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 11977 6987 12035 6993
rect 11977 6953 11989 6987
rect 12023 6984 12035 6987
rect 12342 6984 12348 6996
rect 12023 6956 12348 6984
rect 12023 6953 12035 6956
rect 11977 6947 12035 6953
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 13504 6956 13645 6984
rect 13504 6944 13510 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 16945 6987 17003 6993
rect 16945 6984 16957 6987
rect 16540 6956 16957 6984
rect 16540 6944 16546 6956
rect 16945 6953 16957 6956
rect 16991 6953 17003 6987
rect 17310 6984 17316 6996
rect 17271 6956 17316 6984
rect 16945 6947 17003 6953
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 21910 6944 21916 6996
rect 21968 6984 21974 6996
rect 22186 6984 22192 6996
rect 21968 6956 22192 6984
rect 21968 6944 21974 6956
rect 22186 6944 22192 6956
rect 22244 6944 22250 6996
rect 22649 6987 22707 6993
rect 22649 6953 22661 6987
rect 22695 6984 22707 6987
rect 22922 6984 22928 6996
rect 22695 6956 22928 6984
rect 22695 6953 22707 6956
rect 22649 6947 22707 6953
rect 22922 6944 22928 6956
rect 22980 6984 22986 6996
rect 24121 6987 24179 6993
rect 24121 6984 24133 6987
rect 22980 6956 24133 6984
rect 22980 6944 22986 6956
rect 24121 6953 24133 6956
rect 24167 6984 24179 6987
rect 24302 6984 24308 6996
rect 24167 6956 24308 6984
rect 24167 6953 24179 6956
rect 24121 6947 24179 6953
rect 24302 6944 24308 6956
rect 24360 6944 24366 6996
rect 15749 6919 15807 6925
rect 15749 6916 15761 6919
rect 15120 6888 15761 6916
rect 13081 6851 13139 6857
rect 13081 6817 13093 6851
rect 13127 6848 13139 6851
rect 13538 6848 13544 6860
rect 13127 6820 13544 6848
rect 13127 6817 13139 6820
rect 13081 6811 13139 6817
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 15120 6857 15148 6888
rect 15749 6885 15761 6888
rect 15795 6916 15807 6919
rect 16390 6916 16396 6928
rect 15795 6888 16396 6916
rect 15795 6885 15807 6888
rect 15749 6879 15807 6885
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 16853 6919 16911 6925
rect 16853 6885 16865 6919
rect 16899 6916 16911 6919
rect 17218 6916 17224 6928
rect 16899 6888 17224 6916
rect 16899 6885 16911 6888
rect 16853 6879 16911 6885
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 17586 6876 17592 6928
rect 17644 6876 17650 6928
rect 21545 6919 21603 6925
rect 21545 6885 21557 6919
rect 21591 6916 21603 6919
rect 21591 6888 21956 6916
rect 21591 6885 21603 6888
rect 21545 6879 21603 6885
rect 15105 6851 15163 6857
rect 15105 6817 15117 6851
rect 15151 6817 15163 6851
rect 15105 6811 15163 6817
rect 17405 6851 17463 6857
rect 17405 6817 17417 6851
rect 17451 6848 17463 6851
rect 17604 6848 17632 6876
rect 18874 6848 18880 6860
rect 17451 6820 17632 6848
rect 18835 6820 18880 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 18874 6808 18880 6820
rect 18932 6808 18938 6860
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 20070 6848 20076 6860
rect 19843 6820 20076 6848
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 20070 6808 20076 6820
rect 20128 6808 20134 6860
rect 13630 6740 13636 6792
rect 13688 6780 13694 6792
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 13688 6752 13737 6780
rect 13688 6740 13694 6752
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 15838 6780 15844 6792
rect 15799 6752 15844 6780
rect 13725 6743 13783 6749
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6749 15991 6783
rect 15933 6743 15991 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 17635 6752 18644 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 12713 6715 12771 6721
rect 12713 6681 12725 6715
rect 12759 6712 12771 6715
rect 12759 6684 13768 6712
rect 12759 6681 12771 6684
rect 12713 6675 12771 6681
rect 13740 6656 13768 6684
rect 15562 6672 15568 6724
rect 15620 6712 15626 6724
rect 15948 6712 15976 6743
rect 15620 6684 15976 6712
rect 15620 6672 15626 6684
rect 17954 6672 17960 6724
rect 18012 6712 18018 6724
rect 18509 6715 18567 6721
rect 18509 6712 18521 6715
rect 18012 6684 18521 6712
rect 18012 6672 18018 6684
rect 18509 6681 18521 6684
rect 18555 6681 18567 6715
rect 18616 6712 18644 6752
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 18840 6752 18981 6780
rect 18840 6740 18846 6752
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19116 6752 19161 6780
rect 19116 6740 19122 6752
rect 21542 6740 21548 6792
rect 21600 6780 21606 6792
rect 21637 6783 21695 6789
rect 21637 6780 21649 6783
rect 21600 6752 21649 6780
rect 21600 6740 21606 6752
rect 21637 6749 21649 6752
rect 21683 6749 21695 6783
rect 21637 6743 21695 6749
rect 21726 6740 21732 6792
rect 21784 6780 21790 6792
rect 21928 6780 21956 6888
rect 22554 6808 22560 6860
rect 22612 6848 22618 6860
rect 23014 6857 23020 6860
rect 22741 6851 22799 6857
rect 22741 6848 22753 6851
rect 22612 6820 22753 6848
rect 22612 6808 22618 6820
rect 22741 6817 22753 6820
rect 22787 6817 22799 6851
rect 23008 6848 23020 6857
rect 22975 6820 23020 6848
rect 22741 6811 22799 6817
rect 23008 6811 23020 6820
rect 23014 6808 23020 6811
rect 23072 6808 23078 6860
rect 25222 6848 25228 6860
rect 25183 6820 25228 6848
rect 25222 6808 25228 6820
rect 25280 6808 25286 6860
rect 22002 6780 22008 6792
rect 21784 6752 21829 6780
rect 21928 6752 22008 6780
rect 21784 6740 21790 6752
rect 22002 6740 22008 6752
rect 22060 6740 22066 6792
rect 19076 6712 19104 6740
rect 21174 6712 21180 6724
rect 18616 6684 19104 6712
rect 21135 6684 21180 6712
rect 18509 6675 18567 6681
rect 21174 6672 21180 6684
rect 21232 6672 21238 6724
rect 13170 6644 13176 6656
rect 13131 6616 13176 6644
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 13722 6604 13728 6656
rect 13780 6604 13786 6656
rect 14182 6644 14188 6656
rect 14143 6616 14188 6644
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 15378 6644 15384 6656
rect 15339 6616 15384 6644
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 16482 6644 16488 6656
rect 16443 6616 16488 6644
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 18417 6647 18475 6653
rect 18417 6613 18429 6647
rect 18463 6644 18475 6647
rect 18598 6644 18604 6656
rect 18463 6616 18604 6644
rect 18463 6613 18475 6616
rect 18417 6607 18475 6613
rect 18598 6604 18604 6616
rect 18656 6604 18662 6656
rect 20717 6647 20775 6653
rect 20717 6613 20729 6647
rect 20763 6644 20775 6647
rect 21634 6644 21640 6656
rect 20763 6616 21640 6644
rect 20763 6613 20775 6616
rect 20717 6607 20775 6613
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 22186 6644 22192 6656
rect 22147 6616 22192 6644
rect 22186 6604 22192 6616
rect 22244 6604 22250 6656
rect 25406 6644 25412 6656
rect 25367 6616 25412 6644
rect 25406 6604 25412 6616
rect 25464 6604 25470 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 14734 6400 14740 6452
rect 14792 6440 14798 6452
rect 15197 6443 15255 6449
rect 15197 6440 15209 6443
rect 14792 6412 15209 6440
rect 14792 6400 14798 6412
rect 15197 6409 15209 6412
rect 15243 6440 15255 6443
rect 15289 6443 15347 6449
rect 15289 6440 15301 6443
rect 15243 6412 15301 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 15289 6409 15301 6412
rect 15335 6409 15347 6443
rect 15289 6403 15347 6409
rect 17310 6400 17316 6452
rect 17368 6440 17374 6452
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 17368 6412 17417 6440
rect 17368 6400 17374 6412
rect 17405 6409 17417 6412
rect 17451 6409 17463 6443
rect 17405 6403 17463 6409
rect 17586 6400 17592 6452
rect 17644 6440 17650 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17644 6412 17785 6440
rect 17644 6400 17650 6412
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 17773 6403 17831 6409
rect 18601 6443 18659 6449
rect 18601 6409 18613 6443
rect 18647 6440 18659 6443
rect 18874 6440 18880 6452
rect 18647 6412 18880 6440
rect 18647 6409 18659 6412
rect 18601 6403 18659 6409
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 21634 6400 21640 6452
rect 21692 6440 21698 6452
rect 21821 6443 21879 6449
rect 21821 6440 21833 6443
rect 21692 6412 21833 6440
rect 21692 6400 21698 6412
rect 21821 6409 21833 6412
rect 21867 6409 21879 6443
rect 21821 6403 21879 6409
rect 13630 6304 13636 6316
rect 13591 6276 13636 6304
rect 13630 6264 13636 6276
rect 13688 6304 13694 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13688 6276 14105 6304
rect 13688 6264 13694 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6304 14703 6307
rect 14691 6276 15608 6304
rect 14691 6273 14703 6276
rect 14645 6267 14703 6273
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6236 13599 6239
rect 13722 6236 13728 6248
rect 13587 6208 13728 6236
rect 13587 6205 13599 6208
rect 13541 6199 13599 6205
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 15197 6239 15255 6245
rect 15197 6205 15209 6239
rect 15243 6236 15255 6239
rect 15473 6239 15531 6245
rect 15473 6236 15485 6239
rect 15243 6208 15485 6236
rect 15243 6205 15255 6208
rect 15197 6199 15255 6205
rect 15473 6205 15485 6208
rect 15519 6205 15531 6239
rect 15580 6236 15608 6276
rect 15740 6239 15798 6245
rect 15740 6236 15752 6239
rect 15580 6208 15752 6236
rect 15473 6199 15531 6205
rect 15740 6205 15752 6208
rect 15786 6236 15798 6239
rect 16482 6236 16488 6248
rect 15786 6208 16488 6236
rect 15786 6205 15798 6208
rect 15740 6199 15798 6205
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 19518 6236 19524 6248
rect 19431 6208 19524 6236
rect 19518 6196 19524 6208
rect 19576 6196 19582 6248
rect 19788 6239 19846 6245
rect 19788 6205 19800 6239
rect 19834 6236 19846 6239
rect 20806 6236 20812 6248
rect 19834 6208 20812 6236
rect 19834 6205 19846 6208
rect 19788 6199 19846 6205
rect 12253 6171 12311 6177
rect 12253 6137 12265 6171
rect 12299 6168 12311 6171
rect 12526 6168 12532 6180
rect 12299 6140 12532 6168
rect 12299 6137 12311 6140
rect 12253 6131 12311 6137
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 13449 6171 13507 6177
rect 13449 6168 13461 6171
rect 12912 6140 13461 6168
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12912 6109 12940 6140
rect 13449 6137 13461 6140
rect 13495 6137 13507 6171
rect 13449 6131 13507 6137
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 14921 6171 14979 6177
rect 14921 6168 14933 6171
rect 14240 6140 14933 6168
rect 14240 6128 14246 6140
rect 14921 6137 14933 6140
rect 14967 6168 14979 6171
rect 15562 6168 15568 6180
rect 14967 6140 15568 6168
rect 14967 6137 14979 6140
rect 14921 6131 14979 6137
rect 15562 6128 15568 6140
rect 15620 6128 15626 6180
rect 16666 6128 16672 6180
rect 16724 6168 16730 6180
rect 19337 6171 19395 6177
rect 19337 6168 19349 6171
rect 16724 6140 19349 6168
rect 16724 6128 16730 6140
rect 19337 6137 19349 6140
rect 19383 6168 19395 6171
rect 19536 6168 19564 6196
rect 19383 6140 19564 6168
rect 19383 6137 19395 6140
rect 19337 6131 19395 6137
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12492 6072 12909 6100
rect 12492 6060 12498 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 13078 6100 13084 6112
rect 13039 6072 13084 6100
rect 12897 6063 12955 6069
rect 13078 6060 13084 6072
rect 13136 6060 13142 6112
rect 15580 6100 15608 6128
rect 16853 6103 16911 6109
rect 16853 6100 16865 6103
rect 15580 6072 16865 6100
rect 16853 6069 16865 6072
rect 16899 6069 16911 6103
rect 16853 6063 16911 6069
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 17920 6072 18061 6100
rect 17920 6060 17926 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 18782 6060 18788 6112
rect 18840 6100 18846 6112
rect 18877 6103 18935 6109
rect 18877 6100 18889 6103
rect 18840 6072 18889 6100
rect 18840 6060 18846 6072
rect 18877 6069 18889 6072
rect 18923 6069 18935 6103
rect 18877 6063 18935 6069
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 19803 6100 19831 6199
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 21836 6168 21864 6403
rect 21910 6400 21916 6452
rect 21968 6440 21974 6452
rect 22005 6443 22063 6449
rect 22005 6440 22017 6443
rect 21968 6412 22017 6440
rect 21968 6400 21974 6412
rect 22005 6409 22017 6412
rect 22051 6409 22063 6443
rect 22005 6403 22063 6409
rect 22554 6400 22560 6452
rect 22612 6440 22618 6452
rect 23017 6443 23075 6449
rect 23017 6440 23029 6443
rect 22612 6412 23029 6440
rect 22612 6400 22618 6412
rect 23017 6409 23029 6412
rect 23063 6409 23075 6443
rect 24026 6440 24032 6452
rect 23987 6412 24032 6440
rect 23017 6403 23075 6409
rect 24026 6400 24032 6412
rect 24084 6440 24090 6452
rect 25222 6440 25228 6452
rect 24084 6412 24716 6440
rect 25183 6412 25228 6440
rect 24084 6400 24090 6412
rect 22186 6264 22192 6316
rect 22244 6304 22250 6316
rect 22465 6307 22523 6313
rect 22465 6304 22477 6307
rect 22244 6276 22477 6304
rect 22244 6264 22250 6276
rect 22465 6273 22477 6276
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 22649 6307 22707 6313
rect 22649 6273 22661 6307
rect 22695 6304 22707 6307
rect 22922 6304 22928 6316
rect 22695 6276 22928 6304
rect 22695 6273 22707 6276
rect 22649 6267 22707 6273
rect 22922 6264 22928 6276
rect 22980 6264 22986 6316
rect 23658 6264 23664 6316
rect 23716 6304 23722 6316
rect 23934 6304 23940 6316
rect 23716 6276 23940 6304
rect 23716 6264 23722 6276
rect 23934 6264 23940 6276
rect 23992 6264 23998 6316
rect 24688 6313 24716 6412
rect 25222 6400 25228 6412
rect 25280 6400 25286 6452
rect 24673 6307 24731 6313
rect 24673 6273 24685 6307
rect 24719 6273 24731 6307
rect 24673 6267 24731 6273
rect 24857 6307 24915 6313
rect 24857 6273 24869 6307
rect 24903 6304 24915 6307
rect 25038 6304 25044 6316
rect 24903 6276 25044 6304
rect 24903 6273 24915 6276
rect 24857 6267 24915 6273
rect 25038 6264 25044 6276
rect 25096 6264 25102 6316
rect 22373 6171 22431 6177
rect 22373 6168 22385 6171
rect 21836 6140 22385 6168
rect 22373 6137 22385 6140
rect 22419 6168 22431 6171
rect 23382 6168 23388 6180
rect 22419 6140 23388 6168
rect 22419 6137 22431 6140
rect 22373 6131 22431 6137
rect 23382 6128 23388 6140
rect 23440 6128 23446 6180
rect 23477 6171 23535 6177
rect 23477 6137 23489 6171
rect 23523 6168 23535 6171
rect 24581 6171 24639 6177
rect 24581 6168 24593 6171
rect 23523 6140 24593 6168
rect 23523 6137 23535 6140
rect 23477 6131 23535 6137
rect 24581 6137 24593 6140
rect 24627 6168 24639 6171
rect 25130 6168 25136 6180
rect 24627 6140 25136 6168
rect 24627 6137 24639 6140
rect 24581 6131 24639 6137
rect 25130 6128 25136 6140
rect 25188 6128 25194 6180
rect 20898 6100 20904 6112
rect 19576 6072 19831 6100
rect 20859 6072 20904 6100
rect 19576 6060 19582 6072
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 21542 6100 21548 6112
rect 21503 6072 21548 6100
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 23566 6060 23572 6112
rect 23624 6100 23630 6112
rect 24213 6103 24271 6109
rect 24213 6100 24225 6103
rect 23624 6072 24225 6100
rect 23624 6060 23630 6072
rect 24213 6069 24225 6072
rect 24259 6069 24271 6103
rect 24213 6063 24271 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 14001 5899 14059 5905
rect 14001 5896 14013 5899
rect 13504 5868 14013 5896
rect 13504 5856 13510 5868
rect 14001 5865 14013 5868
rect 14047 5865 14059 5899
rect 14001 5859 14059 5865
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 15838 5896 15844 5908
rect 15151 5868 15844 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 19518 5896 19524 5908
rect 19479 5868 19524 5896
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 20717 5899 20775 5905
rect 20717 5865 20729 5899
rect 20763 5896 20775 5899
rect 21726 5896 21732 5908
rect 20763 5868 21732 5896
rect 20763 5865 20775 5868
rect 20717 5859 20775 5865
rect 21726 5856 21732 5868
rect 21784 5856 21790 5908
rect 22373 5899 22431 5905
rect 22373 5865 22385 5899
rect 22419 5896 22431 5899
rect 22922 5896 22928 5908
rect 22419 5868 22928 5896
rect 22419 5865 22431 5868
rect 22373 5859 22431 5865
rect 22922 5856 22928 5868
rect 22980 5856 22986 5908
rect 25130 5856 25136 5908
rect 25188 5896 25194 5908
rect 25225 5899 25283 5905
rect 25225 5896 25237 5899
rect 25188 5868 25237 5896
rect 25188 5856 25194 5868
rect 25225 5865 25237 5868
rect 25271 5865 25283 5899
rect 25225 5859 25283 5865
rect 12250 5788 12256 5840
rect 12308 5837 12314 5840
rect 12308 5831 12372 5837
rect 12308 5797 12326 5831
rect 12360 5797 12372 5831
rect 12308 5791 12372 5797
rect 12308 5788 12314 5791
rect 12434 5788 12440 5840
rect 12492 5788 12498 5840
rect 15657 5831 15715 5837
rect 15657 5797 15669 5831
rect 15703 5828 15715 5831
rect 16206 5828 16212 5840
rect 15703 5800 16212 5828
rect 15703 5797 15715 5800
rect 15657 5791 15715 5797
rect 16206 5788 16212 5800
rect 16264 5788 16270 5840
rect 16577 5831 16635 5837
rect 16577 5797 16589 5831
rect 16623 5828 16635 5831
rect 16945 5831 17003 5837
rect 16945 5828 16957 5831
rect 16623 5800 16957 5828
rect 16623 5797 16635 5800
rect 16577 5791 16635 5797
rect 16945 5797 16957 5800
rect 16991 5828 17003 5831
rect 17304 5831 17362 5837
rect 17304 5828 17316 5831
rect 16991 5800 17316 5828
rect 16991 5797 17003 5800
rect 16945 5791 17003 5797
rect 17304 5797 17316 5800
rect 17350 5828 17362 5831
rect 19058 5828 19064 5840
rect 17350 5800 19064 5828
rect 17350 5797 17362 5800
rect 17304 5791 17362 5797
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 21358 5828 21364 5840
rect 21319 5800 21364 5828
rect 21358 5788 21364 5800
rect 21416 5788 21422 5840
rect 12452 5760 12480 5788
rect 13630 5760 13636 5772
rect 12452 5732 13636 5760
rect 12066 5692 12072 5704
rect 12027 5664 12072 5692
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 13464 5633 13492 5732
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 15838 5760 15844 5772
rect 15795 5732 15844 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 19705 5763 19763 5769
rect 19705 5729 19717 5763
rect 19751 5760 19763 5763
rect 20070 5760 20076 5772
rect 19751 5732 20076 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 20070 5720 20076 5732
rect 20128 5720 20134 5772
rect 21266 5760 21272 5772
rect 21227 5732 21272 5760
rect 21266 5720 21272 5732
rect 21324 5720 21330 5772
rect 22462 5760 22468 5772
rect 22423 5732 22468 5760
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 24029 5763 24087 5769
rect 24029 5729 24041 5763
rect 24075 5760 24087 5763
rect 24854 5760 24860 5772
rect 24075 5732 24860 5760
rect 24075 5729 24087 5732
rect 24029 5723 24087 5729
rect 24854 5720 24860 5732
rect 24912 5720 24918 5772
rect 15930 5692 15936 5704
rect 15891 5664 15936 5692
rect 15930 5652 15936 5664
rect 15988 5652 15994 5704
rect 16666 5652 16672 5704
rect 16724 5692 16730 5704
rect 17037 5695 17095 5701
rect 17037 5692 17049 5695
rect 16724 5664 17049 5692
rect 16724 5652 16730 5664
rect 17037 5661 17049 5664
rect 17083 5661 17095 5695
rect 17037 5655 17095 5661
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 20864 5664 21465 5692
rect 20864 5652 20870 5664
rect 21453 5661 21465 5664
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 23474 5652 23480 5704
rect 23532 5692 23538 5704
rect 24121 5695 24179 5701
rect 24121 5692 24133 5695
rect 23532 5664 24133 5692
rect 23532 5652 23538 5664
rect 24121 5661 24133 5664
rect 24167 5661 24179 5695
rect 24121 5655 24179 5661
rect 24305 5695 24363 5701
rect 24305 5661 24317 5695
rect 24351 5692 24363 5695
rect 24351 5664 24808 5692
rect 24351 5661 24363 5664
rect 24305 5655 24363 5661
rect 13449 5627 13507 5633
rect 13449 5593 13461 5627
rect 13495 5593 13507 5627
rect 15286 5624 15292 5636
rect 15247 5596 15292 5624
rect 13449 5587 13507 5593
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 22649 5627 22707 5633
rect 22649 5593 22661 5627
rect 22695 5624 22707 5627
rect 23382 5624 23388 5636
rect 22695 5596 23388 5624
rect 22695 5593 22707 5596
rect 22649 5587 22707 5593
rect 23382 5584 23388 5596
rect 23440 5584 23446 5636
rect 23569 5627 23627 5633
rect 23569 5593 23581 5627
rect 23615 5624 23627 5627
rect 24026 5624 24032 5636
rect 23615 5596 24032 5624
rect 23615 5593 23627 5596
rect 23569 5587 23627 5593
rect 24026 5584 24032 5596
rect 24084 5624 24090 5636
rect 24320 5624 24348 5655
rect 24084 5596 24348 5624
rect 24084 5584 24090 5596
rect 11977 5559 12035 5565
rect 11977 5525 11989 5559
rect 12023 5556 12035 5559
rect 13078 5556 13084 5568
rect 12023 5528 13084 5556
rect 12023 5525 12035 5528
rect 11977 5519 12035 5525
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 17770 5516 17776 5568
rect 17828 5556 17834 5568
rect 18417 5559 18475 5565
rect 18417 5556 18429 5559
rect 17828 5528 18429 5556
rect 17828 5516 17834 5528
rect 18417 5525 18429 5528
rect 18463 5525 18475 5559
rect 18417 5519 18475 5525
rect 19889 5559 19947 5565
rect 19889 5525 19901 5559
rect 19935 5556 19947 5559
rect 20254 5556 20260 5568
rect 19935 5528 20260 5556
rect 19935 5525 19947 5528
rect 19889 5519 19947 5525
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20349 5559 20407 5565
rect 20349 5525 20361 5559
rect 20395 5556 20407 5559
rect 20438 5556 20444 5568
rect 20395 5528 20444 5556
rect 20395 5525 20407 5528
rect 20349 5519 20407 5525
rect 20438 5516 20444 5528
rect 20496 5516 20502 5568
rect 20898 5556 20904 5568
rect 20859 5528 20904 5556
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 22002 5556 22008 5568
rect 21963 5528 22008 5556
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 23106 5556 23112 5568
rect 23067 5528 23112 5556
rect 23106 5516 23112 5528
rect 23164 5516 23170 5568
rect 23290 5516 23296 5568
rect 23348 5556 23354 5568
rect 24780 5565 24808 5664
rect 23661 5559 23719 5565
rect 23661 5556 23673 5559
rect 23348 5528 23673 5556
rect 23348 5516 23354 5528
rect 23661 5525 23673 5528
rect 23707 5525 23719 5559
rect 23661 5519 23719 5525
rect 24765 5559 24823 5565
rect 24765 5525 24777 5559
rect 24811 5556 24823 5559
rect 25038 5556 25044 5568
rect 24811 5528 25044 5556
rect 24811 5525 24823 5528
rect 24765 5519 24823 5525
rect 25038 5516 25044 5528
rect 25096 5516 25102 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 12066 5352 12072 5364
rect 12027 5324 12072 5352
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 14274 5312 14280 5364
rect 14332 5352 14338 5364
rect 15473 5355 15531 5361
rect 15473 5352 15485 5355
rect 14332 5324 15485 5352
rect 14332 5312 14338 5324
rect 15120 5296 15148 5324
rect 15473 5321 15485 5324
rect 15519 5352 15531 5355
rect 15930 5352 15936 5364
rect 15519 5324 15936 5352
rect 15519 5321 15531 5324
rect 15473 5315 15531 5321
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 16117 5355 16175 5361
rect 16117 5321 16129 5355
rect 16163 5352 16175 5355
rect 16206 5352 16212 5364
rect 16163 5324 16212 5352
rect 16163 5321 16175 5324
rect 16117 5315 16175 5321
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 19889 5355 19947 5361
rect 19889 5321 19901 5355
rect 19935 5352 19947 5355
rect 20162 5352 20168 5364
rect 19935 5324 20168 5352
rect 19935 5321 19947 5324
rect 19889 5315 19947 5321
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20864 5324 21005 5352
rect 20864 5312 20870 5324
rect 20993 5321 21005 5324
rect 21039 5321 21051 5355
rect 21358 5352 21364 5364
rect 21319 5324 21364 5352
rect 20993 5315 21051 5321
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 21818 5312 21824 5364
rect 21876 5352 21882 5364
rect 22005 5355 22063 5361
rect 22005 5352 22017 5355
rect 21876 5324 22017 5352
rect 21876 5312 21882 5324
rect 22005 5321 22017 5324
rect 22051 5321 22063 5355
rect 22005 5315 22063 5321
rect 22462 5312 22468 5364
rect 22520 5352 22526 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22520 5324 23029 5352
rect 22520 5312 22526 5324
rect 23017 5321 23029 5324
rect 23063 5321 23075 5355
rect 23017 5315 23075 5321
rect 23106 5312 23112 5364
rect 23164 5352 23170 5364
rect 23164 5324 24808 5352
rect 23164 5312 23170 5324
rect 11241 5287 11299 5293
rect 11241 5253 11253 5287
rect 11287 5284 11299 5287
rect 12250 5284 12256 5296
rect 11287 5256 12256 5284
rect 11287 5253 11299 5256
rect 11241 5247 11299 5253
rect 12250 5244 12256 5256
rect 12308 5244 12314 5296
rect 15102 5244 15108 5296
rect 15160 5244 15166 5296
rect 18325 5287 18383 5293
rect 18325 5253 18337 5287
rect 18371 5284 18383 5287
rect 18874 5284 18880 5296
rect 18371 5256 18880 5284
rect 18371 5253 18383 5256
rect 18325 5247 18383 5253
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 19981 5287 20039 5293
rect 19981 5253 19993 5287
rect 20027 5284 20039 5287
rect 20714 5284 20720 5296
rect 20027 5256 20720 5284
rect 20027 5253 20039 5256
rect 19981 5247 20039 5253
rect 20714 5244 20720 5256
rect 20772 5244 20778 5296
rect 23124 5284 23152 5312
rect 22664 5256 23152 5284
rect 24780 5284 24808 5324
rect 24854 5312 24860 5364
rect 24912 5352 24918 5364
rect 25777 5355 25835 5361
rect 25777 5352 25789 5355
rect 24912 5324 25789 5352
rect 24912 5312 24918 5324
rect 25777 5321 25789 5324
rect 25823 5321 25835 5355
rect 25777 5315 25835 5321
rect 25225 5287 25283 5293
rect 25225 5284 25237 5287
rect 24780 5256 25237 5284
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 12342 5216 12348 5228
rect 11379 5188 12348 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5216 13231 5219
rect 13538 5216 13544 5228
rect 13219 5188 13544 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 16868 5188 17417 5216
rect 16868 5160 16896 5188
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 19061 5219 19119 5225
rect 19061 5185 19073 5219
rect 19107 5216 19119 5219
rect 19518 5216 19524 5228
rect 19107 5188 19524 5216
rect 19107 5185 19119 5188
rect 19061 5179 19119 5185
rect 19518 5176 19524 5188
rect 19576 5176 19582 5228
rect 20438 5176 20444 5228
rect 20496 5216 20502 5228
rect 20625 5219 20683 5225
rect 20625 5216 20637 5219
rect 20496 5188 20637 5216
rect 20496 5176 20502 5188
rect 20625 5185 20637 5188
rect 20671 5216 20683 5219
rect 20990 5216 20996 5228
rect 20671 5188 20996 5216
rect 20671 5185 20683 5188
rect 20625 5179 20683 5185
rect 20990 5176 20996 5188
rect 21048 5176 21054 5228
rect 22664 5225 22692 5256
rect 25225 5253 25237 5256
rect 25271 5253 25283 5287
rect 25225 5247 25283 5253
rect 21913 5219 21971 5225
rect 21913 5185 21925 5219
rect 21959 5216 21971 5219
rect 22649 5219 22707 5225
rect 22649 5216 22661 5219
rect 21959 5188 22661 5216
rect 21959 5185 21971 5188
rect 21913 5179 21971 5185
rect 22649 5185 22661 5188
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5216 22891 5219
rect 23566 5216 23572 5228
rect 22879 5188 23572 5216
rect 22879 5185 22891 5188
rect 22833 5179 22891 5185
rect 23566 5176 23572 5188
rect 23624 5176 23630 5228
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 13078 5148 13084 5160
rect 12943 5120 13084 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13906 5108 13912 5160
rect 13964 5148 13970 5160
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13964 5120 14013 5148
rect 13964 5108 13970 5120
rect 14001 5117 14013 5120
rect 14047 5148 14059 5151
rect 14093 5151 14151 5157
rect 14093 5148 14105 5151
rect 14047 5120 14105 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14093 5117 14105 5120
rect 14139 5148 14151 5151
rect 14734 5148 14740 5160
rect 14139 5120 14740 5148
rect 14139 5117 14151 5120
rect 14093 5111 14151 5117
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 16850 5148 16856 5160
rect 16811 5120 16856 5148
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 18877 5151 18935 5157
rect 18877 5148 18889 5151
rect 17788 5120 18889 5148
rect 11422 5040 11428 5092
rect 11480 5080 11486 5092
rect 12989 5083 13047 5089
rect 11480 5052 12940 5080
rect 11480 5040 11486 5052
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12529 5015 12587 5021
rect 12529 5012 12541 5015
rect 12400 4984 12541 5012
rect 12400 4972 12406 4984
rect 12529 4981 12541 4984
rect 12575 4981 12587 5015
rect 12912 5012 12940 5052
rect 12989 5049 13001 5083
rect 13035 5080 13047 5083
rect 13170 5080 13176 5092
rect 13035 5052 13176 5080
rect 13035 5049 13047 5052
rect 12989 5043 13047 5049
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 14182 5040 14188 5092
rect 14240 5080 14246 5092
rect 17788 5089 17816 5120
rect 18877 5117 18889 5120
rect 18923 5117 18935 5151
rect 18877 5111 18935 5117
rect 19978 5108 19984 5160
rect 20036 5148 20042 5160
rect 20349 5151 20407 5157
rect 20349 5148 20361 5151
rect 20036 5120 20361 5148
rect 20036 5108 20042 5120
rect 20349 5117 20361 5120
rect 20395 5117 20407 5151
rect 20349 5111 20407 5117
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22152 5120 22477 5148
rect 22152 5108 22158 5120
rect 22465 5117 22477 5120
rect 22511 5148 22523 5151
rect 23290 5148 23296 5160
rect 22511 5120 23296 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 23290 5108 23296 5120
rect 23348 5108 23354 5160
rect 23845 5151 23903 5157
rect 23845 5148 23857 5151
rect 23400 5120 23857 5148
rect 14338 5083 14396 5089
rect 14338 5080 14350 5083
rect 14240 5052 14350 5080
rect 14240 5040 14246 5052
rect 14338 5049 14350 5052
rect 14384 5049 14396 5083
rect 17773 5083 17831 5089
rect 17773 5080 17785 5083
rect 14338 5043 14396 5049
rect 15028 5052 17785 5080
rect 15028 5012 15056 5052
rect 17773 5049 17785 5052
rect 17819 5049 17831 5083
rect 18966 5080 18972 5092
rect 17773 5043 17831 5049
rect 18432 5052 18972 5080
rect 16666 5012 16672 5024
rect 12912 4984 15056 5012
rect 16627 4984 16672 5012
rect 12529 4975 12587 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 17034 5012 17040 5024
rect 16995 4984 17040 5012
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 18432 5021 18460 5052
rect 18966 5040 18972 5052
rect 19024 5040 19030 5092
rect 20162 5040 20168 5092
rect 20220 5080 20226 5092
rect 20441 5083 20499 5089
rect 20441 5080 20453 5083
rect 20220 5052 20453 5080
rect 20220 5040 20226 5052
rect 20441 5049 20453 5052
rect 20487 5049 20499 5083
rect 20441 5043 20499 5049
rect 22373 5083 22431 5089
rect 22373 5049 22385 5083
rect 22419 5080 22431 5083
rect 22833 5083 22891 5089
rect 22833 5080 22845 5083
rect 22419 5052 22845 5080
rect 22419 5049 22431 5052
rect 22373 5043 22431 5049
rect 22480 5024 22508 5052
rect 22833 5049 22845 5052
rect 22879 5049 22891 5083
rect 22833 5043 22891 5049
rect 18417 5015 18475 5021
rect 18417 4981 18429 5015
rect 18463 4981 18475 5015
rect 18417 4975 18475 4981
rect 18785 5015 18843 5021
rect 18785 4981 18797 5015
rect 18831 5012 18843 5015
rect 18874 5012 18880 5024
rect 18831 4984 18880 5012
rect 18831 4981 18843 4984
rect 18785 4975 18843 4981
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 19518 5012 19524 5024
rect 19479 4984 19524 5012
rect 19518 4972 19524 4984
rect 19576 4972 19582 5024
rect 22462 4972 22468 5024
rect 22520 4972 22526 5024
rect 23106 4972 23112 5024
rect 23164 5012 23170 5024
rect 23400 5021 23428 5120
rect 23845 5117 23857 5120
rect 23891 5117 23903 5151
rect 23845 5111 23903 5117
rect 24026 5040 24032 5092
rect 24084 5089 24090 5092
rect 24084 5083 24148 5089
rect 24084 5049 24102 5083
rect 24136 5049 24148 5083
rect 24084 5043 24148 5049
rect 24084 5040 24090 5043
rect 23385 5015 23443 5021
rect 23385 5012 23397 5015
rect 23164 4984 23397 5012
rect 23164 4972 23170 4984
rect 23385 4981 23397 4984
rect 23431 4981 23443 5015
rect 23385 4975 23443 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 12069 4811 12127 4817
rect 12069 4777 12081 4811
rect 12115 4808 12127 4811
rect 13170 4808 13176 4820
rect 12115 4780 13176 4808
rect 12115 4777 12127 4780
rect 12069 4771 12127 4777
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 13538 4808 13544 4820
rect 13499 4780 13544 4808
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 14182 4808 14188 4820
rect 14143 4780 14188 4808
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 15102 4808 15108 4820
rect 15063 4780 15108 4808
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 16853 4811 16911 4817
rect 16853 4777 16865 4811
rect 16899 4808 16911 4811
rect 17313 4811 17371 4817
rect 17313 4808 17325 4811
rect 16899 4780 17325 4808
rect 16899 4777 16911 4780
rect 16853 4771 16911 4777
rect 17313 4777 17325 4780
rect 17359 4808 17371 4811
rect 17862 4808 17868 4820
rect 17359 4780 17868 4808
rect 17359 4777 17371 4780
rect 17313 4771 17371 4777
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 18138 4808 18144 4820
rect 18099 4780 18144 4808
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18230 4768 18236 4820
rect 18288 4808 18294 4820
rect 18874 4808 18880 4820
rect 18288 4780 18880 4808
rect 18288 4768 18294 4780
rect 18874 4768 18880 4780
rect 18932 4808 18938 4820
rect 19978 4808 19984 4820
rect 18932 4780 19104 4808
rect 19939 4780 19984 4808
rect 18932 4768 18938 4780
rect 17405 4743 17463 4749
rect 17405 4709 17417 4743
rect 17451 4740 17463 4743
rect 17494 4740 17500 4752
rect 17451 4712 17500 4740
rect 17451 4709 17463 4712
rect 17405 4703 17463 4709
rect 17494 4700 17500 4712
rect 17552 4700 17558 4752
rect 17678 4700 17684 4752
rect 17736 4740 17742 4752
rect 19076 4740 19104 4780
rect 19978 4768 19984 4780
rect 20036 4768 20042 4820
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 21266 4808 21272 4820
rect 20763 4780 21272 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 22925 4811 22983 4817
rect 22925 4777 22937 4811
rect 22971 4808 22983 4811
rect 23290 4808 23296 4820
rect 22971 4780 23296 4808
rect 22971 4777 22983 4780
rect 22925 4771 22983 4777
rect 23290 4768 23296 4780
rect 23348 4808 23354 4820
rect 23474 4808 23480 4820
rect 23348 4780 23480 4808
rect 23348 4768 23354 4780
rect 23474 4768 23480 4780
rect 23532 4768 23538 4820
rect 20070 4740 20076 4752
rect 17736 4712 19012 4740
rect 19076 4712 20076 4740
rect 17736 4700 17742 4712
rect 12066 4632 12072 4684
rect 12124 4672 12130 4684
rect 12434 4681 12440 4684
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 12124 4644 12173 4672
rect 12124 4632 12130 4644
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 12428 4635 12440 4681
rect 12492 4672 12498 4684
rect 12492 4644 12528 4672
rect 12434 4632 12440 4635
rect 12492 4632 12498 4644
rect 15470 4632 15476 4684
rect 15528 4672 15534 4684
rect 18984 4681 19012 4712
rect 20070 4700 20076 4712
rect 20128 4700 20134 4752
rect 23842 4700 23848 4752
rect 23900 4740 23906 4752
rect 24946 4740 24952 4752
rect 23900 4712 24952 4740
rect 23900 4700 23906 4712
rect 24946 4700 24952 4712
rect 25004 4700 25010 4752
rect 15841 4675 15899 4681
rect 15841 4672 15853 4675
rect 15528 4644 15853 4672
rect 15528 4632 15534 4644
rect 15841 4641 15853 4644
rect 15887 4641 15899 4675
rect 15841 4635 15899 4641
rect 18969 4675 19027 4681
rect 18969 4641 18981 4675
rect 19015 4672 19027 4675
rect 19150 4672 19156 4684
rect 19015 4644 19156 4672
rect 19015 4641 19027 4644
rect 18969 4635 19027 4641
rect 19150 4632 19156 4644
rect 19208 4632 19214 4684
rect 20990 4632 20996 4684
rect 21048 4672 21054 4684
rect 21157 4675 21215 4681
rect 21157 4672 21169 4675
rect 21048 4644 21169 4672
rect 21048 4632 21054 4644
rect 21157 4641 21169 4644
rect 21203 4641 21215 4675
rect 23198 4672 23204 4684
rect 21157 4635 21215 4641
rect 22296 4644 23204 4672
rect 17494 4564 17500 4616
rect 17552 4604 17558 4616
rect 17770 4604 17776 4616
rect 17552 4576 17776 4604
rect 17552 4564 17558 4576
rect 17770 4564 17776 4576
rect 17828 4564 17834 4616
rect 19058 4604 19064 4616
rect 19019 4576 19064 4604
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 19610 4564 19616 4616
rect 19668 4604 19674 4616
rect 20806 4604 20812 4616
rect 19668 4576 20812 4604
rect 19668 4564 19674 4576
rect 20806 4564 20812 4576
rect 20864 4604 20870 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20864 4576 20913 4604
rect 20864 4564 20870 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 16485 4539 16543 4545
rect 16485 4505 16497 4539
rect 16531 4536 16543 4539
rect 18509 4539 18567 4545
rect 18509 4536 18521 4539
rect 16531 4508 18521 4536
rect 16531 4505 16543 4508
rect 16485 4499 16543 4505
rect 18509 4505 18521 4508
rect 18555 4536 18567 4539
rect 19242 4536 19248 4548
rect 18555 4508 19248 4536
rect 18555 4505 18567 4508
rect 18509 4499 18567 4505
rect 19242 4496 19248 4508
rect 19300 4496 19306 4548
rect 22296 4545 22324 4644
rect 23198 4632 23204 4644
rect 23256 4672 23262 4684
rect 23641 4675 23699 4681
rect 23641 4672 23653 4675
rect 23256 4644 23653 4672
rect 23256 4632 23262 4644
rect 23641 4641 23653 4644
rect 23687 4641 23699 4675
rect 23641 4635 23699 4641
rect 23385 4607 23443 4613
rect 23385 4604 23397 4607
rect 23216 4576 23397 4604
rect 22281 4539 22339 4545
rect 22281 4505 22293 4539
rect 22327 4505 22339 4539
rect 22281 4499 22339 4505
rect 14734 4468 14740 4480
rect 14695 4440 14740 4468
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 15565 4471 15623 4477
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 15838 4468 15844 4480
rect 15611 4440 15844 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 16022 4468 16028 4480
rect 15983 4440 16028 4468
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 16945 4471 17003 4477
rect 16945 4468 16957 4471
rect 16632 4440 16957 4468
rect 16632 4428 16638 4440
rect 16945 4437 16957 4440
rect 16991 4437 17003 4471
rect 16945 4431 17003 4437
rect 19518 4428 19524 4480
rect 19576 4468 19582 4480
rect 19705 4471 19763 4477
rect 19705 4468 19717 4471
rect 19576 4440 19717 4468
rect 19576 4428 19582 4440
rect 19705 4437 19717 4440
rect 19751 4468 19763 4471
rect 19978 4468 19984 4480
rect 19751 4440 19984 4468
rect 19751 4437 19763 4440
rect 19705 4431 19763 4437
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 23106 4428 23112 4480
rect 23164 4468 23170 4480
rect 23216 4477 23244 4576
rect 23385 4573 23397 4576
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 23201 4471 23259 4477
rect 23201 4468 23213 4471
rect 23164 4440 23213 4468
rect 23164 4428 23170 4440
rect 23201 4437 23213 4440
rect 23247 4437 23259 4471
rect 24762 4468 24768 4480
rect 24723 4440 24768 4468
rect 23201 4431 23259 4437
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 12066 4224 12072 4276
rect 12124 4264 12130 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 12124 4236 12173 4264
rect 12124 4224 12130 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 12161 4227 12219 4233
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6822 4128 6828 4140
rect 6420 4100 6828 4128
rect 6420 4088 6426 4100
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 8202 4128 8208 4140
rect 7800 4100 8208 4128
rect 7800 4088 7806 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4029 11391 4063
rect 12176 4060 12204 4227
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 12621 4267 12679 4273
rect 12621 4264 12633 4267
rect 12492 4236 12633 4264
rect 12492 4224 12498 4236
rect 12621 4233 12633 4236
rect 12667 4233 12679 4267
rect 12621 4227 12679 4233
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 12768 4236 15424 4264
rect 12768 4224 12774 4236
rect 15396 4196 15424 4236
rect 15470 4224 15476 4276
rect 15528 4264 15534 4276
rect 15841 4267 15899 4273
rect 15841 4264 15853 4267
rect 15528 4236 15853 4264
rect 15528 4224 15534 4236
rect 15841 4233 15853 4236
rect 15887 4233 15899 4267
rect 15841 4227 15899 4233
rect 17221 4267 17279 4273
rect 17221 4233 17233 4267
rect 17267 4264 17279 4267
rect 17402 4264 17408 4276
rect 17267 4236 17408 4264
rect 17267 4233 17279 4236
rect 17221 4227 17279 4233
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 20530 4224 20536 4276
rect 20588 4264 20594 4276
rect 20990 4264 20996 4276
rect 20588 4236 20996 4264
rect 20588 4224 20594 4236
rect 20990 4224 20996 4236
rect 21048 4264 21054 4276
rect 21913 4267 21971 4273
rect 21913 4264 21925 4267
rect 21048 4236 21925 4264
rect 21048 4224 21054 4236
rect 21913 4233 21925 4236
rect 21959 4233 21971 4267
rect 25038 4264 25044 4276
rect 24999 4236 25044 4264
rect 21913 4227 21971 4233
rect 25038 4224 25044 4236
rect 25096 4224 25102 4276
rect 17681 4199 17739 4205
rect 17681 4196 17693 4199
rect 15396 4168 17693 4196
rect 17681 4165 17693 4168
rect 17727 4196 17739 4199
rect 17773 4199 17831 4205
rect 17773 4196 17785 4199
rect 17727 4168 17785 4196
rect 17727 4165 17739 4168
rect 17681 4159 17739 4165
rect 17773 4165 17785 4168
rect 17819 4165 17831 4199
rect 17773 4159 17831 4165
rect 18049 4199 18107 4205
rect 18049 4165 18061 4199
rect 18095 4165 18107 4199
rect 18049 4159 18107 4165
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 13262 4128 13268 4140
rect 12584 4100 13268 4128
rect 12584 4088 12590 4100
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4128 15623 4131
rect 16666 4128 16672 4140
rect 15611 4100 16672 4128
rect 15611 4097 15623 4100
rect 15565 4091 15623 4097
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 18064 4128 18092 4159
rect 18138 4156 18144 4208
rect 18196 4196 18202 4208
rect 19058 4196 19064 4208
rect 18196 4168 19064 4196
rect 18196 4156 18202 4168
rect 16776 4100 18092 4128
rect 13173 4063 13231 4069
rect 13173 4060 13185 4063
rect 12176 4032 13185 4060
rect 11333 4023 11391 4029
rect 13173 4029 13185 4032
rect 13219 4060 13231 4063
rect 13357 4063 13415 4069
rect 13357 4060 13369 4063
rect 13219 4032 13369 4060
rect 13219 4029 13231 4032
rect 13173 4023 13231 4029
rect 13357 4029 13369 4032
rect 13403 4060 13415 4063
rect 13906 4060 13912 4072
rect 13403 4032 13912 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 11348 3992 11376 4023
rect 13906 4020 13912 4032
rect 13964 4020 13970 4072
rect 16574 4060 16580 4072
rect 16535 4032 16580 4060
rect 16574 4020 16580 4032
rect 16632 4060 16638 4072
rect 16776 4060 16804 4100
rect 18230 4088 18236 4140
rect 18288 4128 18294 4140
rect 18616 4137 18644 4168
rect 19058 4156 19064 4168
rect 19116 4196 19122 4208
rect 19116 4168 19288 4196
rect 19116 4156 19122 4168
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 18288 4100 18521 4128
rect 18288 4088 18294 4100
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 19260 4128 19288 4168
rect 20806 4156 20812 4208
rect 20864 4196 20870 4208
rect 21545 4199 21603 4205
rect 21545 4196 21557 4199
rect 20864 4168 21557 4196
rect 20864 4156 20870 4168
rect 21545 4165 21557 4168
rect 21591 4196 21603 4199
rect 23106 4196 23112 4208
rect 21591 4168 23112 4196
rect 21591 4165 21603 4168
rect 21545 4159 21603 4165
rect 23106 4156 23112 4168
rect 23164 4196 23170 4208
rect 23385 4199 23443 4205
rect 23385 4196 23397 4199
rect 23164 4168 23397 4196
rect 23164 4156 23170 4168
rect 23385 4165 23397 4168
rect 23431 4196 23443 4199
rect 23431 4168 23704 4196
rect 23431 4165 23443 4168
rect 23385 4159 23443 4165
rect 19518 4128 19524 4140
rect 19260 4100 19524 4128
rect 18601 4091 18659 4097
rect 19518 4088 19524 4100
rect 19576 4088 19582 4140
rect 23676 4137 23704 4168
rect 23661 4131 23719 4137
rect 23661 4097 23673 4131
rect 23707 4097 23719 4131
rect 23661 4091 23719 4097
rect 16632 4032 16804 4060
rect 17681 4063 17739 4069
rect 16632 4020 16638 4032
rect 17681 4029 17693 4063
rect 17727 4060 17739 4063
rect 18322 4060 18328 4072
rect 17727 4032 18328 4060
rect 17727 4029 17739 4032
rect 17681 4023 17739 4029
rect 18322 4020 18328 4032
rect 18380 4060 18386 4072
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18380 4032 18429 4060
rect 18380 4020 18386 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 19150 4060 19156 4072
rect 19111 4032 19156 4060
rect 18417 4023 18475 4029
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 19610 4060 19616 4072
rect 19444 4032 19616 4060
rect 11885 3995 11943 4001
rect 11885 3992 11897 3995
rect 11348 3964 11897 3992
rect 11885 3961 11897 3964
rect 11931 3992 11943 3995
rect 12342 3992 12348 4004
rect 11931 3964 12348 3992
rect 11931 3961 11943 3964
rect 11885 3955 11943 3961
rect 12342 3952 12348 3964
rect 12400 3952 12406 4004
rect 13538 3952 13544 4004
rect 13596 4001 13602 4004
rect 13596 3995 13660 4001
rect 13596 3961 13614 3995
rect 13648 3961 13660 3995
rect 13596 3955 13660 3961
rect 13596 3952 13602 3955
rect 16206 3952 16212 4004
rect 16264 3992 16270 4004
rect 16485 3995 16543 4001
rect 16485 3992 16497 3995
rect 16264 3964 16497 3992
rect 16264 3952 16270 3964
rect 16485 3961 16497 3964
rect 16531 3961 16543 3995
rect 16485 3955 16543 3961
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11204 3896 11529 3924
rect 11204 3884 11210 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3924 14795 3927
rect 14826 3924 14832 3936
rect 14783 3896 14832 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 16298 3924 16304 3936
rect 16163 3896 16304 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 19444 3933 19472 4032
rect 19610 4020 19616 4032
rect 19668 4020 19674 4072
rect 22186 4060 22192 4072
rect 22147 4032 22192 4060
rect 22186 4020 22192 4032
rect 22244 4060 22250 4072
rect 22741 4063 22799 4069
rect 22741 4060 22753 4063
rect 22244 4032 22753 4060
rect 22244 4020 22250 4032
rect 22741 4029 22753 4032
rect 22787 4029 22799 4063
rect 22741 4023 22799 4029
rect 19880 3995 19938 4001
rect 19880 3961 19892 3995
rect 19926 3992 19938 3995
rect 19978 3992 19984 4004
rect 19926 3964 19984 3992
rect 19926 3961 19938 3964
rect 19880 3955 19938 3961
rect 19978 3952 19984 3964
rect 20036 3952 20042 4004
rect 23842 3952 23848 4004
rect 23900 4001 23906 4004
rect 23900 3995 23964 4001
rect 23900 3961 23918 3995
rect 23952 3961 23964 3995
rect 23900 3955 23964 3961
rect 23900 3952 23906 3955
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 18288 3896 19441 3924
rect 18288 3884 18294 3896
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 22370 3924 22376 3936
rect 22331 3896 22376 3924
rect 19429 3887 19487 3893
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 12710 3720 12716 3732
rect 12671 3692 12716 3720
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 13449 3723 13507 3729
rect 13449 3689 13461 3723
rect 13495 3720 13507 3723
rect 13538 3720 13544 3732
rect 13495 3692 13544 3720
rect 13495 3689 13507 3692
rect 13449 3683 13507 3689
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 14090 3720 14096 3732
rect 14051 3692 14096 3720
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 18601 3723 18659 3729
rect 18601 3689 18613 3723
rect 18647 3720 18659 3723
rect 18874 3720 18880 3732
rect 18647 3692 18880 3720
rect 18647 3689 18659 3692
rect 18601 3683 18659 3689
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 19242 3720 19248 3732
rect 19203 3692 19248 3720
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 19889 3723 19947 3729
rect 19889 3720 19901 3723
rect 19576 3692 19901 3720
rect 19576 3680 19582 3692
rect 19889 3689 19901 3692
rect 19935 3689 19947 3723
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 19889 3683 19947 3689
rect 20714 3680 20720 3692
rect 20772 3720 20778 3732
rect 21269 3723 21327 3729
rect 21269 3720 21281 3723
rect 20772 3692 21281 3720
rect 20772 3680 20778 3692
rect 21269 3689 21281 3692
rect 21315 3689 21327 3723
rect 21269 3683 21327 3689
rect 22094 3680 22100 3732
rect 22152 3720 22158 3732
rect 22462 3720 22468 3732
rect 22152 3692 22197 3720
rect 22423 3692 22468 3720
rect 22152 3680 22158 3692
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 23290 3720 23296 3732
rect 23251 3692 23296 3720
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 24854 3720 24860 3732
rect 24815 3692 24860 3720
rect 24854 3680 24860 3692
rect 24912 3680 24918 3732
rect 24946 3680 24952 3732
rect 25004 3720 25010 3732
rect 25225 3723 25283 3729
rect 25225 3720 25237 3723
rect 25004 3692 25237 3720
rect 25004 3680 25010 3692
rect 25225 3689 25237 3692
rect 25271 3689 25283 3723
rect 25225 3683 25283 3689
rect 13906 3612 13912 3664
rect 13964 3652 13970 3664
rect 14550 3652 14556 3664
rect 13964 3624 14556 3652
rect 13964 3612 13970 3624
rect 14550 3612 14556 3624
rect 14608 3652 14614 3664
rect 14645 3655 14703 3661
rect 14645 3652 14657 3655
rect 14608 3624 14657 3652
rect 14608 3612 14614 3624
rect 14645 3621 14657 3624
rect 14691 3652 14703 3655
rect 14691 3624 16436 3652
rect 14691 3621 14703 3624
rect 14645 3615 14703 3621
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3584 10471 3587
rect 10686 3584 10692 3596
rect 10459 3556 10692 3584
rect 10459 3553 10471 3556
rect 10413 3547 10471 3553
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 11425 3587 11483 3593
rect 11425 3584 11437 3587
rect 11388 3556 11437 3584
rect 11388 3544 11394 3556
rect 11425 3553 11437 3556
rect 11471 3553 11483 3587
rect 11425 3547 11483 3553
rect 12529 3587 12587 3593
rect 12529 3553 12541 3587
rect 12575 3584 12587 3587
rect 12986 3584 12992 3596
rect 12575 3556 12992 3584
rect 12575 3553 12587 3556
rect 12529 3547 12587 3553
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 14001 3587 14059 3593
rect 14001 3553 14013 3587
rect 14047 3584 14059 3587
rect 14182 3584 14188 3596
rect 14047 3556 14188 3584
rect 14047 3553 14059 3556
rect 14001 3547 14059 3553
rect 14182 3544 14188 3556
rect 14240 3584 14246 3596
rect 15289 3587 15347 3593
rect 14240 3556 15148 3584
rect 14240 3544 14246 3556
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14826 3516 14832 3528
rect 14323 3488 14832 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15120 3516 15148 3556
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 15654 3584 15660 3596
rect 15335 3556 15660 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 16408 3593 16436 3624
rect 21450 3612 21456 3664
rect 21508 3652 21514 3664
rect 22557 3655 22615 3661
rect 22557 3652 22569 3655
rect 21508 3624 22569 3652
rect 21508 3612 21514 3624
rect 22557 3621 22569 3624
rect 22603 3621 22615 3655
rect 22738 3652 22744 3664
rect 22699 3624 22744 3652
rect 22557 3615 22615 3621
rect 22738 3612 22744 3624
rect 22796 3612 22802 3664
rect 23198 3652 23204 3664
rect 23159 3624 23204 3652
rect 23198 3612 23204 3624
rect 23256 3612 23262 3664
rect 16393 3587 16451 3593
rect 16393 3553 16405 3587
rect 16439 3584 16451 3587
rect 16482 3584 16488 3596
rect 16439 3556 16488 3584
rect 16439 3553 16451 3556
rect 16393 3547 16451 3553
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 16666 3593 16672 3596
rect 16660 3584 16672 3593
rect 16627 3556 16672 3584
rect 16660 3547 16672 3556
rect 16666 3544 16672 3547
rect 16724 3544 16730 3596
rect 15378 3516 15384 3528
rect 15120 3488 15384 3516
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 19150 3476 19156 3528
rect 19208 3516 19214 3528
rect 19337 3519 19395 3525
rect 19337 3516 19349 3519
rect 19208 3488 19349 3516
rect 19208 3476 19214 3488
rect 19337 3485 19349 3488
rect 19383 3485 19395 3519
rect 19337 3479 19395 3485
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 13630 3448 13636 3460
rect 13591 3420 13636 3448
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 19058 3408 19064 3460
rect 19116 3448 19122 3460
rect 19444 3448 19472 3479
rect 19610 3476 19616 3528
rect 19668 3516 19674 3528
rect 21358 3516 21364 3528
rect 19668 3488 21364 3516
rect 19668 3476 19674 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21545 3519 21603 3525
rect 21545 3485 21557 3519
rect 21591 3516 21603 3519
rect 21726 3516 21732 3528
rect 21591 3488 21732 3516
rect 21591 3485 21603 3488
rect 21545 3479 21603 3485
rect 21726 3476 21732 3488
rect 21784 3516 21790 3528
rect 23216 3516 23244 3612
rect 23661 3587 23719 3593
rect 23661 3584 23673 3587
rect 21784 3488 23244 3516
rect 23584 3556 23673 3584
rect 21784 3476 21790 3488
rect 20898 3448 20904 3460
rect 19116 3420 19472 3448
rect 20859 3420 20904 3448
rect 19116 3408 19122 3420
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 22557 3451 22615 3457
rect 22557 3417 22569 3451
rect 22603 3448 22615 3451
rect 23290 3448 23296 3460
rect 22603 3420 23296 3448
rect 22603 3417 22615 3420
rect 22557 3411 22615 3417
rect 23290 3408 23296 3420
rect 23348 3448 23354 3460
rect 23584 3448 23612 3556
rect 23661 3553 23673 3556
rect 23707 3553 23719 3587
rect 23661 3547 23719 3553
rect 23750 3516 23756 3528
rect 23711 3488 23756 3516
rect 23750 3476 23756 3488
rect 23808 3476 23814 3528
rect 23842 3476 23848 3528
rect 23900 3516 23906 3528
rect 23937 3519 23995 3525
rect 23937 3516 23949 3519
rect 23900 3488 23949 3516
rect 23900 3476 23906 3488
rect 23937 3485 23949 3488
rect 23983 3516 23995 3519
rect 23983 3488 24440 3516
rect 23983 3485 23995 3488
rect 23937 3479 23995 3485
rect 24412 3457 24440 3488
rect 24854 3476 24860 3528
rect 24912 3516 24918 3528
rect 25317 3519 25375 3525
rect 25317 3516 25329 3519
rect 24912 3488 25329 3516
rect 24912 3476 24918 3488
rect 25317 3485 25329 3488
rect 25363 3485 25375 3519
rect 25498 3516 25504 3528
rect 25459 3488 25504 3516
rect 25317 3479 25375 3485
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 23348 3420 23612 3448
rect 24397 3451 24455 3457
rect 23348 3408 23354 3420
rect 24397 3417 24409 3451
rect 24443 3448 24455 3451
rect 24762 3448 24768 3460
rect 24443 3420 24768 3448
rect 24443 3417 24455 3420
rect 24397 3411 24455 3417
rect 24762 3408 24768 3420
rect 24820 3448 24826 3460
rect 25516 3448 25544 3476
rect 24820 3420 25544 3448
rect 24820 3408 24826 3420
rect 10597 3383 10655 3389
rect 10597 3349 10609 3383
rect 10643 3380 10655 3383
rect 10870 3380 10876 3392
rect 10643 3352 10876 3380
rect 10643 3349 10655 3352
rect 10597 3343 10655 3349
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 11606 3380 11612 3392
rect 11567 3352 11612 3380
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 14826 3340 14832 3392
rect 14884 3380 14890 3392
rect 15013 3383 15071 3389
rect 15013 3380 15025 3383
rect 14884 3352 15025 3380
rect 14884 3340 14890 3352
rect 15013 3349 15025 3352
rect 15059 3349 15071 3383
rect 15470 3380 15476 3392
rect 15431 3352 15476 3380
rect 15013 3343 15071 3349
rect 15470 3340 15476 3352
rect 15528 3340 15534 3392
rect 17402 3340 17408 3392
rect 17460 3380 17466 3392
rect 17773 3383 17831 3389
rect 17773 3380 17785 3383
rect 17460 3352 17785 3380
rect 17460 3340 17466 3352
rect 17773 3349 17785 3352
rect 17819 3349 17831 3383
rect 18874 3380 18880 3392
rect 18835 3352 18880 3380
rect 17773 3343 17831 3349
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 20346 3380 20352 3392
rect 20307 3352 20352 3380
rect 20346 3340 20352 3352
rect 20404 3340 20410 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 10134 3176 10140 3188
rect 10095 3148 10140 3176
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 10686 3176 10692 3188
rect 10647 3148 10692 3176
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 11146 3176 11152 3188
rect 11107 3148 11152 3176
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 12986 3176 12992 3188
rect 12947 3148 12992 3176
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13357 3179 13415 3185
rect 13357 3145 13369 3179
rect 13403 3176 13415 3179
rect 13446 3176 13452 3188
rect 13403 3148 13452 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 14093 3179 14151 3185
rect 14093 3145 14105 3179
rect 14139 3176 14151 3179
rect 14182 3176 14188 3188
rect 14139 3148 14188 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 16482 3176 16488 3188
rect 16443 3148 16488 3176
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 17037 3179 17095 3185
rect 17037 3145 17049 3179
rect 17083 3176 17095 3179
rect 17494 3176 17500 3188
rect 17083 3148 17500 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 20346 3136 20352 3188
rect 20404 3176 20410 3188
rect 20717 3179 20775 3185
rect 20717 3176 20729 3179
rect 20404 3148 20729 3176
rect 20404 3136 20410 3148
rect 20717 3145 20729 3148
rect 20763 3145 20775 3179
rect 21726 3176 21732 3188
rect 21687 3148 21732 3176
rect 20717 3139 20775 3145
rect 21726 3136 21732 3148
rect 21784 3136 21790 3188
rect 23290 3176 23296 3188
rect 23251 3148 23296 3176
rect 23290 3136 23296 3148
rect 23348 3136 23354 3188
rect 23750 3136 23756 3188
rect 23808 3176 23814 3188
rect 23845 3179 23903 3185
rect 23845 3176 23857 3179
rect 23808 3148 23857 3176
rect 23808 3136 23814 3148
rect 23845 3145 23857 3148
rect 23891 3145 23903 3179
rect 23845 3139 23903 3145
rect 24854 3136 24860 3188
rect 24912 3176 24918 3188
rect 25133 3179 25191 3185
rect 25133 3176 25145 3179
rect 24912 3148 25145 3176
rect 24912 3136 24918 3148
rect 25133 3145 25145 3148
rect 25179 3145 25191 3179
rect 25133 3139 25191 3145
rect 25498 3136 25504 3188
rect 25556 3176 25562 3188
rect 25869 3179 25927 3185
rect 25869 3176 25881 3179
rect 25556 3148 25881 3176
rect 25556 3136 25562 3148
rect 25869 3145 25881 3148
rect 25915 3145 25927 3179
rect 25869 3139 25927 3145
rect 10413 3111 10471 3117
rect 10413 3077 10425 3111
rect 10459 3108 10471 3111
rect 11054 3108 11060 3120
rect 10459 3080 11060 3108
rect 10459 3077 10471 3080
rect 10413 3071 10471 3077
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 10778 3040 10784 3052
rect 9815 3012 10784 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9784 2972 9812 3003
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 9263 2944 9812 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 10192 2944 10241 2972
rect 10192 2932 10198 2944
rect 10229 2941 10241 2944
rect 10275 2941 10287 2975
rect 10229 2935 10287 2941
rect 10686 2932 10692 2984
rect 10744 2972 10750 2984
rect 10962 2972 10968 2984
rect 10744 2944 10968 2972
rect 10744 2932 10750 2944
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 11164 2972 11192 3136
rect 11422 3108 11428 3120
rect 11383 3080 11428 3108
rect 11422 3068 11428 3080
rect 11480 3068 11486 3120
rect 15933 3111 15991 3117
rect 15933 3077 15945 3111
rect 15979 3108 15991 3111
rect 16666 3108 16672 3120
rect 15979 3080 16672 3108
rect 15979 3077 15991 3080
rect 15933 3071 15991 3077
rect 16666 3068 16672 3080
rect 16724 3108 16730 3120
rect 17126 3108 17132 3120
rect 16724 3080 17132 3108
rect 16724 3068 16730 3080
rect 17126 3068 17132 3080
rect 17184 3068 17190 3120
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3077 19671 3111
rect 19613 3071 19671 3077
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12492 3012 12537 3040
rect 12492 3000 12498 3012
rect 14090 3000 14096 3052
rect 14148 3040 14154 3052
rect 14369 3043 14427 3049
rect 14369 3040 14381 3043
rect 14148 3012 14381 3040
rect 14148 3000 14154 3012
rect 14369 3009 14381 3012
rect 14415 3009 14427 3043
rect 14550 3040 14556 3052
rect 14511 3012 14556 3040
rect 14369 3003 14427 3009
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 17773 3043 17831 3049
rect 17773 3040 17785 3043
rect 16540 3012 17785 3040
rect 16540 3000 16546 3012
rect 17773 3009 17785 3012
rect 17819 3040 17831 3043
rect 18230 3040 18236 3052
rect 17819 3012 18236 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 19628 3040 19656 3071
rect 21358 3068 21364 3120
rect 21416 3108 21422 3120
rect 22097 3111 22155 3117
rect 22097 3108 22109 3111
rect 21416 3080 22109 3108
rect 21416 3068 21422 3080
rect 22097 3077 22109 3080
rect 22143 3077 22155 3111
rect 23308 3108 23336 3136
rect 24397 3111 24455 3117
rect 24397 3108 24409 3111
rect 23308 3080 24409 3108
rect 22097 3071 22155 3077
rect 24397 3077 24409 3080
rect 24443 3077 24455 3111
rect 24397 3071 24455 3077
rect 19978 3040 19984 3052
rect 19628 3012 19984 3040
rect 19978 3000 19984 3012
rect 20036 3040 20042 3052
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 20036 3012 20269 3040
rect 20036 3000 20042 3012
rect 20257 3009 20269 3012
rect 20303 3040 20315 3043
rect 21269 3043 21327 3049
rect 21269 3040 21281 3043
rect 20303 3012 21281 3040
rect 20303 3009 20315 3012
rect 20257 3003 20315 3009
rect 21269 3009 21281 3012
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 11164 2944 11253 2972
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 13446 2972 13452 2984
rect 13407 2944 13452 2972
rect 11241 2935 11299 2941
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 19484 2944 20545 2972
rect 19484 2932 19490 2944
rect 20533 2941 20545 2944
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 11330 2904 11336 2916
rect 9416 2876 11336 2904
rect 9416 2845 9444 2876
rect 11330 2864 11336 2876
rect 11388 2904 11394 2916
rect 14826 2913 14832 2916
rect 11793 2907 11851 2913
rect 11793 2904 11805 2907
rect 11388 2876 11805 2904
rect 11388 2864 11394 2876
rect 11793 2873 11805 2876
rect 11839 2873 11851 2907
rect 14820 2904 14832 2913
rect 14787 2876 14832 2904
rect 11793 2867 11851 2873
rect 14820 2867 14832 2876
rect 14826 2864 14832 2867
rect 14884 2864 14890 2916
rect 18478 2907 18536 2913
rect 18478 2873 18490 2907
rect 18524 2873 18536 2907
rect 20548 2904 20576 2935
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 21082 2972 21088 2984
rect 20864 2944 21088 2972
rect 20864 2932 20870 2944
rect 21082 2932 21088 2944
rect 21140 2932 21146 2984
rect 22465 2975 22523 2981
rect 22465 2941 22477 2975
rect 22511 2972 22523 2975
rect 22554 2972 22560 2984
rect 22511 2944 22560 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 24412 2972 24440 3071
rect 24946 3000 24952 3052
rect 25004 3040 25010 3052
rect 25501 3043 25559 3049
rect 25501 3040 25513 3043
rect 25004 3012 25513 3040
rect 25004 3000 25010 3012
rect 25501 3009 25513 3012
rect 25547 3009 25559 3043
rect 25501 3003 25559 3009
rect 24581 2975 24639 2981
rect 24581 2972 24593 2975
rect 24412 2944 24593 2972
rect 24581 2941 24593 2944
rect 24627 2941 24639 2975
rect 24581 2935 24639 2941
rect 21177 2907 21235 2913
rect 21177 2904 21189 2907
rect 20548 2876 21189 2904
rect 18478 2867 18536 2873
rect 21177 2873 21189 2876
rect 21223 2904 21235 2907
rect 21450 2904 21456 2916
rect 21223 2876 21456 2904
rect 21223 2873 21235 2876
rect 21177 2867 21235 2873
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2805 9459 2839
rect 13630 2836 13636 2848
rect 13591 2808 13636 2836
rect 9401 2799 9459 2805
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 17402 2836 17408 2848
rect 17363 2808 17408 2836
rect 17402 2796 17408 2808
rect 17460 2836 17466 2848
rect 18493 2836 18521 2867
rect 21450 2864 21456 2876
rect 21508 2864 21514 2916
rect 22646 2836 22652 2848
rect 17460 2808 18521 2836
rect 22607 2808 22652 2836
rect 17460 2796 17466 2808
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 24762 2836 24768 2848
rect 24723 2808 24768 2836
rect 24762 2796 24768 2808
rect 24820 2796 24826 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2958 2632 2964 2644
rect 2919 2604 2964 2632
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 5718 2632 5724 2644
rect 5679 2604 5724 2632
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 13078 2632 13084 2644
rect 13039 2604 13084 2632
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 16025 2635 16083 2641
rect 16025 2632 16037 2635
rect 14792 2604 16037 2632
rect 14792 2592 14798 2604
rect 16025 2601 16037 2604
rect 16071 2601 16083 2635
rect 16025 2595 16083 2601
rect 16114 2592 16120 2644
rect 16172 2632 16178 2644
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 16172 2604 16497 2632
rect 16172 2592 16178 2604
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 17126 2632 17132 2644
rect 17039 2604 17132 2632
rect 16485 2595 16543 2601
rect 17126 2592 17132 2604
rect 17184 2632 17190 2644
rect 19058 2632 19064 2644
rect 17184 2604 19064 2632
rect 17184 2592 17190 2604
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 19518 2632 19524 2644
rect 19479 2604 19524 2632
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 19889 2635 19947 2641
rect 19889 2601 19901 2635
rect 19935 2632 19947 2635
rect 20346 2632 20352 2644
rect 19935 2604 20352 2632
rect 19935 2601 19947 2604
rect 19889 2595 19947 2601
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 20806 2632 20812 2644
rect 20767 2604 20812 2632
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 22462 2592 22468 2644
rect 22520 2632 22526 2644
rect 22649 2635 22707 2641
rect 22649 2632 22661 2635
rect 22520 2604 22661 2632
rect 22520 2592 22526 2604
rect 22649 2601 22661 2604
rect 22695 2601 22707 2635
rect 23842 2632 23848 2644
rect 23803 2604 23848 2632
rect 22649 2595 22707 2601
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 2958 2496 2964 2508
rect 2823 2468 2964 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 2958 2456 2964 2468
rect 3016 2496 3022 2508
rect 3329 2499 3387 2505
rect 3329 2496 3341 2499
rect 3016 2468 3341 2496
rect 3016 2456 3022 2468
rect 3329 2465 3341 2468
rect 3375 2465 3387 2499
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 3329 2459 3387 2465
rect 5534 2456 5540 2468
rect 5592 2496 5598 2508
rect 6089 2499 6147 2505
rect 6089 2496 6101 2499
rect 5592 2468 6101 2496
rect 5592 2456 5598 2468
rect 6089 2465 6101 2468
rect 6135 2465 6147 2499
rect 6089 2459 6147 2465
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8386 2496 8392 2508
rect 8159 2468 8392 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 10888 2496 10916 2592
rect 11514 2524 11520 2576
rect 11572 2564 11578 2576
rect 13725 2567 13783 2573
rect 13725 2564 13737 2567
rect 11572 2536 13737 2564
rect 11572 2524 11578 2536
rect 10367 2468 10916 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 13188 2505 13216 2536
rect 13725 2533 13737 2536
rect 13771 2533 13783 2567
rect 13725 2527 13783 2533
rect 14185 2567 14243 2573
rect 14185 2533 14197 2567
rect 14231 2564 14243 2567
rect 14826 2564 14832 2576
rect 14231 2536 14832 2564
rect 14231 2533 14243 2536
rect 14185 2527 14243 2533
rect 14826 2524 14832 2536
rect 14884 2524 14890 2576
rect 15746 2564 15752 2576
rect 15707 2536 15752 2564
rect 15746 2524 15752 2536
rect 15804 2524 15810 2576
rect 16298 2564 16304 2576
rect 16211 2536 16304 2564
rect 16298 2524 16304 2536
rect 16356 2564 16362 2576
rect 16393 2567 16451 2573
rect 16393 2564 16405 2567
rect 16356 2536 16405 2564
rect 16356 2524 16362 2536
rect 16393 2533 16405 2536
rect 16439 2533 16451 2567
rect 18046 2564 18052 2576
rect 18007 2536 18052 2564
rect 16393 2527 16451 2533
rect 18046 2524 18052 2536
rect 18104 2524 18110 2576
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 11112 2468 11437 2496
rect 11112 2456 11118 2468
rect 11425 2465 11437 2468
rect 11471 2496 11483 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11471 2468 11989 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14642 2496 14648 2508
rect 14323 2468 14648 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 14642 2456 14648 2468
rect 14700 2496 14706 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14700 2468 14933 2496
rect 14700 2456 14706 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 16316 2428 16344 2524
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 18414 2496 18420 2508
rect 17819 2468 18420 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 19429 2499 19487 2505
rect 19429 2465 19441 2499
rect 19475 2496 19487 2499
rect 20530 2496 20536 2508
rect 19475 2468 20536 2496
rect 19475 2465 19487 2468
rect 19429 2459 19487 2465
rect 12483 2400 16344 2428
rect 16577 2431 16635 2437
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 16577 2397 16589 2431
rect 16623 2428 16635 2431
rect 17402 2428 17408 2440
rect 16623 2400 17408 2428
rect 16623 2397 16635 2400
rect 16577 2391 16635 2397
rect 14458 2360 14464 2372
rect 14419 2332 14464 2360
rect 14458 2320 14464 2332
rect 14516 2320 14522 2372
rect 15289 2363 15347 2369
rect 15289 2329 15301 2363
rect 15335 2360 15347 2363
rect 16592 2360 16620 2391
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 18966 2388 18972 2440
rect 19024 2428 19030 2440
rect 20088 2437 20116 2468
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 21634 2456 21640 2508
rect 21692 2496 21698 2508
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 21692 2468 21741 2496
rect 21692 2456 21698 2468
rect 21729 2465 21741 2468
rect 21775 2496 21787 2499
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 21775 2468 22293 2496
rect 21775 2465 21787 2468
rect 21729 2459 21787 2465
rect 22281 2465 22293 2468
rect 22327 2465 22339 2499
rect 22830 2496 22836 2508
rect 22791 2468 22836 2496
rect 22281 2459 22339 2465
rect 22830 2456 22836 2468
rect 22888 2496 22894 2508
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 22888 2468 23397 2496
rect 22888 2456 22894 2468
rect 23385 2465 23397 2468
rect 23431 2465 23443 2499
rect 23385 2459 23443 2465
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 23992 2468 24593 2496
rect 23992 2456 23998 2468
rect 24581 2465 24593 2468
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 19981 2431 20039 2437
rect 19981 2428 19993 2431
rect 19024 2400 19993 2428
rect 19024 2388 19030 2400
rect 19981 2397 19993 2400
rect 20027 2397 20039 2431
rect 19981 2391 20039 2397
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 15335 2332 16620 2360
rect 18601 2363 18659 2369
rect 15335 2329 15347 2332
rect 15289 2323 15347 2329
rect 18601 2329 18613 2363
rect 18647 2360 18659 2363
rect 19886 2360 19892 2372
rect 18647 2332 19892 2360
rect 18647 2329 18659 2332
rect 18601 2323 18659 2329
rect 19886 2320 19892 2332
rect 19944 2320 19950 2372
rect 19996 2360 20024 2391
rect 21361 2363 21419 2369
rect 21361 2360 21373 2363
rect 19996 2332 21373 2360
rect 21361 2329 21373 2332
rect 21407 2329 21419 2363
rect 21361 2323 21419 2329
rect 23017 2363 23075 2369
rect 23017 2329 23029 2363
rect 23063 2360 23075 2363
rect 24670 2360 24676 2372
rect 23063 2332 24676 2360
rect 23063 2329 23075 2332
rect 23017 2323 23075 2329
rect 24670 2320 24676 2332
rect 24728 2320 24734 2372
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 26142 2360 26148 2372
rect 24811 2332 26148 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 26142 2320 26148 2332
rect 26200 2320 26206 2372
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8444 2264 8677 2292
rect 8444 2252 8450 2264
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 8665 2255 8723 2261
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2292 10563 2295
rect 10962 2292 10968 2304
rect 10551 2264 10968 2292
rect 10551 2261 10563 2264
rect 10505 2255 10563 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 13354 2292 13360 2304
rect 13315 2264 13360 2292
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 21910 2292 21916 2304
rect 21871 2264 21916 2292
rect 21910 2252 21916 2264
rect 21968 2252 21974 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 12802 552 12808 604
rect 12860 592 12866 604
rect 13170 592 13176 604
rect 12860 564 13176 592
rect 12860 552 12866 564
rect 13170 552 13176 564
rect 13228 552 13234 604
rect 20438 552 20444 604
rect 20496 592 20502 604
rect 21358 592 21364 604
rect 20496 564 21364 592
rect 20496 552 20502 564
rect 21358 552 21364 564
rect 21416 552 21422 604
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 15292 25440 15344 25492
rect 16580 25440 16632 25492
rect 17960 25440 18012 25492
rect 20076 25440 20128 25492
rect 22744 25440 22796 25492
rect 14372 25304 14424 25356
rect 15568 25304 15620 25356
rect 16672 25347 16724 25356
rect 16672 25313 16681 25347
rect 16681 25313 16715 25347
rect 16715 25313 16724 25347
rect 16672 25304 16724 25313
rect 19340 25304 19392 25356
rect 22008 25347 22060 25356
rect 22008 25313 22017 25347
rect 22017 25313 22051 25347
rect 22051 25313 22060 25347
rect 22008 25304 22060 25313
rect 18420 25236 18472 25288
rect 16396 25100 16448 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 18880 24896 18932 24948
rect 24768 24896 24820 24948
rect 8392 24760 8444 24812
rect 9588 24760 9640 24812
rect 15384 24760 15436 24812
rect 16396 24760 16448 24812
rect 21456 24828 21508 24880
rect 22008 24871 22060 24880
rect 22008 24837 22017 24871
rect 22017 24837 22051 24871
rect 22051 24837 22060 24871
rect 22008 24828 22060 24837
rect 14648 24692 14700 24744
rect 15016 24735 15068 24744
rect 15016 24701 15025 24735
rect 15025 24701 15059 24735
rect 15059 24701 15068 24735
rect 15016 24692 15068 24701
rect 18420 24735 18472 24744
rect 18420 24701 18429 24735
rect 18429 24701 18463 24735
rect 18463 24701 18472 24735
rect 18420 24692 18472 24701
rect 19984 24735 20036 24744
rect 19984 24701 19993 24735
rect 19993 24701 20027 24735
rect 20027 24701 20036 24735
rect 19984 24692 20036 24701
rect 15568 24624 15620 24676
rect 17500 24624 17552 24676
rect 21180 24760 21232 24812
rect 23664 24828 23716 24880
rect 21088 24735 21140 24744
rect 21088 24701 21097 24735
rect 21097 24701 21131 24735
rect 21131 24701 21140 24735
rect 21088 24692 21140 24701
rect 21732 24692 21784 24744
rect 21824 24624 21876 24676
rect 12992 24599 13044 24608
rect 12992 24565 13001 24599
rect 13001 24565 13035 24599
rect 13035 24565 13044 24599
rect 12992 24556 13044 24565
rect 13268 24556 13320 24608
rect 14372 24556 14424 24608
rect 14556 24599 14608 24608
rect 14556 24565 14565 24599
rect 14565 24565 14599 24599
rect 14599 24565 14608 24599
rect 14556 24556 14608 24565
rect 15476 24599 15528 24608
rect 15476 24565 15485 24599
rect 15485 24565 15519 24599
rect 15519 24565 15528 24599
rect 15476 24556 15528 24565
rect 16672 24556 16724 24608
rect 17132 24556 17184 24608
rect 18328 24556 18380 24608
rect 19340 24556 19392 24608
rect 20168 24599 20220 24608
rect 20168 24565 20177 24599
rect 20177 24565 20211 24599
rect 20211 24565 20220 24599
rect 20168 24556 20220 24565
rect 21272 24599 21324 24608
rect 21272 24565 21281 24599
rect 21281 24565 21315 24599
rect 21315 24565 21324 24599
rect 21272 24556 21324 24565
rect 24124 24556 24176 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 12348 24395 12400 24404
rect 12348 24361 12357 24395
rect 12357 24361 12391 24395
rect 12391 24361 12400 24395
rect 12348 24352 12400 24361
rect 15476 24352 15528 24404
rect 16304 24395 16356 24404
rect 16304 24361 16313 24395
rect 16313 24361 16347 24395
rect 16347 24361 16356 24395
rect 16304 24352 16356 24361
rect 20628 24352 20680 24404
rect 23664 24395 23716 24404
rect 23664 24361 23673 24395
rect 23673 24361 23707 24395
rect 23707 24361 23716 24395
rect 23664 24352 23716 24361
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 11520 24216 11572 24268
rect 13820 24259 13872 24268
rect 13820 24225 13829 24259
rect 13829 24225 13863 24259
rect 13863 24225 13872 24259
rect 13820 24216 13872 24225
rect 14464 24216 14516 24268
rect 15384 24216 15436 24268
rect 16028 24216 16080 24268
rect 18052 24216 18104 24268
rect 18604 24216 18656 24268
rect 21272 24259 21324 24268
rect 21272 24225 21281 24259
rect 21281 24225 21315 24259
rect 21315 24225 21324 24259
rect 21272 24216 21324 24225
rect 23848 24216 23900 24268
rect 24124 24216 24176 24268
rect 12716 24148 12768 24200
rect 14004 24191 14056 24200
rect 14004 24157 14013 24191
rect 14013 24157 14047 24191
rect 14047 24157 14056 24191
rect 14004 24148 14056 24157
rect 16120 24148 16172 24200
rect 16488 24148 16540 24200
rect 18420 24191 18472 24200
rect 12348 24012 12400 24064
rect 13452 24055 13504 24064
rect 13452 24021 13461 24055
rect 13461 24021 13495 24055
rect 13495 24021 13504 24055
rect 13452 24012 13504 24021
rect 14556 24080 14608 24132
rect 15016 24080 15068 24132
rect 18420 24157 18429 24191
rect 18429 24157 18463 24191
rect 18463 24157 18472 24191
rect 18420 24148 18472 24157
rect 21180 24148 21232 24200
rect 21824 24148 21876 24200
rect 23572 24148 23624 24200
rect 15660 24012 15712 24064
rect 17776 24055 17828 24064
rect 17776 24021 17785 24055
rect 17785 24021 17819 24055
rect 17819 24021 17828 24055
rect 17776 24012 17828 24021
rect 18972 24055 19024 24064
rect 18972 24021 18981 24055
rect 18981 24021 19015 24055
rect 19015 24021 19024 24055
rect 18972 24012 19024 24021
rect 20904 24055 20956 24064
rect 20904 24021 20913 24055
rect 20913 24021 20947 24055
rect 20947 24021 20956 24055
rect 20904 24012 20956 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 11520 23851 11572 23860
rect 11520 23817 11529 23851
rect 11529 23817 11563 23851
rect 11563 23817 11572 23851
rect 11520 23808 11572 23817
rect 12256 23808 12308 23860
rect 13820 23808 13872 23860
rect 16120 23808 16172 23860
rect 16304 23851 16356 23860
rect 16304 23817 16313 23851
rect 16313 23817 16347 23851
rect 16347 23817 16356 23851
rect 16304 23808 16356 23817
rect 17040 23851 17092 23860
rect 17040 23817 17049 23851
rect 17049 23817 17083 23851
rect 17083 23817 17092 23851
rect 17040 23808 17092 23817
rect 20996 23808 21048 23860
rect 21272 23851 21324 23860
rect 21272 23817 21281 23851
rect 21281 23817 21315 23851
rect 21315 23817 21324 23851
rect 21272 23808 21324 23817
rect 22652 23851 22704 23860
rect 22652 23817 22661 23851
rect 22661 23817 22695 23851
rect 22695 23817 22704 23851
rect 22652 23808 22704 23817
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 15660 23672 15712 23724
rect 24124 23672 24176 23724
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12716 23647 12768 23656
rect 12440 23604 12492 23613
rect 12716 23613 12750 23647
rect 12750 23613 12768 23647
rect 12716 23604 12768 23613
rect 18972 23647 19024 23656
rect 14280 23536 14332 23588
rect 18972 23613 18981 23647
rect 18981 23613 19015 23647
rect 19015 23613 19024 23647
rect 18972 23604 19024 23613
rect 18420 23536 18472 23588
rect 19432 23536 19484 23588
rect 13820 23511 13872 23520
rect 13820 23477 13829 23511
rect 13829 23477 13863 23511
rect 13863 23477 13872 23511
rect 13820 23468 13872 23477
rect 14004 23468 14056 23520
rect 15292 23511 15344 23520
rect 15292 23477 15301 23511
rect 15301 23477 15335 23511
rect 15335 23477 15344 23511
rect 15292 23468 15344 23477
rect 16028 23468 16080 23520
rect 18604 23468 18656 23520
rect 20628 23468 20680 23520
rect 21180 23468 21232 23520
rect 21548 23468 21600 23520
rect 21824 23468 21876 23520
rect 23112 23511 23164 23520
rect 23112 23477 23121 23511
rect 23121 23477 23155 23511
rect 23155 23477 23164 23511
rect 23112 23468 23164 23477
rect 23848 23511 23900 23520
rect 23848 23477 23857 23511
rect 23857 23477 23891 23511
rect 23891 23477 23900 23511
rect 23848 23468 23900 23477
rect 24032 23468 24084 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 13452 23264 13504 23316
rect 15660 23264 15712 23316
rect 16580 23264 16632 23316
rect 17776 23264 17828 23316
rect 18144 23307 18196 23316
rect 18144 23273 18153 23307
rect 18153 23273 18187 23307
rect 18187 23273 18196 23307
rect 18144 23264 18196 23273
rect 19432 23264 19484 23316
rect 21640 23264 21692 23316
rect 23296 23307 23348 23316
rect 23296 23273 23305 23307
rect 23305 23273 23339 23307
rect 23339 23273 23348 23307
rect 23296 23264 23348 23273
rect 23572 23264 23624 23316
rect 15936 23196 15988 23248
rect 16396 23196 16448 23248
rect 24676 23307 24728 23316
rect 24676 23273 24685 23307
rect 24685 23273 24719 23307
rect 24719 23273 24728 23307
rect 24676 23264 24728 23273
rect 23848 23196 23900 23248
rect 11060 23171 11112 23180
rect 11060 23137 11094 23171
rect 11094 23137 11112 23171
rect 11060 23128 11112 23137
rect 12900 23128 12952 23180
rect 13452 23128 13504 23180
rect 18972 23128 19024 23180
rect 21272 23171 21324 23180
rect 21272 23137 21281 23171
rect 21281 23137 21315 23171
rect 21315 23137 21324 23171
rect 21272 23128 21324 23137
rect 24768 23128 24820 23180
rect 10784 23103 10836 23112
rect 10784 23069 10793 23103
rect 10793 23069 10827 23103
rect 10827 23069 10836 23103
rect 10784 23060 10836 23069
rect 13820 23103 13872 23112
rect 13820 23069 13829 23103
rect 13829 23069 13863 23103
rect 13863 23069 13872 23103
rect 13820 23060 13872 23069
rect 14464 23060 14516 23112
rect 15844 23103 15896 23112
rect 15844 23069 15853 23103
rect 15853 23069 15887 23103
rect 15887 23069 15896 23103
rect 15844 23060 15896 23069
rect 20812 23060 20864 23112
rect 22928 23060 22980 23112
rect 12440 22992 12492 23044
rect 20720 22992 20772 23044
rect 11796 22924 11848 22976
rect 13084 22924 13136 22976
rect 14832 22924 14884 22976
rect 15292 22924 15344 22976
rect 22468 22924 22520 22976
rect 24216 22924 24268 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10784 22763 10836 22772
rect 10784 22729 10793 22763
rect 10793 22729 10827 22763
rect 10827 22729 10836 22763
rect 10784 22720 10836 22729
rect 11060 22720 11112 22772
rect 13820 22763 13872 22772
rect 13820 22729 13829 22763
rect 13829 22729 13863 22763
rect 13863 22729 13872 22763
rect 13820 22720 13872 22729
rect 15844 22720 15896 22772
rect 16396 22763 16448 22772
rect 16396 22729 16405 22763
rect 16405 22729 16439 22763
rect 16439 22729 16448 22763
rect 16396 22720 16448 22729
rect 17040 22763 17092 22772
rect 17040 22729 17049 22763
rect 17049 22729 17083 22763
rect 17083 22729 17092 22763
rect 17040 22720 17092 22729
rect 17500 22763 17552 22772
rect 17500 22729 17509 22763
rect 17509 22729 17543 22763
rect 17543 22729 17552 22763
rect 17500 22720 17552 22729
rect 17776 22763 17828 22772
rect 17776 22729 17785 22763
rect 17785 22729 17819 22763
rect 17819 22729 17828 22763
rect 17776 22720 17828 22729
rect 18052 22763 18104 22772
rect 18052 22729 18061 22763
rect 18061 22729 18095 22763
rect 18095 22729 18104 22763
rect 18052 22720 18104 22729
rect 21824 22720 21876 22772
rect 22928 22763 22980 22772
rect 22928 22729 22937 22763
rect 22937 22729 22971 22763
rect 22971 22729 22980 22763
rect 22928 22720 22980 22729
rect 25412 22763 25464 22772
rect 25412 22729 25421 22763
rect 25421 22729 25455 22763
rect 25455 22729 25464 22763
rect 25412 22720 25464 22729
rect 11520 22652 11572 22704
rect 18420 22652 18472 22704
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 15660 22584 15712 22636
rect 18144 22584 18196 22636
rect 23296 22652 23348 22704
rect 21272 22584 21324 22636
rect 23204 22584 23256 22636
rect 23388 22584 23440 22636
rect 24216 22627 24268 22636
rect 24216 22593 24225 22627
rect 24225 22593 24259 22627
rect 24259 22593 24268 22627
rect 24216 22584 24268 22593
rect 17500 22516 17552 22568
rect 18328 22516 18380 22568
rect 12716 22491 12768 22500
rect 12716 22457 12750 22491
rect 12750 22457 12768 22491
rect 12716 22448 12768 22457
rect 14924 22423 14976 22432
rect 14924 22389 14933 22423
rect 14933 22389 14967 22423
rect 14967 22389 14976 22423
rect 14924 22380 14976 22389
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 15384 22423 15436 22432
rect 15384 22389 15393 22423
rect 15393 22389 15427 22423
rect 15427 22389 15436 22423
rect 15384 22380 15436 22389
rect 18972 22380 19024 22432
rect 23848 22516 23900 22568
rect 20260 22448 20312 22500
rect 20720 22380 20772 22432
rect 23296 22380 23348 22432
rect 23664 22423 23716 22432
rect 23664 22389 23673 22423
rect 23673 22389 23707 22423
rect 23707 22389 23716 22423
rect 23664 22380 23716 22389
rect 24768 22423 24820 22432
rect 24768 22389 24777 22423
rect 24777 22389 24811 22423
rect 24811 22389 24820 22423
rect 24768 22380 24820 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 11428 22219 11480 22228
rect 11428 22185 11437 22219
rect 11437 22185 11471 22219
rect 11471 22185 11480 22219
rect 11428 22176 11480 22185
rect 12900 22219 12952 22228
rect 12900 22185 12909 22219
rect 12909 22185 12943 22219
rect 12943 22185 12952 22219
rect 12900 22176 12952 22185
rect 14924 22176 14976 22228
rect 17408 22176 17460 22228
rect 18420 22219 18472 22228
rect 18420 22185 18429 22219
rect 18429 22185 18463 22219
rect 18463 22185 18472 22219
rect 18420 22176 18472 22185
rect 18512 22176 18564 22228
rect 18880 22219 18932 22228
rect 18880 22185 18889 22219
rect 18889 22185 18923 22219
rect 18923 22185 18932 22219
rect 18880 22176 18932 22185
rect 20260 22219 20312 22228
rect 20260 22185 20269 22219
rect 20269 22185 20303 22219
rect 20303 22185 20312 22219
rect 20260 22176 20312 22185
rect 20812 22176 20864 22228
rect 21640 22219 21692 22228
rect 21640 22185 21649 22219
rect 21649 22185 21683 22219
rect 21683 22185 21692 22219
rect 21640 22176 21692 22185
rect 23388 22176 23440 22228
rect 12716 22040 12768 22092
rect 11060 21972 11112 22024
rect 11796 21972 11848 22024
rect 12440 21972 12492 22024
rect 13360 22015 13412 22024
rect 13360 21981 13369 22015
rect 13369 21981 13403 22015
rect 13403 21981 13412 22015
rect 13360 21972 13412 21981
rect 13728 21972 13780 22024
rect 15292 21972 15344 22024
rect 15660 21972 15712 22024
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 15936 22015 15988 22024
rect 15936 21981 15945 22015
rect 15945 21981 15979 22015
rect 15979 21981 15988 22015
rect 15936 21972 15988 21981
rect 16672 21972 16724 22024
rect 17684 21972 17736 22024
rect 18420 21972 18472 22024
rect 16028 21904 16080 21956
rect 22100 22083 22152 22092
rect 22100 22049 22109 22083
rect 22109 22049 22143 22083
rect 22143 22049 22152 22083
rect 23664 22108 23716 22160
rect 23388 22083 23440 22092
rect 22100 22040 22152 22049
rect 22376 21972 22428 22024
rect 23388 22049 23422 22083
rect 23422 22049 23440 22083
rect 23388 22040 23440 22049
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 19156 21904 19208 21956
rect 21088 21904 21140 21956
rect 21916 21904 21968 21956
rect 12348 21836 12400 21888
rect 13452 21836 13504 21888
rect 16396 21879 16448 21888
rect 16396 21845 16405 21879
rect 16405 21845 16439 21879
rect 16439 21845 16448 21879
rect 16396 21836 16448 21845
rect 16948 21879 17000 21888
rect 16948 21845 16957 21879
rect 16957 21845 16991 21879
rect 16991 21845 17000 21879
rect 16948 21836 17000 21845
rect 17592 21836 17644 21888
rect 19524 21879 19576 21888
rect 19524 21845 19533 21879
rect 19533 21845 19567 21879
rect 19567 21845 19576 21879
rect 19524 21836 19576 21845
rect 23296 21836 23348 21888
rect 24216 21836 24268 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 11060 21675 11112 21684
rect 11060 21641 11069 21675
rect 11069 21641 11103 21675
rect 11103 21641 11112 21675
rect 11060 21632 11112 21641
rect 13728 21632 13780 21684
rect 15844 21632 15896 21684
rect 16028 21632 16080 21684
rect 17316 21632 17368 21684
rect 18972 21632 19024 21684
rect 20260 21632 20312 21684
rect 22100 21632 22152 21684
rect 12164 21564 12216 21616
rect 11336 21496 11388 21548
rect 11520 21496 11572 21548
rect 15844 21496 15896 21548
rect 16580 21496 16632 21548
rect 18052 21496 18104 21548
rect 22468 21539 22520 21548
rect 22468 21505 22477 21539
rect 22477 21505 22511 21539
rect 22511 21505 22520 21539
rect 22468 21496 22520 21505
rect 23756 21496 23808 21548
rect 15200 21471 15252 21480
rect 15200 21437 15209 21471
rect 15209 21437 15243 21471
rect 15243 21437 15252 21471
rect 15200 21428 15252 21437
rect 16396 21471 16448 21480
rect 16396 21437 16405 21471
rect 16405 21437 16439 21471
rect 16439 21437 16448 21471
rect 16396 21428 16448 21437
rect 19524 21428 19576 21480
rect 22376 21471 22428 21480
rect 22376 21437 22385 21471
rect 22385 21437 22419 21471
rect 22419 21437 22428 21471
rect 22376 21428 22428 21437
rect 12532 21360 12584 21412
rect 11520 21335 11572 21344
rect 11520 21301 11529 21335
rect 11529 21301 11563 21335
rect 11563 21301 11572 21335
rect 11520 21292 11572 21301
rect 11796 21335 11848 21344
rect 11796 21301 11805 21335
rect 11805 21301 11839 21335
rect 11839 21301 11848 21335
rect 11796 21292 11848 21301
rect 12164 21335 12216 21344
rect 12164 21301 12173 21335
rect 12173 21301 12207 21335
rect 12207 21301 12216 21335
rect 12164 21292 12216 21301
rect 12624 21292 12676 21344
rect 12808 21335 12860 21344
rect 12808 21301 12817 21335
rect 12817 21301 12851 21335
rect 12851 21301 12860 21335
rect 12808 21292 12860 21301
rect 13820 21292 13872 21344
rect 17408 21403 17460 21412
rect 17408 21369 17417 21403
rect 17417 21369 17451 21403
rect 17451 21369 17460 21403
rect 17408 21360 17460 21369
rect 17868 21360 17920 21412
rect 14740 21292 14792 21344
rect 15752 21292 15804 21344
rect 17040 21292 17092 21344
rect 17684 21292 17736 21344
rect 17960 21292 18012 21344
rect 18420 21335 18472 21344
rect 18420 21301 18429 21335
rect 18429 21301 18463 21335
rect 18463 21301 18472 21335
rect 18420 21292 18472 21301
rect 21180 21292 21232 21344
rect 23112 21292 23164 21344
rect 23848 21292 23900 21344
rect 24216 21428 24268 21480
rect 25504 21335 25556 21344
rect 25504 21301 25513 21335
rect 25513 21301 25547 21335
rect 25547 21301 25556 21335
rect 25504 21292 25556 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 13360 21088 13412 21140
rect 14832 21088 14884 21140
rect 15936 21088 15988 21140
rect 16948 21088 17000 21140
rect 17684 21131 17736 21140
rect 17684 21097 17693 21131
rect 17693 21097 17727 21131
rect 17727 21097 17736 21131
rect 17684 21088 17736 21097
rect 18880 21088 18932 21140
rect 22100 21088 22152 21140
rect 23388 21088 23440 21140
rect 23756 21131 23808 21140
rect 23756 21097 23765 21131
rect 23765 21097 23799 21131
rect 23799 21097 23808 21131
rect 23756 21088 23808 21097
rect 15384 21020 15436 21072
rect 17592 21063 17644 21072
rect 17592 21029 17601 21063
rect 17601 21029 17635 21063
rect 17635 21029 17644 21063
rect 17592 21020 17644 21029
rect 1952 20952 2004 21004
rect 11244 20952 11296 21004
rect 11796 20995 11848 21004
rect 11796 20961 11819 20995
rect 11819 20961 11848 20995
rect 15660 20995 15712 21004
rect 11796 20952 11848 20961
rect 15660 20961 15669 20995
rect 15669 20961 15703 20995
rect 15703 20961 15712 20995
rect 15660 20952 15712 20961
rect 11336 20884 11388 20936
rect 15844 20927 15896 20936
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 19524 21020 19576 21072
rect 20720 21020 20772 21072
rect 20904 21020 20956 21072
rect 23112 21020 23164 21072
rect 23572 21020 23624 21072
rect 24032 21020 24084 21072
rect 19156 20995 19208 21004
rect 19156 20961 19165 20995
rect 19165 20961 19199 20995
rect 19199 20961 19208 20995
rect 19156 20952 19208 20961
rect 21824 20995 21876 21004
rect 21824 20961 21833 20995
rect 21833 20961 21867 20995
rect 21867 20961 21876 20995
rect 21824 20952 21876 20961
rect 22100 20995 22152 21004
rect 22100 20961 22134 20995
rect 22134 20961 22152 20995
rect 22100 20952 22152 20961
rect 23480 20952 23532 21004
rect 24676 20995 24728 21004
rect 24676 20961 24685 20995
rect 24685 20961 24719 20995
rect 24719 20961 24728 20995
rect 24676 20952 24728 20961
rect 1584 20859 1636 20868
rect 1584 20825 1593 20859
rect 1593 20825 1627 20859
rect 1627 20825 1636 20859
rect 1584 20816 1636 20825
rect 12808 20816 12860 20868
rect 20260 20884 20312 20936
rect 24216 20884 24268 20936
rect 12900 20791 12952 20800
rect 12900 20757 12909 20791
rect 12909 20757 12943 20791
rect 12943 20757 12952 20791
rect 12900 20748 12952 20757
rect 14832 20748 14884 20800
rect 15292 20791 15344 20800
rect 15292 20757 15301 20791
rect 15301 20757 15335 20791
rect 15335 20757 15344 20791
rect 15292 20748 15344 20757
rect 17040 20791 17092 20800
rect 17040 20757 17049 20791
rect 17049 20757 17083 20791
rect 17083 20757 17092 20791
rect 17040 20748 17092 20757
rect 18420 20748 18472 20800
rect 18788 20791 18840 20800
rect 18788 20757 18797 20791
rect 18797 20757 18831 20791
rect 18831 20757 18840 20791
rect 18788 20748 18840 20757
rect 20444 20748 20496 20800
rect 24124 20791 24176 20800
rect 24124 20757 24133 20791
rect 24133 20757 24167 20791
rect 24167 20757 24176 20791
rect 24124 20748 24176 20757
rect 24216 20748 24268 20800
rect 25504 20884 25556 20936
rect 24952 20748 25004 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 11244 20587 11296 20596
rect 11244 20553 11253 20587
rect 11253 20553 11287 20587
rect 11287 20553 11296 20587
rect 11244 20544 11296 20553
rect 11336 20544 11388 20596
rect 10048 20476 10100 20528
rect 12532 20544 12584 20596
rect 15844 20544 15896 20596
rect 19524 20544 19576 20596
rect 20260 20544 20312 20596
rect 21824 20587 21876 20596
rect 21824 20553 21833 20587
rect 21833 20553 21867 20587
rect 21867 20553 21876 20587
rect 21824 20544 21876 20553
rect 22100 20544 22152 20596
rect 23480 20587 23532 20596
rect 23480 20553 23489 20587
rect 23489 20553 23523 20587
rect 23523 20553 23532 20587
rect 23480 20544 23532 20553
rect 25504 20587 25556 20596
rect 25504 20553 25513 20587
rect 25513 20553 25547 20587
rect 25547 20553 25556 20587
rect 25504 20544 25556 20553
rect 13360 20476 13412 20528
rect 16580 20519 16632 20528
rect 16580 20485 16589 20519
rect 16589 20485 16623 20519
rect 16623 20485 16632 20519
rect 16580 20476 16632 20485
rect 10324 20451 10376 20460
rect 10324 20417 10333 20451
rect 10333 20417 10367 20451
rect 10367 20417 10376 20451
rect 10324 20408 10376 20417
rect 12900 20408 12952 20460
rect 18052 20451 18104 20460
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 20720 20408 20772 20460
rect 25044 20408 25096 20460
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 14648 20383 14700 20392
rect 14648 20349 14657 20383
rect 14657 20349 14691 20383
rect 14691 20349 14700 20383
rect 14648 20340 14700 20349
rect 21640 20340 21692 20392
rect 24124 20340 24176 20392
rect 12532 20272 12584 20324
rect 14832 20272 14884 20324
rect 17040 20272 17092 20324
rect 18696 20272 18748 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 1952 20247 2004 20256
rect 1952 20213 1961 20247
rect 1961 20213 1995 20247
rect 1995 20213 2004 20247
rect 1952 20204 2004 20213
rect 11796 20204 11848 20256
rect 13176 20204 13228 20256
rect 14188 20204 14240 20256
rect 15384 20204 15436 20256
rect 20536 20247 20588 20256
rect 20536 20213 20545 20247
rect 20545 20213 20579 20247
rect 20579 20213 20588 20247
rect 20536 20204 20588 20213
rect 20628 20204 20680 20256
rect 21364 20204 21416 20256
rect 23480 20204 23532 20256
rect 24860 20272 24912 20324
rect 24124 20247 24176 20256
rect 24124 20213 24133 20247
rect 24133 20213 24167 20247
rect 24167 20213 24176 20247
rect 24124 20204 24176 20213
rect 24952 20204 25004 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 12164 20000 12216 20052
rect 17684 20043 17736 20052
rect 17684 20009 17693 20043
rect 17693 20009 17727 20043
rect 17727 20009 17736 20043
rect 17684 20000 17736 20009
rect 18420 20043 18472 20052
rect 18420 20009 18429 20043
rect 18429 20009 18463 20043
rect 18463 20009 18472 20043
rect 18420 20000 18472 20009
rect 19156 20000 19208 20052
rect 22100 20000 22152 20052
rect 24124 20000 24176 20052
rect 12900 19932 12952 19984
rect 15844 19932 15896 19984
rect 19064 19975 19116 19984
rect 19064 19941 19073 19975
rect 19073 19941 19107 19975
rect 19107 19941 19116 19975
rect 19064 19932 19116 19941
rect 20536 19932 20588 19984
rect 21088 19932 21140 19984
rect 25044 19932 25096 19984
rect 10048 19907 10100 19916
rect 10048 19873 10057 19907
rect 10057 19873 10091 19907
rect 10091 19873 10100 19907
rect 10048 19864 10100 19873
rect 10140 19864 10192 19916
rect 12164 19864 12216 19916
rect 13360 19864 13412 19916
rect 14188 19864 14240 19916
rect 14648 19864 14700 19916
rect 16212 19864 16264 19916
rect 18972 19907 19024 19916
rect 18972 19873 18981 19907
rect 18981 19873 19015 19907
rect 19015 19873 19024 19907
rect 18972 19864 19024 19873
rect 20904 19907 20956 19916
rect 20904 19873 20913 19907
rect 20913 19873 20947 19907
rect 20947 19873 20956 19907
rect 20904 19864 20956 19873
rect 19524 19796 19576 19848
rect 23848 19796 23900 19848
rect 20260 19728 20312 19780
rect 1400 19660 1452 19712
rect 11428 19703 11480 19712
rect 11428 19669 11437 19703
rect 11437 19669 11471 19703
rect 11471 19669 11480 19703
rect 11428 19660 11480 19669
rect 11796 19660 11848 19712
rect 12532 19660 12584 19712
rect 16764 19703 16816 19712
rect 16764 19669 16773 19703
rect 16773 19669 16807 19703
rect 16807 19669 16816 19703
rect 16764 19660 16816 19669
rect 18144 19703 18196 19712
rect 18144 19669 18153 19703
rect 18153 19669 18187 19703
rect 18187 19669 18196 19703
rect 18144 19660 18196 19669
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 22008 19660 22060 19712
rect 25320 19703 25372 19712
rect 25320 19669 25329 19703
rect 25329 19669 25363 19703
rect 25363 19669 25372 19703
rect 25320 19660 25372 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 10048 19456 10100 19508
rect 11796 19499 11848 19508
rect 11796 19465 11805 19499
rect 11805 19465 11839 19499
rect 11839 19465 11848 19499
rect 11796 19456 11848 19465
rect 15844 19456 15896 19508
rect 19524 19456 19576 19508
rect 20904 19499 20956 19508
rect 20904 19465 20913 19499
rect 20913 19465 20947 19499
rect 20947 19465 20956 19499
rect 20904 19456 20956 19465
rect 22100 19456 22152 19508
rect 25044 19499 25096 19508
rect 25044 19465 25053 19499
rect 25053 19465 25087 19499
rect 25087 19465 25096 19499
rect 25044 19456 25096 19465
rect 18972 19388 19024 19440
rect 10140 19320 10192 19372
rect 10876 19363 10928 19372
rect 10876 19329 10885 19363
rect 10885 19329 10919 19363
rect 10919 19329 10928 19363
rect 10876 19320 10928 19329
rect 11428 19320 11480 19372
rect 12440 19320 12492 19372
rect 12900 19320 12952 19372
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 9680 19252 9732 19304
rect 18144 19252 18196 19304
rect 19248 19252 19300 19304
rect 21180 19388 21232 19440
rect 20260 19363 20312 19372
rect 20260 19329 20269 19363
rect 20269 19329 20303 19363
rect 20303 19329 20312 19363
rect 20260 19320 20312 19329
rect 20904 19320 20956 19372
rect 24584 19363 24636 19372
rect 21180 19252 21232 19304
rect 22008 19252 22060 19304
rect 24584 19329 24593 19363
rect 24593 19329 24627 19363
rect 24627 19329 24636 19363
rect 24584 19320 24636 19329
rect 25320 19320 25372 19372
rect 23940 19252 23992 19304
rect 10140 19116 10192 19168
rect 10784 19116 10836 19168
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12440 19116 12492 19125
rect 15752 19184 15804 19236
rect 17132 19184 17184 19236
rect 13176 19116 13228 19168
rect 14188 19116 14240 19168
rect 14832 19116 14884 19168
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 16948 19116 17000 19168
rect 23848 19184 23900 19236
rect 18512 19159 18564 19168
rect 18512 19125 18521 19159
rect 18521 19125 18555 19159
rect 18555 19125 18564 19159
rect 18512 19116 18564 19125
rect 19524 19159 19576 19168
rect 19524 19125 19533 19159
rect 19533 19125 19567 19159
rect 19567 19125 19576 19159
rect 19524 19116 19576 19125
rect 20168 19159 20220 19168
rect 20168 19125 20177 19159
rect 20177 19125 20211 19159
rect 20211 19125 20220 19159
rect 20168 19116 20220 19125
rect 20628 19116 20680 19168
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 21732 19159 21784 19168
rect 21732 19125 21741 19159
rect 21741 19125 21775 19159
rect 21775 19125 21784 19159
rect 21732 19116 21784 19125
rect 22284 19116 22336 19168
rect 23940 19159 23992 19168
rect 23940 19125 23949 19159
rect 23949 19125 23983 19159
rect 23983 19125 23992 19159
rect 23940 19116 23992 19125
rect 24124 19252 24176 19304
rect 25504 19295 25556 19304
rect 25504 19261 25513 19295
rect 25513 19261 25547 19295
rect 25547 19261 25556 19295
rect 25504 19252 25556 19261
rect 24216 19184 24268 19236
rect 24124 19116 24176 19168
rect 25688 19159 25740 19168
rect 25688 19125 25697 19159
rect 25697 19125 25731 19159
rect 25731 19125 25740 19159
rect 25688 19116 25740 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 12900 18955 12952 18964
rect 12900 18921 12909 18955
rect 12909 18921 12943 18955
rect 12943 18921 12952 18955
rect 12900 18912 12952 18921
rect 13728 18912 13780 18964
rect 13912 18912 13964 18964
rect 14096 18955 14148 18964
rect 14096 18921 14105 18955
rect 14105 18921 14139 18955
rect 14139 18921 14148 18955
rect 14096 18912 14148 18921
rect 15292 18912 15344 18964
rect 18972 18912 19024 18964
rect 21180 18955 21232 18964
rect 21180 18921 21189 18955
rect 21189 18921 21223 18955
rect 21223 18921 21232 18955
rect 21180 18912 21232 18921
rect 21548 18955 21600 18964
rect 21548 18921 21557 18955
rect 21557 18921 21591 18955
rect 21591 18921 21600 18955
rect 21548 18912 21600 18921
rect 21732 18912 21784 18964
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 14740 18844 14792 18896
rect 16672 18844 16724 18896
rect 19064 18887 19116 18896
rect 19064 18853 19073 18887
rect 19073 18853 19107 18887
rect 19107 18853 19116 18887
rect 19064 18844 19116 18853
rect 24216 18844 24268 18896
rect 24584 18844 24636 18896
rect 10324 18776 10376 18828
rect 10876 18819 10928 18828
rect 10876 18785 10899 18819
rect 10899 18785 10928 18819
rect 10876 18776 10928 18785
rect 17684 18776 17736 18828
rect 19800 18819 19852 18828
rect 19800 18785 19809 18819
rect 19809 18785 19843 18819
rect 19843 18785 19852 18819
rect 19800 18776 19852 18785
rect 22284 18819 22336 18828
rect 22284 18785 22293 18819
rect 22293 18785 22327 18819
rect 22327 18785 22336 18819
rect 22284 18776 22336 18785
rect 10048 18708 10100 18760
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 10600 18708 10652 18717
rect 14188 18751 14240 18760
rect 14188 18717 14197 18751
rect 14197 18717 14231 18751
rect 14231 18717 14240 18751
rect 16028 18751 16080 18760
rect 14188 18708 14240 18717
rect 16028 18717 16037 18751
rect 16037 18717 16071 18751
rect 16071 18717 16080 18751
rect 16028 18708 16080 18717
rect 16948 18708 17000 18760
rect 21180 18708 21232 18760
rect 21640 18751 21692 18760
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 21088 18640 21140 18692
rect 23388 18708 23440 18760
rect 23848 18751 23900 18760
rect 23848 18717 23857 18751
rect 23857 18717 23891 18751
rect 23891 18717 23900 18751
rect 23848 18708 23900 18717
rect 22928 18640 22980 18692
rect 23480 18640 23532 18692
rect 10784 18572 10836 18624
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 14004 18572 14056 18624
rect 14648 18615 14700 18624
rect 14648 18581 14657 18615
rect 14657 18581 14691 18615
rect 14691 18581 14700 18615
rect 14648 18572 14700 18581
rect 15384 18615 15436 18624
rect 15384 18581 15393 18615
rect 15393 18581 15427 18615
rect 15427 18581 15436 18615
rect 15384 18572 15436 18581
rect 16580 18572 16632 18624
rect 19984 18615 20036 18624
rect 19984 18581 19993 18615
rect 19993 18581 20027 18615
rect 20027 18581 20036 18615
rect 19984 18572 20036 18581
rect 25228 18615 25280 18624
rect 25228 18581 25237 18615
rect 25237 18581 25271 18615
rect 25271 18581 25280 18615
rect 25228 18572 25280 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 10600 18411 10652 18420
rect 10600 18377 10609 18411
rect 10609 18377 10643 18411
rect 10643 18377 10652 18411
rect 10600 18368 10652 18377
rect 13912 18368 13964 18420
rect 15752 18411 15804 18420
rect 15752 18377 15761 18411
rect 15761 18377 15795 18411
rect 15795 18377 15804 18411
rect 15752 18368 15804 18377
rect 16028 18368 16080 18420
rect 16764 18368 16816 18420
rect 17684 18411 17736 18420
rect 17684 18377 17693 18411
rect 17693 18377 17727 18411
rect 17727 18377 17736 18411
rect 17684 18368 17736 18377
rect 18604 18411 18656 18420
rect 18604 18377 18613 18411
rect 18613 18377 18647 18411
rect 18647 18377 18656 18411
rect 18604 18368 18656 18377
rect 20444 18411 20496 18420
rect 20444 18377 20453 18411
rect 20453 18377 20487 18411
rect 20487 18377 20496 18411
rect 20444 18368 20496 18377
rect 21732 18368 21784 18420
rect 23204 18368 23256 18420
rect 11152 18300 11204 18352
rect 10140 18232 10192 18284
rect 14096 18300 14148 18352
rect 16672 18343 16724 18352
rect 16672 18309 16681 18343
rect 16681 18309 16715 18343
rect 16715 18309 16724 18343
rect 16672 18300 16724 18309
rect 11428 18275 11480 18284
rect 11428 18241 11437 18275
rect 11437 18241 11471 18275
rect 11471 18241 11480 18275
rect 11428 18232 11480 18241
rect 11980 18232 12032 18284
rect 14188 18232 14240 18284
rect 22100 18232 22152 18284
rect 22284 18232 22336 18284
rect 23848 18368 23900 18420
rect 24768 18232 24820 18284
rect 25228 18368 25280 18420
rect 13360 18207 13412 18216
rect 13360 18173 13369 18207
rect 13369 18173 13403 18207
rect 13403 18173 13412 18207
rect 13360 18164 13412 18173
rect 14004 18164 14056 18216
rect 14648 18207 14700 18216
rect 14648 18173 14682 18207
rect 14682 18173 14700 18207
rect 14648 18164 14700 18173
rect 16580 18164 16632 18216
rect 18604 18164 18656 18216
rect 14740 18096 14792 18148
rect 16948 18096 17000 18148
rect 21548 18164 21600 18216
rect 23664 18164 23716 18216
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 19340 18139 19392 18148
rect 19340 18105 19374 18139
rect 19374 18105 19392 18139
rect 19340 18096 19392 18105
rect 21364 18096 21416 18148
rect 22560 18139 22612 18148
rect 22560 18105 22569 18139
rect 22569 18105 22603 18139
rect 22603 18105 22612 18139
rect 22560 18096 22612 18105
rect 23572 18096 23624 18148
rect 23848 18096 23900 18148
rect 11060 18028 11112 18080
rect 13544 18071 13596 18080
rect 13544 18037 13553 18071
rect 13553 18037 13587 18071
rect 13587 18037 13596 18071
rect 13544 18028 13596 18037
rect 17224 18028 17276 18080
rect 18052 18028 18104 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 21272 18071 21324 18080
rect 21272 18037 21281 18071
rect 21281 18037 21315 18071
rect 21315 18037 21324 18071
rect 21272 18028 21324 18037
rect 23664 18071 23716 18080
rect 23664 18037 23673 18071
rect 23673 18037 23707 18071
rect 23707 18037 23716 18071
rect 23664 18028 23716 18037
rect 25412 18071 25464 18080
rect 25412 18037 25421 18071
rect 25421 18037 25455 18071
rect 25455 18037 25464 18071
rect 25412 18028 25464 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 13360 17867 13412 17876
rect 13360 17833 13369 17867
rect 13369 17833 13403 17867
rect 13403 17833 13412 17867
rect 13360 17824 13412 17833
rect 20076 17824 20128 17876
rect 20352 17867 20404 17876
rect 20352 17833 20361 17867
rect 20361 17833 20395 17867
rect 20395 17833 20404 17867
rect 20352 17824 20404 17833
rect 20720 17824 20772 17876
rect 20996 17824 21048 17876
rect 23664 17867 23716 17876
rect 23664 17833 23673 17867
rect 23673 17833 23707 17867
rect 23707 17833 23716 17867
rect 23664 17824 23716 17833
rect 24216 17867 24268 17876
rect 24216 17833 24225 17867
rect 24225 17833 24259 17867
rect 24259 17833 24268 17867
rect 24216 17824 24268 17833
rect 11428 17799 11480 17808
rect 11428 17765 11462 17799
rect 11462 17765 11480 17799
rect 11428 17756 11480 17765
rect 14004 17799 14056 17808
rect 14004 17765 14013 17799
rect 14013 17765 14047 17799
rect 14047 17765 14056 17799
rect 14004 17756 14056 17765
rect 14280 17756 14332 17808
rect 14740 17799 14792 17808
rect 14740 17765 14749 17799
rect 14749 17765 14783 17799
rect 14783 17765 14792 17799
rect 14740 17756 14792 17765
rect 17408 17756 17460 17808
rect 23296 17756 23348 17808
rect 20 17688 72 17740
rect 9588 17688 9640 17740
rect 10692 17688 10744 17740
rect 11796 17688 11848 17740
rect 14648 17688 14700 17740
rect 15660 17731 15712 17740
rect 14832 17620 14884 17672
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 19800 17731 19852 17740
rect 19800 17697 19809 17731
rect 19809 17697 19843 17731
rect 19843 17697 19852 17731
rect 19800 17688 19852 17697
rect 20720 17688 20772 17740
rect 20904 17688 20956 17740
rect 21364 17688 21416 17740
rect 23572 17731 23624 17740
rect 23572 17697 23581 17731
rect 23581 17697 23615 17731
rect 23615 17697 23624 17731
rect 23572 17688 23624 17697
rect 25596 17688 25648 17740
rect 16304 17663 16356 17672
rect 16304 17629 16313 17663
rect 16313 17629 16347 17663
rect 16347 17629 16356 17663
rect 16304 17620 16356 17629
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 23296 17620 23348 17672
rect 23204 17595 23256 17604
rect 23204 17561 23213 17595
rect 23213 17561 23247 17595
rect 23247 17561 23256 17595
rect 23204 17552 23256 17561
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 15292 17527 15344 17536
rect 15292 17493 15301 17527
rect 15301 17493 15335 17527
rect 15335 17493 15344 17527
rect 15292 17484 15344 17493
rect 18328 17527 18380 17536
rect 18328 17493 18337 17527
rect 18337 17493 18371 17527
rect 18371 17493 18380 17527
rect 18328 17484 18380 17493
rect 19156 17527 19208 17536
rect 19156 17493 19165 17527
rect 19165 17493 19199 17527
rect 19199 17493 19208 17527
rect 19156 17484 19208 17493
rect 19340 17484 19392 17536
rect 21088 17484 21140 17536
rect 22100 17484 22152 17536
rect 24952 17527 25004 17536
rect 24952 17493 24961 17527
rect 24961 17493 24995 17527
rect 24995 17493 25004 17527
rect 24952 17484 25004 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 16304 17323 16356 17332
rect 16304 17289 16313 17323
rect 16313 17289 16347 17323
rect 16347 17289 16356 17323
rect 16304 17280 16356 17289
rect 22560 17323 22612 17332
rect 22560 17289 22569 17323
rect 22569 17289 22603 17323
rect 22603 17289 22612 17323
rect 22560 17280 22612 17289
rect 23296 17280 23348 17332
rect 25596 17323 25648 17332
rect 25596 17289 25605 17323
rect 25605 17289 25639 17323
rect 25639 17289 25648 17323
rect 25596 17280 25648 17289
rect 11244 17144 11296 17196
rect 11428 17187 11480 17196
rect 11428 17153 11437 17187
rect 11437 17153 11471 17187
rect 11471 17153 11480 17187
rect 11428 17144 11480 17153
rect 23664 17212 23716 17264
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 10968 17076 11020 17128
rect 11336 17008 11388 17060
rect 11060 16940 11112 16992
rect 12532 17076 12584 17128
rect 16028 17076 16080 17128
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 14832 17008 14884 17060
rect 14280 16940 14332 16992
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 20904 17076 20956 17128
rect 24768 17076 24820 17128
rect 19064 17008 19116 17060
rect 19340 17008 19392 17060
rect 21364 17008 21416 17060
rect 22560 17008 22612 17060
rect 16948 16940 17000 16949
rect 19156 16940 19208 16992
rect 21180 16983 21232 16992
rect 21180 16949 21189 16983
rect 21189 16949 21223 16983
rect 21223 16949 21232 16983
rect 21180 16940 21232 16949
rect 21640 16983 21692 16992
rect 21640 16949 21649 16983
rect 21649 16949 21683 16983
rect 21683 16949 21692 16983
rect 21640 16940 21692 16949
rect 23020 16983 23072 16992
rect 23020 16949 23029 16983
rect 23029 16949 23063 16983
rect 23063 16949 23072 16983
rect 23020 16940 23072 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 11244 16779 11296 16788
rect 11244 16745 11253 16779
rect 11253 16745 11287 16779
rect 11287 16745 11296 16779
rect 11244 16736 11296 16745
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 14004 16736 14056 16788
rect 14832 16736 14884 16788
rect 15660 16736 15712 16788
rect 15844 16736 15896 16788
rect 11060 16668 11112 16720
rect 14648 16711 14700 16720
rect 11336 16600 11388 16652
rect 14648 16677 14657 16711
rect 14657 16677 14691 16711
rect 14691 16677 14700 16711
rect 14648 16668 14700 16677
rect 15292 16668 15344 16720
rect 11152 16532 11204 16584
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 11980 16575 12032 16584
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 14648 16532 14700 16584
rect 14740 16532 14792 16584
rect 19064 16736 19116 16788
rect 19524 16736 19576 16788
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 20996 16736 21048 16788
rect 22284 16779 22336 16788
rect 22284 16745 22293 16779
rect 22293 16745 22327 16779
rect 22327 16745 22336 16779
rect 22284 16736 22336 16745
rect 23572 16736 23624 16788
rect 23664 16736 23716 16788
rect 24124 16736 24176 16788
rect 21088 16668 21140 16720
rect 23204 16711 23256 16720
rect 23204 16677 23213 16711
rect 23213 16677 23247 16711
rect 23247 16677 23256 16711
rect 23204 16668 23256 16677
rect 15752 16532 15804 16584
rect 16948 16600 17000 16652
rect 17132 16643 17184 16652
rect 17132 16609 17166 16643
rect 17166 16609 17184 16643
rect 17132 16600 17184 16609
rect 18328 16600 18380 16652
rect 20904 16643 20956 16652
rect 20904 16609 20913 16643
rect 20913 16609 20947 16643
rect 20947 16609 20956 16643
rect 20904 16600 20956 16609
rect 23480 16600 23532 16652
rect 24216 16600 24268 16652
rect 16764 16532 16816 16584
rect 23664 16532 23716 16584
rect 24032 16532 24084 16584
rect 24768 16736 24820 16788
rect 25228 16779 25280 16788
rect 25228 16745 25237 16779
rect 25237 16745 25271 16779
rect 25271 16745 25280 16779
rect 25228 16736 25280 16745
rect 25044 16643 25096 16652
rect 25044 16609 25053 16643
rect 25053 16609 25087 16643
rect 25087 16609 25096 16643
rect 25044 16600 25096 16609
rect 14280 16464 14332 16516
rect 12440 16396 12492 16448
rect 18236 16439 18288 16448
rect 18236 16405 18245 16439
rect 18245 16405 18279 16439
rect 18279 16405 18288 16439
rect 18236 16396 18288 16405
rect 21088 16396 21140 16448
rect 21824 16396 21876 16448
rect 23020 16396 23072 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 11060 16192 11112 16244
rect 11980 16192 12032 16244
rect 14740 16192 14792 16244
rect 15752 16235 15804 16244
rect 15752 16201 15761 16235
rect 15761 16201 15795 16235
rect 15795 16201 15804 16235
rect 15752 16192 15804 16201
rect 19156 16192 19208 16244
rect 20904 16192 20956 16244
rect 21916 16192 21968 16244
rect 24032 16192 24084 16244
rect 24216 16235 24268 16244
rect 24216 16201 24225 16235
rect 24225 16201 24259 16235
rect 24259 16201 24268 16235
rect 24216 16192 24268 16201
rect 25044 16192 25096 16244
rect 11796 16124 11848 16176
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 14832 16056 14884 16108
rect 17132 16124 17184 16176
rect 19156 16099 19208 16108
rect 19156 16065 19165 16099
rect 19165 16065 19199 16099
rect 19199 16065 19208 16099
rect 19156 16056 19208 16065
rect 21088 16056 21140 16108
rect 21824 16056 21876 16108
rect 22284 16099 22336 16108
rect 22284 16065 22293 16099
rect 22293 16065 22327 16099
rect 22327 16065 22336 16099
rect 22284 16056 22336 16065
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 14648 15988 14700 16040
rect 16764 16031 16816 16040
rect 16764 15997 16773 16031
rect 16773 15997 16807 16031
rect 16807 15997 16816 16031
rect 16764 15988 16816 15997
rect 19248 15988 19300 16040
rect 16120 15920 16172 15972
rect 18696 15920 18748 15972
rect 21180 15988 21232 16040
rect 24584 16031 24636 16040
rect 24584 15997 24593 16031
rect 24593 15997 24627 16031
rect 24627 15997 24636 16031
rect 24584 15988 24636 15997
rect 13728 15852 13780 15904
rect 14188 15852 14240 15904
rect 15200 15852 15252 15904
rect 16396 15895 16448 15904
rect 16396 15861 16405 15895
rect 16405 15861 16439 15895
rect 16439 15861 16448 15895
rect 16396 15852 16448 15861
rect 16948 15852 17000 15904
rect 19156 15852 19208 15904
rect 20076 15895 20128 15904
rect 20076 15861 20085 15895
rect 20085 15861 20119 15895
rect 20119 15861 20128 15895
rect 20076 15852 20128 15861
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 20536 15852 20588 15861
rect 23664 15852 23716 15904
rect 24768 15895 24820 15904
rect 24768 15861 24777 15895
rect 24777 15861 24811 15895
rect 24811 15861 24820 15895
rect 24768 15852 24820 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 14648 15691 14700 15700
rect 14648 15657 14657 15691
rect 14657 15657 14691 15691
rect 14691 15657 14700 15691
rect 14648 15648 14700 15657
rect 15108 15691 15160 15700
rect 15108 15657 15117 15691
rect 15117 15657 15151 15691
rect 15151 15657 15160 15691
rect 15108 15648 15160 15657
rect 17040 15691 17092 15700
rect 17040 15657 17049 15691
rect 17049 15657 17083 15691
rect 17083 15657 17092 15691
rect 17040 15648 17092 15657
rect 19248 15648 19300 15700
rect 20536 15648 20588 15700
rect 21180 15648 21232 15700
rect 21824 15691 21876 15700
rect 21824 15657 21833 15691
rect 21833 15657 21867 15691
rect 21867 15657 21876 15691
rect 21824 15648 21876 15657
rect 23020 15648 23072 15700
rect 14280 15512 14332 15564
rect 15752 15512 15804 15564
rect 14832 15444 14884 15496
rect 16396 15512 16448 15564
rect 17408 15555 17460 15564
rect 17408 15521 17442 15555
rect 17442 15521 17460 15555
rect 17408 15512 17460 15521
rect 21364 15512 21416 15564
rect 21916 15555 21968 15564
rect 21916 15521 21925 15555
rect 21925 15521 21959 15555
rect 21959 15521 21968 15555
rect 21916 15512 21968 15521
rect 22192 15555 22244 15564
rect 22192 15521 22226 15555
rect 22226 15521 22244 15555
rect 24584 15555 24636 15564
rect 22192 15512 22244 15521
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 16212 15487 16264 15496
rect 16212 15453 16221 15487
rect 16221 15453 16255 15487
rect 16255 15453 16264 15487
rect 16212 15444 16264 15453
rect 16948 15444 17000 15496
rect 19432 15444 19484 15496
rect 15108 15376 15160 15428
rect 24768 15419 24820 15428
rect 24768 15385 24777 15419
rect 24777 15385 24811 15419
rect 24811 15385 24820 15419
rect 24768 15376 24820 15385
rect 15292 15308 15344 15360
rect 16488 15308 16540 15360
rect 18604 15308 18656 15360
rect 21548 15308 21600 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 14280 15147 14332 15156
rect 14280 15113 14289 15147
rect 14289 15113 14323 15147
rect 14323 15113 14332 15147
rect 14280 15104 14332 15113
rect 14832 15104 14884 15156
rect 15752 15147 15804 15156
rect 15752 15113 15761 15147
rect 15761 15113 15795 15147
rect 15795 15113 15804 15147
rect 15752 15104 15804 15113
rect 16396 15104 16448 15156
rect 20812 15147 20864 15156
rect 20812 15113 20821 15147
rect 20821 15113 20855 15147
rect 20855 15113 20864 15147
rect 20812 15104 20864 15113
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 22192 15104 22244 15156
rect 22744 15147 22796 15156
rect 22744 15113 22753 15147
rect 22753 15113 22787 15147
rect 22787 15113 22796 15147
rect 22744 15104 22796 15113
rect 24676 15104 24728 15156
rect 16580 14968 16632 15020
rect 12624 14900 12676 14952
rect 17408 14900 17460 14952
rect 16212 14832 16264 14884
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 15200 14807 15252 14816
rect 15200 14773 15209 14807
rect 15209 14773 15243 14807
rect 15243 14773 15252 14807
rect 15200 14764 15252 14773
rect 16580 14807 16632 14816
rect 16580 14773 16589 14807
rect 16589 14773 16623 14807
rect 16623 14773 16632 14807
rect 16580 14764 16632 14773
rect 16948 14764 17000 14816
rect 18604 14900 18656 14952
rect 20812 14900 20864 14952
rect 24584 14943 24636 14952
rect 21364 14832 21416 14884
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 19984 14764 20036 14816
rect 20904 14764 20956 14816
rect 21916 14764 21968 14816
rect 22744 14764 22796 14816
rect 23112 14807 23164 14816
rect 23112 14773 23121 14807
rect 23121 14773 23155 14807
rect 23155 14773 23164 14807
rect 23112 14764 23164 14773
rect 24768 14807 24820 14816
rect 24768 14773 24777 14807
rect 24777 14773 24811 14807
rect 24811 14773 24820 14807
rect 24768 14764 24820 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 15200 14560 15252 14612
rect 16120 14560 16172 14612
rect 17408 14603 17460 14612
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 18604 14603 18656 14612
rect 18604 14569 18613 14603
rect 18613 14569 18647 14603
rect 18647 14569 18656 14603
rect 18604 14560 18656 14569
rect 19064 14603 19116 14612
rect 19064 14569 19073 14603
rect 19073 14569 19107 14603
rect 19107 14569 19116 14603
rect 19064 14560 19116 14569
rect 19432 14603 19484 14612
rect 19432 14569 19441 14603
rect 19441 14569 19475 14603
rect 19475 14569 19484 14603
rect 19432 14560 19484 14569
rect 24860 14560 24912 14612
rect 15292 14492 15344 14544
rect 16212 14492 16264 14544
rect 16396 14492 16448 14544
rect 20996 14492 21048 14544
rect 13084 14467 13136 14476
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 13176 14424 13228 14476
rect 14648 14424 14700 14476
rect 16856 14424 16908 14476
rect 20904 14467 20956 14476
rect 20904 14433 20913 14467
rect 20913 14433 20947 14467
rect 20947 14433 20956 14467
rect 20904 14424 20956 14433
rect 23296 14424 23348 14476
rect 25780 14424 25832 14476
rect 18052 14356 18104 14408
rect 22744 14399 22796 14408
rect 14280 14331 14332 14340
rect 14280 14297 14289 14331
rect 14289 14297 14323 14331
rect 14323 14297 14332 14331
rect 14280 14288 14332 14297
rect 19340 14288 19392 14340
rect 22744 14365 22753 14399
rect 22753 14365 22787 14399
rect 22787 14365 22796 14399
rect 22744 14356 22796 14365
rect 19984 14288 20036 14340
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 21088 14263 21140 14272
rect 21088 14229 21097 14263
rect 21097 14229 21131 14263
rect 21131 14229 21140 14263
rect 21088 14220 21140 14229
rect 24124 14263 24176 14272
rect 24124 14229 24133 14263
rect 24133 14229 24167 14263
rect 24167 14229 24176 14263
rect 24124 14220 24176 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 13084 14059 13136 14068
rect 13084 14025 13093 14059
rect 13093 14025 13127 14059
rect 13127 14025 13136 14059
rect 13084 14016 13136 14025
rect 14648 14059 14700 14068
rect 14648 14025 14657 14059
rect 14657 14025 14691 14059
rect 14691 14025 14700 14059
rect 14648 14016 14700 14025
rect 16580 14016 16632 14068
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 19432 14016 19484 14068
rect 20904 14016 20956 14068
rect 22744 14016 22796 14068
rect 23112 14016 23164 14068
rect 25780 14059 25832 14068
rect 25780 14025 25789 14059
rect 25789 14025 25823 14059
rect 25823 14025 25832 14059
rect 25780 14016 25832 14025
rect 14556 13948 14608 14000
rect 22284 13948 22336 14000
rect 24124 13948 24176 14000
rect 25412 13991 25464 14000
rect 16396 13923 16448 13932
rect 16396 13889 16405 13923
rect 16405 13889 16439 13923
rect 16439 13889 16448 13923
rect 16396 13880 16448 13889
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 19340 13880 19392 13932
rect 25412 13957 25421 13991
rect 25421 13957 25455 13991
rect 25455 13957 25464 13991
rect 25412 13948 25464 13957
rect 13820 13812 13872 13864
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 16120 13855 16172 13864
rect 16120 13821 16129 13855
rect 16129 13821 16163 13855
rect 16163 13821 16172 13855
rect 16120 13812 16172 13821
rect 16948 13812 17000 13864
rect 17960 13812 18012 13864
rect 19064 13812 19116 13864
rect 25044 13923 25096 13932
rect 25044 13889 25053 13923
rect 25053 13889 25087 13923
rect 25087 13889 25096 13923
rect 25044 13880 25096 13889
rect 11244 13744 11296 13796
rect 22744 13812 22796 13864
rect 23296 13744 23348 13796
rect 15936 13676 15988 13728
rect 16396 13676 16448 13728
rect 19984 13676 20036 13728
rect 20996 13719 21048 13728
rect 20996 13685 21005 13719
rect 21005 13685 21039 13719
rect 21039 13685 21048 13719
rect 20996 13676 21048 13685
rect 22560 13719 22612 13728
rect 22560 13685 22569 13719
rect 22569 13685 22603 13719
rect 22603 13685 22612 13719
rect 22560 13676 22612 13685
rect 24032 13719 24084 13728
rect 24032 13685 24041 13719
rect 24041 13685 24075 13719
rect 24075 13685 24084 13719
rect 24032 13676 24084 13685
rect 24124 13719 24176 13728
rect 24124 13685 24133 13719
rect 24133 13685 24167 13719
rect 24167 13685 24176 13719
rect 24124 13676 24176 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 13912 13472 13964 13524
rect 14832 13472 14884 13524
rect 17960 13472 18012 13524
rect 19340 13472 19392 13524
rect 19524 13472 19576 13524
rect 20168 13472 20220 13524
rect 22192 13515 22244 13524
rect 22192 13481 22201 13515
rect 22201 13481 22235 13515
rect 22235 13481 22244 13515
rect 22192 13472 22244 13481
rect 22560 13472 22612 13524
rect 23020 13515 23072 13524
rect 23020 13481 23029 13515
rect 23029 13481 23063 13515
rect 23063 13481 23072 13515
rect 23020 13472 23072 13481
rect 23112 13515 23164 13524
rect 23112 13481 23121 13515
rect 23121 13481 23155 13515
rect 23155 13481 23164 13515
rect 23112 13472 23164 13481
rect 23848 13472 23900 13524
rect 24124 13472 24176 13524
rect 24216 13472 24268 13524
rect 13544 13404 13596 13456
rect 14464 13404 14516 13456
rect 16580 13447 16632 13456
rect 16580 13413 16589 13447
rect 16589 13413 16623 13447
rect 16623 13413 16632 13447
rect 16580 13404 16632 13413
rect 17592 13404 17644 13456
rect 13912 13336 13964 13388
rect 14188 13336 14240 13388
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 17776 13268 17828 13320
rect 18880 13268 18932 13320
rect 20076 13336 20128 13388
rect 21088 13336 21140 13388
rect 24584 13379 24636 13388
rect 24584 13345 24593 13379
rect 24593 13345 24627 13379
rect 24627 13345 24636 13379
rect 24584 13336 24636 13345
rect 19800 13311 19852 13320
rect 19800 13277 19809 13311
rect 19809 13277 19843 13311
rect 19843 13277 19852 13311
rect 21364 13311 21416 13320
rect 19800 13268 19852 13277
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 23296 13311 23348 13320
rect 16672 13200 16724 13252
rect 19524 13200 19576 13252
rect 20996 13200 21048 13252
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 21548 13200 21600 13252
rect 24032 13243 24084 13252
rect 24032 13209 24041 13243
rect 24041 13209 24075 13243
rect 24075 13209 24084 13243
rect 24032 13200 24084 13209
rect 14280 13132 14332 13184
rect 14464 13132 14516 13184
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 20904 13175 20956 13184
rect 20904 13141 20913 13175
rect 20913 13141 20947 13175
rect 20947 13141 20956 13175
rect 20904 13132 20956 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 14188 12928 14240 12980
rect 15844 12928 15896 12980
rect 16212 12928 16264 12980
rect 16304 12928 16356 12980
rect 19800 12928 19852 12980
rect 20168 12971 20220 12980
rect 20168 12937 20177 12971
rect 20177 12937 20211 12971
rect 20211 12937 20220 12971
rect 20168 12928 20220 12937
rect 21180 12928 21232 12980
rect 21364 12928 21416 12980
rect 23020 12971 23072 12980
rect 23020 12937 23029 12971
rect 23029 12937 23063 12971
rect 23063 12937 23072 12971
rect 23020 12928 23072 12937
rect 24676 12928 24728 12980
rect 11980 12860 12032 12912
rect 13912 12860 13964 12912
rect 18972 12860 19024 12912
rect 18880 12835 18932 12844
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 14464 12767 14516 12776
rect 14464 12733 14498 12767
rect 14498 12733 14516 12767
rect 14464 12724 14516 12733
rect 16672 12767 16724 12776
rect 16672 12733 16681 12767
rect 16681 12733 16715 12767
rect 16715 12733 16724 12767
rect 16672 12724 16724 12733
rect 17776 12724 17828 12776
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 19340 12792 19392 12844
rect 21732 12792 21784 12844
rect 23480 12860 23532 12912
rect 22468 12792 22520 12844
rect 23112 12792 23164 12844
rect 19524 12767 19576 12776
rect 13912 12656 13964 12708
rect 14832 12656 14884 12708
rect 18328 12656 18380 12708
rect 19524 12733 19533 12767
rect 19533 12733 19567 12767
rect 19567 12733 19576 12767
rect 19524 12724 19576 12733
rect 20720 12724 20772 12776
rect 20904 12656 20956 12708
rect 21088 12724 21140 12776
rect 22192 12767 22244 12776
rect 22192 12733 22201 12767
rect 22201 12733 22235 12767
rect 22235 12733 22244 12767
rect 22192 12724 22244 12733
rect 23756 12724 23808 12776
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 15476 12588 15528 12640
rect 16580 12631 16632 12640
rect 16580 12597 16589 12631
rect 16589 12597 16623 12631
rect 16623 12597 16632 12631
rect 16580 12588 16632 12597
rect 19156 12588 19208 12640
rect 20536 12588 20588 12640
rect 20996 12631 21048 12640
rect 20996 12597 21005 12631
rect 21005 12597 21039 12631
rect 21039 12597 21048 12631
rect 20996 12588 21048 12597
rect 21272 12588 21324 12640
rect 21548 12588 21600 12640
rect 23204 12588 23256 12640
rect 23296 12588 23348 12640
rect 24032 12588 24084 12640
rect 24768 12631 24820 12640
rect 24768 12597 24777 12631
rect 24777 12597 24811 12631
rect 24811 12597 24820 12631
rect 24768 12588 24820 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 12164 12384 12216 12436
rect 13176 12384 13228 12436
rect 13728 12384 13780 12436
rect 14280 12384 14332 12436
rect 17040 12427 17092 12436
rect 17040 12393 17049 12427
rect 17049 12393 17083 12427
rect 17083 12393 17092 12427
rect 17040 12384 17092 12393
rect 19248 12384 19300 12436
rect 20812 12384 20864 12436
rect 21272 12384 21324 12436
rect 23756 12427 23808 12436
rect 23756 12393 23765 12427
rect 23765 12393 23799 12427
rect 23799 12393 23808 12427
rect 23756 12384 23808 12393
rect 24216 12384 24268 12436
rect 24952 12384 25004 12436
rect 11428 12316 11480 12368
rect 13912 12316 13964 12368
rect 18144 12359 18196 12368
rect 18144 12325 18153 12359
rect 18153 12325 18187 12359
rect 18187 12325 18196 12359
rect 18144 12316 18196 12325
rect 21732 12316 21784 12368
rect 23480 12316 23532 12368
rect 11704 12248 11756 12300
rect 12072 12248 12124 12300
rect 12808 12180 12860 12232
rect 17132 12248 17184 12300
rect 19524 12248 19576 12300
rect 20536 12248 20588 12300
rect 23572 12291 23624 12300
rect 23572 12257 23581 12291
rect 23581 12257 23615 12291
rect 23615 12257 23624 12291
rect 23572 12248 23624 12257
rect 24676 12248 24728 12300
rect 13636 12180 13688 12232
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 15476 12180 15528 12232
rect 15660 12223 15712 12232
rect 15660 12189 15676 12223
rect 15676 12189 15710 12223
rect 15710 12189 15712 12223
rect 15660 12180 15712 12189
rect 19432 12180 19484 12232
rect 20076 12180 20128 12232
rect 20720 12180 20772 12232
rect 18052 12155 18104 12164
rect 18052 12121 18061 12155
rect 18061 12121 18095 12155
rect 18095 12121 18104 12155
rect 18052 12112 18104 12121
rect 13544 12044 13596 12096
rect 14188 12044 14240 12096
rect 15292 12044 15344 12096
rect 15476 12087 15528 12096
rect 15476 12053 15485 12087
rect 15485 12053 15519 12087
rect 15519 12053 15528 12087
rect 15476 12044 15528 12053
rect 16028 12044 16080 12096
rect 17592 12087 17644 12096
rect 17592 12053 17601 12087
rect 17601 12053 17635 12087
rect 17635 12053 17644 12087
rect 17592 12044 17644 12053
rect 17684 12044 17736 12096
rect 17868 12044 17920 12096
rect 18236 12044 18288 12096
rect 21364 12044 21416 12096
rect 22100 12044 22152 12096
rect 22836 12044 22888 12096
rect 24124 12087 24176 12096
rect 24124 12053 24133 12087
rect 24133 12053 24167 12087
rect 24167 12053 24176 12087
rect 24124 12044 24176 12053
rect 24768 12087 24820 12096
rect 24768 12053 24777 12087
rect 24777 12053 24811 12087
rect 24811 12053 24820 12087
rect 24768 12044 24820 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 11428 11883 11480 11892
rect 11428 11849 11437 11883
rect 11437 11849 11471 11883
rect 11471 11849 11480 11883
rect 11428 11840 11480 11849
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 14280 11840 14332 11892
rect 14648 11840 14700 11892
rect 15292 11840 15344 11892
rect 15660 11883 15712 11892
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 17960 11840 18012 11892
rect 18972 11840 19024 11892
rect 21732 11840 21784 11892
rect 23664 11840 23716 11892
rect 24676 11883 24728 11892
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 12808 11704 12860 11756
rect 13544 11747 13596 11756
rect 13544 11713 13553 11747
rect 13553 11713 13587 11747
rect 13587 11713 13596 11747
rect 13544 11704 13596 11713
rect 16304 11704 16356 11756
rect 16488 11679 16540 11688
rect 16488 11645 16497 11679
rect 16497 11645 16531 11679
rect 16531 11645 16540 11679
rect 16488 11636 16540 11645
rect 14648 11568 14700 11620
rect 15752 11500 15804 11552
rect 16672 11500 16724 11552
rect 16948 11500 17000 11552
rect 19064 11636 19116 11688
rect 18236 11568 18288 11620
rect 20076 11543 20128 11552
rect 20076 11509 20085 11543
rect 20085 11509 20119 11543
rect 20119 11509 20128 11543
rect 20076 11500 20128 11509
rect 20628 11568 20680 11620
rect 20720 11500 20772 11552
rect 21732 11500 21784 11552
rect 22744 11500 22796 11552
rect 24124 11568 24176 11620
rect 23480 11500 23532 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 12072 11339 12124 11348
rect 12072 11305 12081 11339
rect 12081 11305 12115 11339
rect 12115 11305 12124 11339
rect 12072 11296 12124 11305
rect 13636 11339 13688 11348
rect 13636 11305 13645 11339
rect 13645 11305 13679 11339
rect 13679 11305 13688 11339
rect 13636 11296 13688 11305
rect 14648 11339 14700 11348
rect 14648 11305 14657 11339
rect 14657 11305 14691 11339
rect 14691 11305 14700 11339
rect 14648 11296 14700 11305
rect 15752 11339 15804 11348
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 15752 11296 15804 11305
rect 18236 11296 18288 11348
rect 18972 11339 19024 11348
rect 18972 11305 18981 11339
rect 18981 11305 19015 11339
rect 19015 11305 19024 11339
rect 18972 11296 19024 11305
rect 20996 11296 21048 11348
rect 21456 11339 21508 11348
rect 21456 11305 21465 11339
rect 21465 11305 21499 11339
rect 21499 11305 21508 11339
rect 21456 11296 21508 11305
rect 25228 11339 25280 11348
rect 25228 11305 25237 11339
rect 25237 11305 25271 11339
rect 25271 11305 25280 11339
rect 25228 11296 25280 11305
rect 14464 11228 14516 11280
rect 14740 11228 14792 11280
rect 17040 11228 17092 11280
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 15292 11160 15344 11212
rect 16580 11160 16632 11212
rect 21272 11203 21324 11212
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 22836 11160 22888 11212
rect 25596 11160 25648 11212
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12532 11092 12584 11101
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 12808 11024 12860 11076
rect 13728 11024 13780 11076
rect 14556 11092 14608 11144
rect 15384 11092 15436 11144
rect 16948 11135 17000 11144
rect 1492 10956 1544 11008
rect 11888 10999 11940 11008
rect 11888 10965 11897 10999
rect 11897 10965 11931 10999
rect 11931 10965 11940 10999
rect 11888 10956 11940 10965
rect 12624 10956 12676 11008
rect 12900 10956 12952 11008
rect 14740 10956 14792 11008
rect 15660 11024 15712 11076
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 20536 11092 20588 11144
rect 22008 11092 22060 11144
rect 25412 11135 25464 11144
rect 16304 11067 16356 11076
rect 16304 11033 16313 11067
rect 16313 11033 16347 11067
rect 16347 11033 16356 11067
rect 16304 11024 16356 11033
rect 16672 11067 16724 11076
rect 16672 11033 16681 11067
rect 16681 11033 16715 11067
rect 16715 11033 16724 11067
rect 16672 11024 16724 11033
rect 19432 11067 19484 11076
rect 19432 11033 19441 11067
rect 19441 11033 19475 11067
rect 19475 11033 19484 11067
rect 19432 11024 19484 11033
rect 20168 10956 20220 11008
rect 20536 10999 20588 11008
rect 20536 10965 20545 10999
rect 20545 10965 20579 10999
rect 20579 10965 20588 10999
rect 20536 10956 20588 10965
rect 20720 11024 20772 11076
rect 22192 11024 22244 11076
rect 25412 11101 25421 11135
rect 25421 11101 25455 11135
rect 25455 11101 25464 11135
rect 25412 11092 25464 11101
rect 23572 11024 23624 11076
rect 20904 10956 20956 11008
rect 23848 10956 23900 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 11612 10752 11664 10804
rect 12624 10752 12676 10804
rect 13636 10752 13688 10804
rect 13912 10752 13964 10804
rect 14464 10752 14516 10804
rect 16948 10795 17000 10804
rect 16948 10761 16957 10795
rect 16957 10761 16991 10795
rect 16991 10761 17000 10795
rect 16948 10752 17000 10761
rect 17040 10752 17092 10804
rect 18880 10752 18932 10804
rect 22836 10795 22888 10804
rect 22836 10761 22845 10795
rect 22845 10761 22879 10795
rect 22879 10761 22888 10795
rect 22836 10752 22888 10761
rect 25412 10752 25464 10804
rect 10876 10727 10928 10736
rect 10876 10693 10885 10727
rect 10885 10693 10919 10727
rect 10919 10693 10928 10727
rect 10876 10684 10928 10693
rect 8208 10616 8260 10668
rect 9404 10616 9456 10668
rect 1492 10548 1544 10600
rect 1676 10591 1728 10600
rect 1676 10557 1710 10591
rect 1710 10557 1728 10591
rect 1676 10548 1728 10557
rect 16764 10684 16816 10736
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 14648 10659 14700 10668
rect 12624 10548 12676 10600
rect 14648 10625 14657 10659
rect 14657 10625 14691 10659
rect 14691 10625 14700 10659
rect 16212 10659 16264 10668
rect 14648 10616 14700 10625
rect 16212 10625 16221 10659
rect 16221 10625 16255 10659
rect 16255 10625 16264 10659
rect 16212 10616 16264 10625
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 13544 10548 13596 10600
rect 14556 10548 14608 10600
rect 15752 10548 15804 10600
rect 19064 10548 19116 10600
rect 21916 10591 21968 10600
rect 21916 10557 21925 10591
rect 21925 10557 21959 10591
rect 21959 10557 21968 10591
rect 21916 10548 21968 10557
rect 11888 10480 11940 10532
rect 13912 10480 13964 10532
rect 16488 10480 16540 10532
rect 20812 10480 20864 10532
rect 23848 10480 23900 10532
rect 2780 10455 2832 10464
rect 2780 10421 2789 10455
rect 2789 10421 2823 10455
rect 2823 10421 2832 10455
rect 2780 10412 2832 10421
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 15568 10412 15620 10464
rect 20168 10412 20220 10464
rect 21548 10412 21600 10464
rect 22192 10412 22244 10464
rect 23664 10412 23716 10464
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 25596 10455 25648 10464
rect 25596 10421 25605 10455
rect 25605 10421 25639 10455
rect 25639 10421 25648 10455
rect 25596 10412 25648 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 11888 10208 11940 10260
rect 12900 10208 12952 10260
rect 13728 10251 13780 10260
rect 13728 10217 13737 10251
rect 13737 10217 13771 10251
rect 13771 10217 13780 10251
rect 13728 10208 13780 10217
rect 14280 10208 14332 10260
rect 15292 10251 15344 10260
rect 15292 10217 15301 10251
rect 15301 10217 15335 10251
rect 15335 10217 15344 10251
rect 15292 10208 15344 10217
rect 16212 10208 16264 10260
rect 16580 10208 16632 10260
rect 18420 10251 18472 10260
rect 18420 10217 18429 10251
rect 18429 10217 18463 10251
rect 18463 10217 18472 10251
rect 18420 10208 18472 10217
rect 13636 10140 13688 10192
rect 14096 10183 14148 10192
rect 14096 10149 14105 10183
rect 14105 10149 14139 10183
rect 14139 10149 14148 10183
rect 14096 10140 14148 10149
rect 15568 10140 15620 10192
rect 16120 10140 16172 10192
rect 17868 10140 17920 10192
rect 19248 10208 19300 10260
rect 19524 10251 19576 10260
rect 19524 10217 19533 10251
rect 19533 10217 19567 10251
rect 19567 10217 19576 10251
rect 19524 10208 19576 10217
rect 20904 10251 20956 10260
rect 20904 10217 20913 10251
rect 20913 10217 20947 10251
rect 20947 10217 20956 10251
rect 20904 10208 20956 10217
rect 21272 10208 21324 10260
rect 22284 10208 22336 10260
rect 22744 10208 22796 10260
rect 23020 10251 23072 10260
rect 23020 10217 23029 10251
rect 23029 10217 23063 10251
rect 23063 10217 23072 10251
rect 23020 10208 23072 10217
rect 23388 10208 23440 10260
rect 25228 10208 25280 10260
rect 23480 10140 23532 10192
rect 24124 10140 24176 10192
rect 25044 10140 25096 10192
rect 11336 10072 11388 10124
rect 13728 10072 13780 10124
rect 14280 10072 14332 10124
rect 14740 10072 14792 10124
rect 15292 10072 15344 10124
rect 16764 10072 16816 10124
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 11612 10004 11664 10056
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 16212 10004 16264 10056
rect 16948 10004 17000 10056
rect 17776 10072 17828 10124
rect 19064 10072 19116 10124
rect 21548 10072 21600 10124
rect 22100 10072 22152 10124
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 18972 10047 19024 10056
rect 17408 10004 17460 10013
rect 18972 10013 18981 10047
rect 18981 10013 19015 10047
rect 19015 10013 19024 10047
rect 18972 10004 19024 10013
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 21732 10004 21784 10056
rect 12440 9936 12492 9988
rect 15844 9936 15896 9988
rect 12900 9868 12952 9920
rect 13268 9868 13320 9920
rect 14832 9868 14884 9920
rect 15384 9868 15436 9920
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 23664 9868 23716 9920
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 11520 9664 11572 9716
rect 11612 9596 11664 9648
rect 15936 9664 15988 9716
rect 16212 9664 16264 9716
rect 15752 9596 15804 9648
rect 10140 9503 10192 9512
rect 10140 9469 10174 9503
rect 10174 9469 10192 9503
rect 13636 9528 13688 9580
rect 16028 9528 16080 9580
rect 16396 9664 16448 9716
rect 20168 9664 20220 9716
rect 16580 9596 16632 9648
rect 16764 9528 16816 9580
rect 17500 9596 17552 9648
rect 17868 9639 17920 9648
rect 17868 9605 17877 9639
rect 17877 9605 17911 9639
rect 17911 9605 17920 9639
rect 17868 9596 17920 9605
rect 18052 9639 18104 9648
rect 18052 9605 18061 9639
rect 18061 9605 18095 9639
rect 18095 9605 18104 9639
rect 18052 9596 18104 9605
rect 17684 9528 17736 9580
rect 18236 9528 18288 9580
rect 18880 9528 18932 9580
rect 21364 9664 21416 9716
rect 21732 9639 21784 9648
rect 21732 9605 21741 9639
rect 21741 9605 21775 9639
rect 21775 9605 21784 9639
rect 21732 9596 21784 9605
rect 23664 9596 23716 9648
rect 24124 9596 24176 9648
rect 22100 9528 22152 9580
rect 10140 9460 10192 9469
rect 12716 9460 12768 9512
rect 14740 9460 14792 9512
rect 15752 9460 15804 9512
rect 21088 9503 21140 9512
rect 21088 9469 21097 9503
rect 21097 9469 21131 9503
rect 21131 9469 21140 9503
rect 21088 9460 21140 9469
rect 21180 9503 21232 9512
rect 21180 9469 21189 9503
rect 21189 9469 21223 9503
rect 21223 9469 21232 9503
rect 21180 9460 21232 9469
rect 14924 9435 14976 9444
rect 14924 9401 14958 9435
rect 14958 9401 14976 9435
rect 14924 9392 14976 9401
rect 18144 9392 18196 9444
rect 18788 9392 18840 9444
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 11336 9324 11388 9376
rect 12256 9367 12308 9376
rect 12256 9333 12265 9367
rect 12265 9333 12299 9367
rect 12299 9333 12308 9367
rect 12256 9324 12308 9333
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 13728 9324 13780 9376
rect 13912 9367 13964 9376
rect 13912 9333 13921 9367
rect 13921 9333 13955 9367
rect 13955 9333 13964 9367
rect 13912 9324 13964 9333
rect 16764 9324 16816 9376
rect 16948 9367 17000 9376
rect 16948 9333 16957 9367
rect 16957 9333 16991 9367
rect 16991 9333 17000 9367
rect 16948 9324 17000 9333
rect 18880 9324 18932 9376
rect 19064 9367 19116 9376
rect 19064 9333 19073 9367
rect 19073 9333 19107 9367
rect 19107 9333 19116 9367
rect 19064 9324 19116 9333
rect 22008 9324 22060 9376
rect 23480 9392 23532 9444
rect 23388 9367 23440 9376
rect 23388 9333 23397 9367
rect 23397 9333 23431 9367
rect 23431 9333 23440 9367
rect 23388 9324 23440 9333
rect 23572 9324 23624 9376
rect 24768 9460 24820 9512
rect 24860 9324 24912 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 10140 9120 10192 9172
rect 12624 9163 12676 9172
rect 12624 9129 12633 9163
rect 12633 9129 12667 9163
rect 12667 9129 12676 9163
rect 12624 9120 12676 9129
rect 13176 9163 13228 9172
rect 13176 9129 13185 9163
rect 13185 9129 13219 9163
rect 13219 9129 13228 9163
rect 13176 9120 13228 9129
rect 14280 9163 14332 9172
rect 14280 9129 14289 9163
rect 14289 9129 14323 9163
rect 14323 9129 14332 9163
rect 14280 9120 14332 9129
rect 14924 9120 14976 9172
rect 17776 9163 17828 9172
rect 17776 9129 17785 9163
rect 17785 9129 17819 9163
rect 17819 9129 17828 9163
rect 17776 9120 17828 9129
rect 18236 9163 18288 9172
rect 18236 9129 18245 9163
rect 18245 9129 18279 9163
rect 18279 9129 18288 9163
rect 18236 9120 18288 9129
rect 19984 9163 20036 9172
rect 19984 9129 19993 9163
rect 19993 9129 20027 9163
rect 20027 9129 20036 9163
rect 19984 9120 20036 9129
rect 23940 9120 23992 9172
rect 11152 9095 11204 9104
rect 11152 9061 11161 9095
rect 11161 9061 11195 9095
rect 11195 9061 11204 9095
rect 11152 9052 11204 9061
rect 11612 9052 11664 9104
rect 16212 9052 16264 9104
rect 21732 9052 21784 9104
rect 23020 9095 23072 9104
rect 23020 9061 23029 9095
rect 23029 9061 23063 9095
rect 23063 9061 23072 9095
rect 23020 9052 23072 9061
rect 9680 8984 9732 9036
rect 11796 8984 11848 9036
rect 16304 8984 16356 9036
rect 17408 8984 17460 9036
rect 17868 8984 17920 9036
rect 19432 8984 19484 9036
rect 17040 8916 17092 8968
rect 17776 8916 17828 8968
rect 19524 8959 19576 8968
rect 19524 8925 19533 8959
rect 19533 8925 19567 8959
rect 19567 8925 19576 8959
rect 19524 8916 19576 8925
rect 21088 8916 21140 8968
rect 22008 8916 22060 8968
rect 22928 8916 22980 8968
rect 24768 9052 24820 9104
rect 24584 9027 24636 9036
rect 24584 8993 24593 9027
rect 24593 8993 24627 9027
rect 24627 8993 24636 9027
rect 24584 8984 24636 8993
rect 24676 9027 24728 9036
rect 24676 8993 24685 9027
rect 24685 8993 24719 9027
rect 24719 8993 24728 9027
rect 24676 8984 24728 8993
rect 16580 8848 16632 8900
rect 17224 8891 17276 8900
rect 17224 8857 17233 8891
rect 17233 8857 17267 8891
rect 17267 8857 17276 8891
rect 17224 8848 17276 8857
rect 22284 8848 22336 8900
rect 24032 8848 24084 8900
rect 24952 8848 25004 8900
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 18696 8780 18748 8832
rect 22192 8823 22244 8832
rect 22192 8789 22201 8823
rect 22201 8789 22235 8823
rect 22235 8789 22244 8823
rect 22192 8780 22244 8789
rect 22376 8780 22428 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 17868 8576 17920 8628
rect 18328 8576 18380 8628
rect 20996 8576 21048 8628
rect 22008 8576 22060 8628
rect 22928 8619 22980 8628
rect 22928 8585 22937 8619
rect 22937 8585 22971 8619
rect 22971 8585 22980 8619
rect 22928 8576 22980 8585
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 21732 8508 21784 8560
rect 22560 8551 22612 8560
rect 22560 8517 22569 8551
rect 22569 8517 22603 8551
rect 22603 8517 22612 8551
rect 22560 8508 22612 8517
rect 17868 8440 17920 8492
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 14740 8415 14792 8424
rect 14740 8381 14749 8415
rect 14749 8381 14783 8415
rect 14783 8381 14792 8415
rect 14740 8372 14792 8381
rect 18144 8372 18196 8424
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 12624 8304 12676 8356
rect 18420 8347 18472 8356
rect 16304 8279 16356 8288
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 16304 8236 16356 8245
rect 18420 8313 18429 8347
rect 18429 8313 18463 8347
rect 18463 8313 18472 8347
rect 18420 8304 18472 8313
rect 17224 8236 17276 8288
rect 19984 8372 20036 8424
rect 22100 8372 22152 8424
rect 23388 8372 23440 8424
rect 19984 8236 20036 8288
rect 22560 8236 22612 8288
rect 24032 8347 24084 8356
rect 24032 8313 24041 8347
rect 24041 8313 24075 8347
rect 24075 8313 24084 8347
rect 24676 8372 24728 8424
rect 24032 8304 24084 8313
rect 24400 8347 24452 8356
rect 24400 8313 24434 8347
rect 24434 8313 24452 8347
rect 24400 8304 24452 8313
rect 24860 8304 24912 8356
rect 24952 8236 25004 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 12624 8032 12676 8084
rect 13820 8032 13872 8084
rect 14740 8032 14792 8084
rect 16488 8032 16540 8084
rect 16672 8032 16724 8084
rect 17040 8032 17092 8084
rect 17684 8032 17736 8084
rect 17960 8032 18012 8084
rect 19340 8032 19392 8084
rect 21088 8075 21140 8084
rect 21088 8041 21097 8075
rect 21097 8041 21131 8075
rect 21131 8041 21140 8075
rect 21088 8032 21140 8041
rect 24952 8075 25004 8084
rect 24952 8041 24961 8075
rect 24961 8041 24995 8075
rect 24995 8041 25004 8075
rect 24952 8032 25004 8041
rect 16304 7964 16356 8016
rect 21640 7964 21692 8016
rect 22284 7964 22336 8016
rect 24400 7964 24452 8016
rect 12256 7939 12308 7948
rect 12256 7905 12265 7939
rect 12265 7905 12299 7939
rect 12299 7905 12308 7939
rect 12256 7896 12308 7905
rect 13912 7896 13964 7948
rect 17684 7896 17736 7948
rect 18512 7939 18564 7948
rect 18512 7905 18521 7939
rect 18521 7905 18555 7939
rect 18555 7905 18564 7939
rect 18512 7896 18564 7905
rect 21456 7939 21508 7948
rect 21456 7905 21465 7939
rect 21465 7905 21499 7939
rect 21499 7905 21508 7939
rect 21456 7896 21508 7905
rect 22928 7939 22980 7948
rect 22928 7905 22962 7939
rect 22962 7905 22980 7939
rect 22928 7896 22980 7905
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 12716 7828 12768 7880
rect 12808 7828 12860 7880
rect 13452 7828 13504 7880
rect 14188 7828 14240 7880
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 17868 7828 17920 7880
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 12532 7760 12584 7812
rect 17776 7760 17828 7812
rect 19984 7828 20036 7880
rect 21916 7828 21968 7880
rect 19892 7760 19944 7812
rect 22560 7760 22612 7812
rect 11888 7735 11940 7744
rect 11888 7701 11897 7735
rect 11897 7701 11931 7735
rect 11931 7701 11940 7735
rect 11888 7692 11940 7701
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 16488 7735 16540 7744
rect 16488 7701 16497 7735
rect 16497 7701 16531 7735
rect 16531 7701 16540 7735
rect 16488 7692 16540 7701
rect 22100 7692 22152 7744
rect 22652 7692 22704 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 12256 7488 12308 7540
rect 13820 7488 13872 7540
rect 15476 7488 15528 7540
rect 12992 7420 13044 7472
rect 13912 7420 13964 7472
rect 16856 7488 16908 7540
rect 17776 7531 17828 7540
rect 17776 7497 17785 7531
rect 17785 7497 17819 7531
rect 17819 7497 17828 7531
rect 17776 7488 17828 7497
rect 18512 7488 18564 7540
rect 18604 7488 18656 7540
rect 21456 7531 21508 7540
rect 21456 7497 21465 7531
rect 21465 7497 21499 7531
rect 21499 7497 21508 7531
rect 21456 7488 21508 7497
rect 21732 7488 21784 7540
rect 22652 7488 22704 7540
rect 15844 7420 15896 7472
rect 22284 7420 22336 7472
rect 22376 7420 22428 7472
rect 12716 7352 12768 7404
rect 14188 7352 14240 7404
rect 16488 7352 16540 7404
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 15108 7284 15160 7336
rect 17040 7284 17092 7336
rect 18236 7284 18288 7336
rect 18604 7284 18656 7336
rect 21732 7352 21784 7404
rect 22192 7352 22244 7404
rect 22652 7395 22704 7404
rect 22652 7361 22661 7395
rect 22661 7361 22695 7395
rect 22695 7361 22704 7395
rect 22652 7352 22704 7361
rect 24124 7395 24176 7404
rect 19524 7284 19576 7336
rect 22376 7327 22428 7336
rect 22376 7293 22385 7327
rect 22385 7293 22419 7327
rect 22419 7293 22428 7327
rect 22376 7284 22428 7293
rect 22560 7284 22612 7336
rect 12624 7148 12676 7200
rect 17868 7216 17920 7268
rect 19340 7216 19392 7268
rect 19892 7216 19944 7268
rect 21456 7216 21508 7268
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 13820 7148 13872 7200
rect 17684 7148 17736 7200
rect 18420 7148 18472 7200
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 22008 7191 22060 7200
rect 22008 7157 22017 7191
rect 22017 7157 22051 7191
rect 22051 7157 22060 7191
rect 22008 7148 22060 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 12348 6944 12400 6996
rect 13452 6944 13504 6996
rect 16488 6944 16540 6996
rect 17316 6987 17368 6996
rect 17316 6953 17325 6987
rect 17325 6953 17359 6987
rect 17359 6953 17368 6987
rect 17316 6944 17368 6953
rect 21916 6944 21968 6996
rect 22192 6944 22244 6996
rect 22928 6944 22980 6996
rect 24308 6944 24360 6996
rect 13544 6851 13596 6860
rect 13544 6817 13553 6851
rect 13553 6817 13587 6851
rect 13587 6817 13596 6851
rect 13544 6808 13596 6817
rect 16396 6876 16448 6928
rect 17224 6876 17276 6928
rect 17592 6876 17644 6928
rect 18880 6851 18932 6860
rect 18880 6817 18889 6851
rect 18889 6817 18923 6851
rect 18923 6817 18932 6851
rect 18880 6808 18932 6817
rect 20076 6808 20128 6860
rect 13636 6740 13688 6792
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 15568 6672 15620 6724
rect 17960 6672 18012 6724
rect 18788 6740 18840 6792
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19064 6740 19116 6749
rect 21548 6740 21600 6792
rect 21732 6783 21784 6792
rect 21732 6749 21741 6783
rect 21741 6749 21775 6783
rect 21775 6749 21784 6783
rect 22560 6808 22612 6860
rect 23020 6851 23072 6860
rect 23020 6817 23054 6851
rect 23054 6817 23072 6851
rect 23020 6808 23072 6817
rect 25228 6851 25280 6860
rect 25228 6817 25237 6851
rect 25237 6817 25271 6851
rect 25271 6817 25280 6851
rect 25228 6808 25280 6817
rect 21732 6740 21784 6749
rect 22008 6740 22060 6792
rect 21180 6715 21232 6724
rect 21180 6681 21189 6715
rect 21189 6681 21223 6715
rect 21223 6681 21232 6715
rect 21180 6672 21232 6681
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 13728 6604 13780 6656
rect 14188 6647 14240 6656
rect 14188 6613 14197 6647
rect 14197 6613 14231 6647
rect 14231 6613 14240 6647
rect 14188 6604 14240 6613
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 16488 6647 16540 6656
rect 16488 6613 16497 6647
rect 16497 6613 16531 6647
rect 16531 6613 16540 6647
rect 16488 6604 16540 6613
rect 18604 6604 18656 6656
rect 21640 6604 21692 6656
rect 22192 6647 22244 6656
rect 22192 6613 22201 6647
rect 22201 6613 22235 6647
rect 22235 6613 22244 6647
rect 22192 6604 22244 6613
rect 25412 6647 25464 6656
rect 25412 6613 25421 6647
rect 25421 6613 25455 6647
rect 25455 6613 25464 6647
rect 25412 6604 25464 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 14740 6400 14792 6452
rect 17316 6400 17368 6452
rect 17592 6400 17644 6452
rect 18880 6400 18932 6452
rect 21640 6400 21692 6452
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 13728 6196 13780 6248
rect 16488 6196 16540 6248
rect 19524 6239 19576 6248
rect 19524 6205 19533 6239
rect 19533 6205 19567 6239
rect 19567 6205 19576 6239
rect 19524 6196 19576 6205
rect 12532 6128 12584 6180
rect 12440 6060 12492 6112
rect 14188 6128 14240 6180
rect 15568 6128 15620 6180
rect 16672 6128 16724 6180
rect 13084 6103 13136 6112
rect 13084 6069 13093 6103
rect 13093 6069 13127 6103
rect 13127 6069 13136 6103
rect 13084 6060 13136 6069
rect 17868 6060 17920 6112
rect 18788 6060 18840 6112
rect 19524 6060 19576 6112
rect 20812 6196 20864 6248
rect 21916 6400 21968 6452
rect 22560 6400 22612 6452
rect 24032 6443 24084 6452
rect 24032 6409 24041 6443
rect 24041 6409 24075 6443
rect 24075 6409 24084 6443
rect 25228 6443 25280 6452
rect 24032 6400 24084 6409
rect 22192 6264 22244 6316
rect 22928 6264 22980 6316
rect 23664 6264 23716 6316
rect 23940 6264 23992 6316
rect 25228 6409 25237 6443
rect 25237 6409 25271 6443
rect 25271 6409 25280 6443
rect 25228 6400 25280 6409
rect 25044 6264 25096 6316
rect 23388 6128 23440 6180
rect 25136 6128 25188 6180
rect 20904 6103 20956 6112
rect 20904 6069 20913 6103
rect 20913 6069 20947 6103
rect 20947 6069 20956 6103
rect 20904 6060 20956 6069
rect 21548 6103 21600 6112
rect 21548 6069 21557 6103
rect 21557 6069 21591 6103
rect 21591 6069 21600 6103
rect 21548 6060 21600 6069
rect 23572 6060 23624 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 13452 5856 13504 5908
rect 15844 5856 15896 5908
rect 19524 5899 19576 5908
rect 19524 5865 19533 5899
rect 19533 5865 19567 5899
rect 19567 5865 19576 5899
rect 19524 5856 19576 5865
rect 21732 5856 21784 5908
rect 22928 5856 22980 5908
rect 25136 5856 25188 5908
rect 12256 5788 12308 5840
rect 12440 5788 12492 5840
rect 16212 5788 16264 5840
rect 19064 5831 19116 5840
rect 19064 5797 19073 5831
rect 19073 5797 19107 5831
rect 19107 5797 19116 5831
rect 19064 5788 19116 5797
rect 21364 5831 21416 5840
rect 21364 5797 21373 5831
rect 21373 5797 21407 5831
rect 21407 5797 21416 5831
rect 21364 5788 21416 5797
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 13636 5720 13688 5772
rect 15844 5720 15896 5772
rect 20076 5720 20128 5772
rect 21272 5763 21324 5772
rect 21272 5729 21281 5763
rect 21281 5729 21315 5763
rect 21315 5729 21324 5763
rect 21272 5720 21324 5729
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 24860 5720 24912 5772
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 16672 5652 16724 5704
rect 20812 5652 20864 5704
rect 23480 5652 23532 5704
rect 15292 5627 15344 5636
rect 15292 5593 15301 5627
rect 15301 5593 15335 5627
rect 15335 5593 15344 5627
rect 15292 5584 15344 5593
rect 23388 5584 23440 5636
rect 24032 5584 24084 5636
rect 13084 5516 13136 5568
rect 17776 5516 17828 5568
rect 20260 5516 20312 5568
rect 20444 5516 20496 5568
rect 20904 5559 20956 5568
rect 20904 5525 20913 5559
rect 20913 5525 20947 5559
rect 20947 5525 20956 5559
rect 20904 5516 20956 5525
rect 22008 5559 22060 5568
rect 22008 5525 22017 5559
rect 22017 5525 22051 5559
rect 22051 5525 22060 5559
rect 22008 5516 22060 5525
rect 23112 5559 23164 5568
rect 23112 5525 23121 5559
rect 23121 5525 23155 5559
rect 23155 5525 23164 5559
rect 23112 5516 23164 5525
rect 23296 5516 23348 5568
rect 25044 5559 25096 5568
rect 25044 5525 25053 5559
rect 25053 5525 25087 5559
rect 25087 5525 25096 5559
rect 25044 5516 25096 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 14280 5312 14332 5364
rect 15936 5312 15988 5364
rect 16212 5312 16264 5364
rect 20168 5312 20220 5364
rect 20812 5312 20864 5364
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 21824 5312 21876 5364
rect 22468 5312 22520 5364
rect 23112 5312 23164 5364
rect 12256 5244 12308 5296
rect 15108 5244 15160 5296
rect 18880 5244 18932 5296
rect 20720 5244 20772 5296
rect 24860 5312 24912 5364
rect 12348 5176 12400 5228
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 19524 5176 19576 5228
rect 20444 5176 20496 5228
rect 20996 5176 21048 5228
rect 23572 5176 23624 5228
rect 13084 5108 13136 5160
rect 13912 5108 13964 5160
rect 14740 5108 14792 5160
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 11428 5040 11480 5092
rect 12348 4972 12400 5024
rect 13176 5040 13228 5092
rect 14188 5040 14240 5092
rect 19984 5108 20036 5160
rect 22100 5108 22152 5160
rect 23296 5108 23348 5160
rect 16672 5015 16724 5024
rect 16672 4981 16681 5015
rect 16681 4981 16715 5015
rect 16715 4981 16724 5015
rect 16672 4972 16724 4981
rect 17040 5015 17092 5024
rect 17040 4981 17049 5015
rect 17049 4981 17083 5015
rect 17083 4981 17092 5015
rect 17040 4972 17092 4981
rect 18972 5040 19024 5092
rect 20168 5040 20220 5092
rect 18880 4972 18932 5024
rect 19524 5015 19576 5024
rect 19524 4981 19533 5015
rect 19533 4981 19567 5015
rect 19567 4981 19576 5015
rect 19524 4972 19576 4981
rect 22468 4972 22520 5024
rect 23112 4972 23164 5024
rect 24032 5040 24084 5092
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 13176 4768 13228 4820
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 14188 4811 14240 4820
rect 14188 4777 14197 4811
rect 14197 4777 14231 4811
rect 14231 4777 14240 4811
rect 14188 4768 14240 4777
rect 15108 4811 15160 4820
rect 15108 4777 15117 4811
rect 15117 4777 15151 4811
rect 15151 4777 15160 4811
rect 15108 4768 15160 4777
rect 17868 4768 17920 4820
rect 18144 4811 18196 4820
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 18236 4768 18288 4820
rect 18880 4811 18932 4820
rect 18880 4777 18889 4811
rect 18889 4777 18923 4811
rect 18923 4777 18932 4811
rect 19984 4811 20036 4820
rect 18880 4768 18932 4777
rect 17500 4700 17552 4752
rect 17684 4700 17736 4752
rect 19984 4777 19993 4811
rect 19993 4777 20027 4811
rect 20027 4777 20036 4811
rect 19984 4768 20036 4777
rect 21272 4768 21324 4820
rect 23296 4768 23348 4820
rect 23480 4768 23532 4820
rect 12072 4632 12124 4684
rect 12440 4675 12492 4684
rect 12440 4641 12474 4675
rect 12474 4641 12492 4675
rect 12440 4632 12492 4641
rect 15476 4632 15528 4684
rect 20076 4700 20128 4752
rect 23848 4700 23900 4752
rect 24952 4700 25004 4752
rect 19156 4632 19208 4684
rect 20996 4632 21048 4684
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 17776 4564 17828 4616
rect 19064 4607 19116 4616
rect 19064 4573 19073 4607
rect 19073 4573 19107 4607
rect 19107 4573 19116 4607
rect 19064 4564 19116 4573
rect 19616 4564 19668 4616
rect 20812 4564 20864 4616
rect 19248 4496 19300 4548
rect 23204 4632 23256 4684
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 15844 4428 15896 4480
rect 16028 4471 16080 4480
rect 16028 4437 16037 4471
rect 16037 4437 16071 4471
rect 16071 4437 16080 4471
rect 16028 4428 16080 4437
rect 16580 4428 16632 4480
rect 19524 4428 19576 4480
rect 19984 4428 20036 4480
rect 23112 4428 23164 4480
rect 24768 4471 24820 4480
rect 24768 4437 24777 4471
rect 24777 4437 24811 4471
rect 24811 4437 24820 4471
rect 24768 4428 24820 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 12072 4224 12124 4276
rect 6368 4088 6420 4140
rect 6828 4088 6880 4140
rect 7748 4088 7800 4140
rect 8208 4088 8260 4140
rect 12440 4224 12492 4276
rect 12716 4224 12768 4276
rect 15476 4224 15528 4276
rect 17408 4224 17460 4276
rect 20536 4224 20588 4276
rect 20996 4267 21048 4276
rect 20996 4233 21005 4267
rect 21005 4233 21039 4267
rect 21039 4233 21048 4267
rect 20996 4224 21048 4233
rect 25044 4267 25096 4276
rect 25044 4233 25053 4267
rect 25053 4233 25087 4267
rect 25087 4233 25096 4267
rect 25044 4224 25096 4233
rect 12532 4088 12584 4140
rect 13268 4088 13320 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 18144 4156 18196 4208
rect 13912 4020 13964 4072
rect 16580 4063 16632 4072
rect 16580 4029 16589 4063
rect 16589 4029 16623 4063
rect 16623 4029 16632 4063
rect 18236 4088 18288 4140
rect 19064 4156 19116 4208
rect 20812 4156 20864 4208
rect 23112 4156 23164 4208
rect 19524 4088 19576 4140
rect 16580 4020 16632 4029
rect 18328 4020 18380 4072
rect 19156 4063 19208 4072
rect 19156 4029 19165 4063
rect 19165 4029 19199 4063
rect 19199 4029 19208 4063
rect 19156 4020 19208 4029
rect 19616 4063 19668 4072
rect 12348 3952 12400 4004
rect 13544 3952 13596 4004
rect 16212 3952 16264 4004
rect 11152 3884 11204 3936
rect 14832 3884 14884 3936
rect 16304 3884 16356 3936
rect 18236 3884 18288 3936
rect 19616 4029 19625 4063
rect 19625 4029 19659 4063
rect 19659 4029 19668 4063
rect 19616 4020 19668 4029
rect 22192 4063 22244 4072
rect 22192 4029 22201 4063
rect 22201 4029 22235 4063
rect 22235 4029 22244 4063
rect 22192 4020 22244 4029
rect 19984 3952 20036 4004
rect 23848 3952 23900 4004
rect 22376 3927 22428 3936
rect 22376 3893 22385 3927
rect 22385 3893 22419 3927
rect 22419 3893 22428 3927
rect 22376 3884 22428 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 12716 3723 12768 3732
rect 12716 3689 12725 3723
rect 12725 3689 12759 3723
rect 12759 3689 12768 3723
rect 12716 3680 12768 3689
rect 13544 3680 13596 3732
rect 14096 3723 14148 3732
rect 14096 3689 14105 3723
rect 14105 3689 14139 3723
rect 14139 3689 14148 3723
rect 14096 3680 14148 3689
rect 18880 3680 18932 3732
rect 19248 3723 19300 3732
rect 19248 3689 19257 3723
rect 19257 3689 19291 3723
rect 19291 3689 19300 3723
rect 19248 3680 19300 3689
rect 19524 3680 19576 3732
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 22100 3723 22152 3732
rect 22100 3689 22109 3723
rect 22109 3689 22143 3723
rect 22143 3689 22152 3723
rect 22468 3723 22520 3732
rect 22100 3680 22152 3689
rect 22468 3689 22477 3723
rect 22477 3689 22511 3723
rect 22511 3689 22520 3723
rect 22468 3680 22520 3689
rect 23296 3723 23348 3732
rect 23296 3689 23305 3723
rect 23305 3689 23339 3723
rect 23339 3689 23348 3723
rect 23296 3680 23348 3689
rect 24860 3723 24912 3732
rect 24860 3689 24869 3723
rect 24869 3689 24903 3723
rect 24903 3689 24912 3723
rect 24860 3680 24912 3689
rect 24952 3680 25004 3732
rect 13912 3612 13964 3664
rect 14556 3612 14608 3664
rect 10692 3544 10744 3596
rect 11336 3544 11388 3596
rect 12992 3544 13044 3596
rect 14188 3544 14240 3596
rect 14832 3476 14884 3528
rect 15660 3544 15712 3596
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 21456 3612 21508 3664
rect 22744 3655 22796 3664
rect 22744 3621 22753 3655
rect 22753 3621 22787 3655
rect 22787 3621 22796 3655
rect 22744 3612 22796 3621
rect 23204 3655 23256 3664
rect 23204 3621 23213 3655
rect 23213 3621 23247 3655
rect 23247 3621 23256 3655
rect 23204 3612 23256 3621
rect 16488 3544 16540 3596
rect 16672 3587 16724 3596
rect 16672 3553 16706 3587
rect 16706 3553 16724 3587
rect 16672 3544 16724 3553
rect 15384 3476 15436 3528
rect 19156 3476 19208 3528
rect 13636 3451 13688 3460
rect 13636 3417 13645 3451
rect 13645 3417 13679 3451
rect 13679 3417 13688 3451
rect 13636 3408 13688 3417
rect 19064 3408 19116 3460
rect 19616 3476 19668 3528
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 21732 3476 21784 3528
rect 20904 3451 20956 3460
rect 20904 3417 20913 3451
rect 20913 3417 20947 3451
rect 20947 3417 20956 3451
rect 20904 3408 20956 3417
rect 23296 3408 23348 3460
rect 23756 3519 23808 3528
rect 23756 3485 23765 3519
rect 23765 3485 23799 3519
rect 23799 3485 23808 3519
rect 23756 3476 23808 3485
rect 23848 3476 23900 3528
rect 24860 3476 24912 3528
rect 25504 3519 25556 3528
rect 25504 3485 25513 3519
rect 25513 3485 25547 3519
rect 25547 3485 25556 3519
rect 25504 3476 25556 3485
rect 24768 3408 24820 3460
rect 10876 3340 10928 3392
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 14832 3340 14884 3392
rect 15476 3383 15528 3392
rect 15476 3349 15485 3383
rect 15485 3349 15519 3383
rect 15519 3349 15528 3383
rect 15476 3340 15528 3349
rect 17408 3340 17460 3392
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 18880 3340 18932 3349
rect 20352 3383 20404 3392
rect 20352 3349 20361 3383
rect 20361 3349 20395 3383
rect 20395 3349 20404 3383
rect 20352 3340 20404 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 10692 3179 10744 3188
rect 10692 3145 10701 3179
rect 10701 3145 10735 3179
rect 10735 3145 10744 3179
rect 10692 3136 10744 3145
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 12992 3179 13044 3188
rect 12992 3145 13001 3179
rect 13001 3145 13035 3179
rect 13035 3145 13044 3179
rect 12992 3136 13044 3145
rect 13452 3136 13504 3188
rect 14188 3136 14240 3188
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 17500 3136 17552 3188
rect 20352 3136 20404 3188
rect 21732 3179 21784 3188
rect 21732 3145 21741 3179
rect 21741 3145 21775 3179
rect 21775 3145 21784 3179
rect 21732 3136 21784 3145
rect 23296 3179 23348 3188
rect 23296 3145 23305 3179
rect 23305 3145 23339 3179
rect 23339 3145 23348 3179
rect 23296 3136 23348 3145
rect 23756 3136 23808 3188
rect 24860 3136 24912 3188
rect 25504 3136 25556 3188
rect 11060 3068 11112 3120
rect 10784 3000 10836 3052
rect 10140 2932 10192 2984
rect 10692 2932 10744 2984
rect 10968 2932 11020 2984
rect 11428 3111 11480 3120
rect 11428 3077 11437 3111
rect 11437 3077 11471 3111
rect 11471 3077 11480 3111
rect 11428 3068 11480 3077
rect 16672 3068 16724 3120
rect 17132 3068 17184 3120
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 14096 3000 14148 3052
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 16488 3000 16540 3052
rect 18236 3043 18288 3052
rect 18236 3009 18245 3043
rect 18245 3009 18279 3043
rect 18279 3009 18288 3043
rect 18236 3000 18288 3009
rect 21364 3068 21416 3120
rect 19984 3000 20036 3052
rect 13452 2975 13504 2984
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 13452 2932 13504 2941
rect 19432 2932 19484 2984
rect 11336 2864 11388 2916
rect 14832 2907 14884 2916
rect 14832 2873 14866 2907
rect 14866 2873 14884 2907
rect 14832 2864 14884 2873
rect 20812 2932 20864 2984
rect 21088 2975 21140 2984
rect 21088 2941 21097 2975
rect 21097 2941 21131 2975
rect 21131 2941 21140 2975
rect 21088 2932 21140 2941
rect 22560 2932 22612 2984
rect 24952 3000 25004 3052
rect 13636 2839 13688 2848
rect 13636 2805 13645 2839
rect 13645 2805 13679 2839
rect 13679 2805 13688 2839
rect 13636 2796 13688 2805
rect 17408 2839 17460 2848
rect 17408 2805 17417 2839
rect 17417 2805 17451 2839
rect 17451 2805 17460 2839
rect 21456 2864 21508 2916
rect 22652 2839 22704 2848
rect 17408 2796 17460 2805
rect 22652 2805 22661 2839
rect 22661 2805 22695 2839
rect 22695 2805 22704 2839
rect 22652 2796 22704 2805
rect 24768 2839 24820 2848
rect 24768 2805 24777 2839
rect 24777 2805 24811 2839
rect 24811 2805 24820 2839
rect 24768 2796 24820 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2964 2635 3016 2644
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 13084 2635 13136 2644
rect 13084 2601 13093 2635
rect 13093 2601 13127 2635
rect 13127 2601 13136 2635
rect 13084 2592 13136 2601
rect 14740 2592 14792 2644
rect 16120 2592 16172 2644
rect 17132 2635 17184 2644
rect 17132 2601 17141 2635
rect 17141 2601 17175 2635
rect 17175 2601 17184 2635
rect 19064 2635 19116 2644
rect 17132 2592 17184 2601
rect 19064 2601 19073 2635
rect 19073 2601 19107 2635
rect 19107 2601 19116 2635
rect 19064 2592 19116 2601
rect 19524 2635 19576 2644
rect 19524 2601 19533 2635
rect 19533 2601 19567 2635
rect 19567 2601 19576 2635
rect 19524 2592 19576 2601
rect 20352 2592 20404 2644
rect 20812 2635 20864 2644
rect 20812 2601 20821 2635
rect 20821 2601 20855 2635
rect 20855 2601 20864 2635
rect 20812 2592 20864 2601
rect 22468 2592 22520 2644
rect 23848 2635 23900 2644
rect 23848 2601 23857 2635
rect 23857 2601 23891 2635
rect 23891 2601 23900 2635
rect 23848 2592 23900 2601
rect 2964 2456 3016 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 8392 2456 8444 2508
rect 11520 2524 11572 2576
rect 11060 2456 11112 2508
rect 14832 2524 14884 2576
rect 15752 2567 15804 2576
rect 15752 2533 15761 2567
rect 15761 2533 15795 2567
rect 15795 2533 15804 2567
rect 15752 2524 15804 2533
rect 16304 2524 16356 2576
rect 18052 2567 18104 2576
rect 18052 2533 18061 2567
rect 18061 2533 18095 2567
rect 18095 2533 18104 2567
rect 18052 2524 18104 2533
rect 14648 2456 14700 2508
rect 18420 2499 18472 2508
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18420 2456 18472 2465
rect 14464 2363 14516 2372
rect 14464 2329 14473 2363
rect 14473 2329 14507 2363
rect 14507 2329 14516 2363
rect 14464 2320 14516 2329
rect 17408 2388 17460 2440
rect 18972 2388 19024 2440
rect 20536 2456 20588 2508
rect 21640 2456 21692 2508
rect 22836 2499 22888 2508
rect 22836 2465 22845 2499
rect 22845 2465 22879 2499
rect 22879 2465 22888 2499
rect 22836 2456 22888 2465
rect 23940 2456 23992 2508
rect 19892 2320 19944 2372
rect 24676 2320 24728 2372
rect 26148 2320 26200 2372
rect 8392 2252 8444 2304
rect 10968 2252 11020 2304
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 21916 2295 21968 2304
rect 21916 2261 21925 2295
rect 21925 2261 21959 2295
rect 21959 2261 21968 2295
rect 21916 2252 21968 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 12808 552 12860 604
rect 13176 552 13228 604
rect 20444 552 20496 604
rect 21364 552 21416 604
<< metal2 >>
rect 294 27520 350 28000
rect 938 27520 994 28000
rect 1582 27520 1638 28000
rect 2318 27520 2374 28000
rect 2962 27520 3018 28000
rect 3698 27520 3754 28000
rect 4342 27520 4398 28000
rect 4986 27520 5042 28000
rect 5722 27520 5778 28000
rect 6366 27520 6422 28000
rect 7102 27520 7158 28000
rect 7746 27520 7802 28000
rect 8390 27520 8446 28000
rect 9126 27520 9182 28000
rect 9770 27520 9826 28000
rect 10506 27520 10562 28000
rect 11150 27520 11206 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13174 27520 13230 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15290 27520 15346 28000
rect 15934 27520 15990 28000
rect 16578 27520 16634 28000
rect 17314 27520 17370 28000
rect 17958 27520 18014 28000
rect 18694 27520 18750 28000
rect 19338 27520 19394 28000
rect 20074 27520 20130 28000
rect 20718 27520 20774 28000
rect 21362 27520 21418 28000
rect 22098 27520 22154 28000
rect 22742 27520 22798 28000
rect 23202 27704 23258 27713
rect 23202 27639 23258 27648
rect 308 27418 336 27520
rect 32 27390 336 27418
rect 32 17746 60 27390
rect 952 22658 980 27520
rect 1596 24721 1624 27520
rect 1582 24712 1638 24721
rect 1582 24647 1638 24656
rect 1490 22672 1546 22681
rect 952 22630 1490 22658
rect 1490 22607 1546 22616
rect 1952 21004 2004 21010
rect 1952 20946 2004 20952
rect 1582 20904 1638 20913
rect 1582 20839 1584 20848
rect 1636 20839 1638 20848
rect 1584 20810 1636 20816
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1582 20360 1638 20369
rect 1412 19718 1440 20334
rect 1582 20295 1638 20304
rect 1596 20262 1624 20295
rect 1964 20262 1992 20946
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 1400 19712 1452 19718
rect 1400 19654 1452 19660
rect 20 17740 72 17746
rect 20 17682 72 17688
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 294 1728 350 1737
rect 294 1663 350 1672
rect 308 480 336 1663
rect 952 480 980 3431
rect 1412 3346 1440 19654
rect 1674 13968 1730 13977
rect 1674 13903 1730 13912
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10606 1532 10950
rect 1688 10606 1716 13903
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1504 9761 1532 10542
rect 1688 10266 1716 10542
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1490 9752 1546 9761
rect 1490 9687 1546 9696
rect 1964 3505 1992 20198
rect 2332 13297 2360 27520
rect 2976 24857 3004 27520
rect 2962 24848 3018 24857
rect 2962 24783 3018 24792
rect 3712 22545 3740 27520
rect 4356 23769 4384 27520
rect 5000 24177 5028 27520
rect 5736 25242 5764 27520
rect 5736 25214 6040 25242
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 4986 24168 5042 24177
rect 4986 24103 5042 24112
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 4342 23760 4398 23769
rect 4342 23695 4398 23704
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 3698 22536 3754 22545
rect 3698 22471 3754 22480
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21729 6040 25214
rect 6380 23905 6408 27520
rect 6366 23896 6422 23905
rect 6366 23831 6422 23840
rect 5998 21720 6054 21729
rect 5998 21655 6054 21664
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 7116 19281 7144 27520
rect 7102 19272 7158 19281
rect 7102 19207 7158 19216
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 7760 17785 7788 27520
rect 8404 24818 8432 27520
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 9140 20777 9168 27520
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9126 20768 9182 20777
rect 9126 20703 9182 20712
rect 9600 19258 9628 24754
rect 9784 21049 9812 27520
rect 10520 25786 10548 27520
rect 10520 25758 10732 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10704 23225 10732 25758
rect 10690 23216 10746 23225
rect 10690 23151 10746 23160
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10796 22778 10824 23054
rect 11072 22778 11100 23122
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 9954 22264 10010 22273
rect 10289 22256 10585 22276
rect 9954 22199 10010 22208
rect 9770 21040 9826 21049
rect 9770 20975 9826 20984
rect 9968 19825 9996 22199
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11072 21729 11100 21966
rect 11058 21720 11114 21729
rect 11058 21655 11060 21664
rect 11112 21655 11114 21664
rect 11060 21626 11112 21632
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10048 20528 10100 20534
rect 10048 20470 10100 20476
rect 10322 20496 10378 20505
rect 10060 19922 10088 20470
rect 11164 20482 11192 27520
rect 11900 24449 11928 27520
rect 12346 24848 12402 24857
rect 12346 24783 12402 24792
rect 11886 24440 11942 24449
rect 12360 24410 12388 24783
rect 11886 24375 11942 24384
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11532 24177 11560 24210
rect 11518 24168 11574 24177
rect 12360 24154 12388 24346
rect 11518 24103 11574 24112
rect 12268 24126 12388 24154
rect 11426 23896 11482 23905
rect 11532 23866 11560 24103
rect 12268 23866 12296 24126
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 11426 23831 11482 23840
rect 11520 23860 11572 23866
rect 11440 22234 11468 23831
rect 11520 23802 11572 23808
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 11532 23746 11560 23802
rect 11532 23718 11652 23746
rect 11520 22704 11572 22710
rect 11520 22646 11572 22652
rect 11428 22228 11480 22234
rect 11428 22170 11480 22176
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11256 20602 11284 20946
rect 11348 20942 11376 21490
rect 11440 21332 11468 22170
rect 11532 21554 11560 22646
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11520 21344 11572 21350
rect 11440 21304 11520 21332
rect 11520 21286 11572 21292
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11348 20602 11376 20878
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11164 20454 11284 20482
rect 10322 20431 10324 20440
rect 10376 20431 10378 20440
rect 10324 20402 10376 20408
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 9954 19816 10010 19825
rect 9954 19751 10010 19760
rect 10060 19514 10088 19858
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9680 19304 9732 19310
rect 9600 19252 9680 19258
rect 9600 19246 9732 19252
rect 9600 19230 9720 19246
rect 10060 18766 10088 19450
rect 10152 19378 10180 19858
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10782 19272 10838 19281
rect 10782 19207 10838 19216
rect 10796 19174 10824 19207
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10152 18290 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10336 18426 10364 18770
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10612 18426 10640 18702
rect 10796 18630 10824 19110
rect 10888 18834 10916 19314
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10600 18420 10652 18426
rect 10652 18380 10732 18408
rect 10600 18362 10652 18368
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 7746 17776 7802 17785
rect 10704 17746 10732 18380
rect 7746 17711 7802 17720
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 9600 16153 9628 17682
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 9586 16144 9642 16153
rect 9586 16079 9642 16088
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 9494 15192 9550 15201
rect 9416 15150 9494 15178
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 2318 13288 2374 13297
rect 2318 13223 2374 13232
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 4986 11656 5042 11665
rect 4986 11591 5042 11600
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 9625 2820 10406
rect 4342 10160 4398 10169
rect 4342 10095 4398 10104
rect 2870 9752 2926 9761
rect 2870 9687 2926 9696
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 2884 9353 2912 9687
rect 2870 9344 2926 9353
rect 2870 9279 2926 9288
rect 2318 6352 2374 6361
rect 2318 6287 2374 6296
rect 1950 3496 2006 3505
rect 1950 3431 2006 3440
rect 1412 3318 1624 3346
rect 1596 480 1624 3318
rect 2332 480 2360 6287
rect 2884 4729 2912 9279
rect 3698 7984 3754 7993
rect 3698 7919 3754 7928
rect 2962 5128 3018 5137
rect 2962 5063 3018 5072
rect 2870 4720 2926 4729
rect 2870 4655 2926 4664
rect 2976 2650 3004 5063
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2976 480 3004 2450
rect 3712 480 3740 7919
rect 4356 480 4384 10095
rect 5000 480 5028 11591
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 9416 10674 9444 15150
rect 9494 15127 9550 15136
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10796 14657 10824 18566
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10876 17536 10928 17542
rect 11072 17524 11100 18022
rect 10928 17496 11100 17524
rect 10876 17478 10928 17484
rect 10888 17241 10916 17478
rect 10874 17232 10930 17241
rect 10874 17167 10930 17176
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10782 14648 10838 14657
rect 10782 14583 10838 14592
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10876 10736 10928 10742
rect 10874 10704 10876 10713
rect 10928 10704 10930 10713
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 9404 10668 9456 10674
rect 10874 10639 10930 10648
rect 9404 10610 9456 10616
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6918 7576 6974 7585
rect 6918 7511 6974 7520
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6828 4140 6880 4146
rect 6932 4128 6960 7511
rect 8220 4146 8248 10610
rect 10980 10452 11008 17070
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16726 11100 16934
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11072 16250 11100 16662
rect 11164 16590 11192 18294
rect 11256 17921 11284 20454
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11440 19378 11468 19654
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11242 17912 11298 17921
rect 11242 17847 11298 17856
rect 11440 17814 11468 18226
rect 11428 17808 11480 17814
rect 11428 17750 11480 17756
rect 11440 17202 11468 17750
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11256 16794 11284 17138
rect 11336 17060 11388 17066
rect 11336 17002 11388 17008
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11348 16658 11376 17002
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11348 16114 11376 16594
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 10980 10424 11100 10452
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10138 9616 10194 9625
rect 10138 9551 10194 9560
rect 10966 9616 11022 9625
rect 10966 9551 11022 9560
rect 10152 9518 10180 9551
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 9680 9376 9732 9382
rect 9678 9344 9680 9353
rect 9732 9344 9734 9353
rect 9678 9279 9734 9288
rect 9692 9042 9720 9279
rect 10152 9178 10180 9454
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9126 8936 9182 8945
rect 9126 8871 9182 8880
rect 8298 4720 8354 4729
rect 8298 4655 8354 4664
rect 6880 4100 6960 4128
rect 7748 4140 7800 4146
rect 6828 4082 6880 4088
rect 7748 4082 7800 4088
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5736 2553 5764 2586
rect 5722 2544 5778 2553
rect 5540 2508 5592 2514
rect 5722 2479 5778 2488
rect 5540 2450 5592 2456
rect 5552 1578 5580 2450
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5552 1550 5764 1578
rect 5736 480 5764 1550
rect 6380 480 6408 4082
rect 7102 4040 7158 4049
rect 7102 3975 7158 3984
rect 7116 480 7144 3975
rect 7760 480 7788 4082
rect 8312 2650 8340 4655
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8404 2310 8432 2450
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8404 480 8432 2246
rect 9140 480 9168 8871
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10782 4992 10838 5001
rect 10289 4924 10585 4944
rect 10782 4927 10838 4936
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 9770 4584 9826 4593
rect 9770 4519 9826 4528
rect 9784 480 9812 4519
rect 10690 4176 10746 4185
rect 10690 4111 10746 4120
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3602 10732 4111
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10138 3224 10194 3233
rect 10704 3194 10732 3538
rect 10138 3159 10140 3168
rect 10192 3159 10194 3168
rect 10692 3188 10744 3194
rect 10140 3130 10192 3136
rect 10692 3130 10744 3136
rect 10152 2990 10180 3130
rect 10796 3058 10824 4927
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 1442 10732 2926
rect 10888 2650 10916 3334
rect 10980 2990 11008 9551
rect 11072 8537 11100 10424
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11164 8634 11192 9046
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11058 8528 11114 8537
rect 11058 8463 11114 8472
rect 11072 4049 11100 8463
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11164 3194 11192 3878
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11072 2514 11100 3062
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 1465 11008 2246
rect 10520 1414 10732 1442
rect 10966 1456 11022 1465
rect 10520 480 10548 1414
rect 10966 1391 11022 1400
rect 11256 626 11284 13738
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11440 11898 11468 12310
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11532 10146 11560 21286
rect 11624 14521 11652 23718
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11808 22030 11836 22918
rect 12360 22114 12388 24006
rect 12440 23656 12492 23662
rect 12544 23633 12572 27520
rect 12990 24712 13046 24721
rect 12990 24647 13046 24656
rect 13004 24614 13032 24647
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12728 23662 12756 24142
rect 13188 23769 13216 27520
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13174 23760 13230 23769
rect 13174 23695 13230 23704
rect 12716 23656 12768 23662
rect 12440 23598 12492 23604
rect 12530 23624 12586 23633
rect 12452 23050 12480 23598
rect 12716 23598 12768 23604
rect 12530 23559 12586 23568
rect 12530 23216 12586 23225
rect 12530 23151 12586 23160
rect 12900 23180 12952 23186
rect 12440 23044 12492 23050
rect 12440 22986 12492 22992
rect 12452 22642 12480 22986
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12360 22086 12480 22114
rect 12452 22030 12480 22086
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 11808 21350 11836 21966
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 12176 21350 12204 21558
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 11702 21040 11758 21049
rect 11808 21010 11836 21286
rect 11702 20975 11758 20984
rect 11796 21004 11848 21010
rect 11716 18193 11744 20975
rect 11796 20946 11848 20952
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11808 19718 11836 20198
rect 12176 20058 12204 21286
rect 12360 20346 12388 21830
rect 12544 21570 12572 23151
rect 12900 23122 12952 23128
rect 12716 22500 12768 22506
rect 12716 22442 12768 22448
rect 12728 22098 12756 22442
rect 12912 22234 12940 23122
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 12544 21542 13032 21570
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12544 20602 12572 21354
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12360 20330 12572 20346
rect 12360 20324 12584 20330
rect 12360 20318 12532 20324
rect 12532 20266 12584 20272
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12070 19952 12126 19961
rect 12176 19922 12204 19994
rect 12070 19887 12126 19896
rect 12164 19916 12216 19922
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11808 19514 11836 19654
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 18290 12020 18566
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11702 18184 11758 18193
rect 11702 18119 11758 18128
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11808 17338 11836 17682
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11808 16182 11836 16526
rect 11992 16250 12020 16526
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11610 14512 11666 14521
rect 11610 14447 11666 14456
rect 11610 14376 11666 14385
rect 11610 14311 11666 14320
rect 11624 10810 11652 14311
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11440 10118 11560 10146
rect 11348 9382 11376 10066
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 8498 11376 9318
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11440 5098 11468 10118
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11532 9722 11560 9998
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11624 9654 11652 9998
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11624 9110 11652 9590
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11348 2922 11376 3538
rect 11440 3210 11468 5034
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11440 3182 11560 3210
rect 11428 3120 11480 3126
rect 11426 3088 11428 3097
rect 11480 3088 11482 3097
rect 11426 3023 11482 3032
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11532 2582 11560 3182
rect 11624 2825 11652 3334
rect 11610 2816 11666 2825
rect 11610 2751 11666 2760
rect 11520 2576 11572 2582
rect 11716 2553 11744 12242
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10538 11928 10950
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11900 10266 11928 10474
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11808 8634 11836 8978
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 5681 11928 7686
rect 11886 5672 11942 5681
rect 11886 5607 11942 5616
rect 11992 5522 12020 12854
rect 12084 12306 12112 19887
rect 12164 19858 12216 19864
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12440 19372 12492 19378
rect 12544 19360 12572 19654
rect 12492 19332 12572 19360
rect 12440 19314 12492 19320
rect 12438 19272 12494 19281
rect 12438 19207 12494 19216
rect 12452 19174 12480 19207
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17134 12572 17478
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12544 16794 12572 17070
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16046 12480 16390
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12636 14958 12664 21286
rect 12820 20874 12848 21286
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12714 20224 12770 20233
rect 12714 20159 12770 20168
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12346 12608 12402 12617
rect 12346 12543 12402 12552
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12176 11898 12204 12378
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12070 11792 12126 11801
rect 12070 11727 12126 11736
rect 12084 11354 12112 11727
rect 12360 11665 12388 12543
rect 12346 11656 12402 11665
rect 12346 11591 12402 11600
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12452 10713 12480 11154
rect 12532 11144 12584 11150
rect 12530 11112 12532 11121
rect 12584 11112 12586 11121
rect 12530 11047 12586 11056
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12636 10810 12664 10950
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12438 10704 12494 10713
rect 12438 10639 12494 10648
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 8945 12296 9318
rect 12254 8936 12310 8945
rect 12254 8871 12310 8880
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12268 7721 12296 7890
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12254 7712 12310 7721
rect 12254 7647 12310 7656
rect 12268 7546 12296 7647
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12360 7002 12388 7822
rect 12452 7585 12480 9930
rect 12636 9178 12664 10542
rect 12728 9518 12756 20159
rect 12820 19281 12848 20810
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12912 20466 12940 20742
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12912 19990 12940 20402
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12912 19378 12940 19926
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12806 19272 12862 19281
rect 12806 19207 12862 19216
rect 12912 18970 12940 19314
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12820 11762 12848 12174
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12820 11082 12848 11698
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10674 12940 10950
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12912 10266 12940 10610
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12912 9382 12940 9862
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12636 8362 12664 9114
rect 12714 9072 12770 9081
rect 12714 9007 12770 9016
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12636 8090 12664 8298
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12530 7984 12586 7993
rect 12530 7919 12586 7928
rect 12544 7818 12572 7919
rect 12728 7886 12756 9007
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12438 7576 12494 7585
rect 12438 7511 12494 7520
rect 12728 7410 12756 7822
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12254 6624 12310 6633
rect 12254 6559 12310 6568
rect 12268 5846 12296 6559
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12440 6112 12492 6118
rect 12360 6060 12440 6066
rect 12360 6054 12492 6060
rect 12360 6038 12480 6054
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11900 5494 12020 5522
rect 11520 2518 11572 2524
rect 11702 2544 11758 2553
rect 11702 2479 11758 2488
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1601 11652 2246
rect 11610 1592 11666 1601
rect 11610 1527 11666 1536
rect 11164 598 11284 626
rect 11164 480 11192 598
rect 11900 480 11928 5494
rect 12084 5370 12112 5646
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 12084 4690 12112 5306
rect 12268 5302 12296 5782
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12360 5234 12388 6038
rect 12544 5930 12572 6122
rect 12452 5902 12572 5930
rect 12452 5846 12480 5902
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12084 4282 12112 4626
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12360 4010 12388 4966
rect 12452 4690 12480 5782
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12452 4282 12480 4626
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12636 4264 12664 7142
rect 12716 4276 12768 4282
rect 12636 4236 12716 4264
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12438 3632 12494 3641
rect 12438 3567 12494 3576
rect 12452 3058 12480 3567
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12544 480 12572 4082
rect 12636 1737 12664 4236
rect 12716 4218 12768 4224
rect 12714 3768 12770 3777
rect 12714 3703 12716 3712
rect 12768 3703 12770 3712
rect 12716 3674 12768 3680
rect 12622 1728 12678 1737
rect 12622 1663 12678 1672
rect 12820 610 12848 7822
rect 12912 6361 12940 9318
rect 13004 7478 13032 21542
rect 13096 14482 13124 22918
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13188 20097 13216 20198
rect 13174 20088 13230 20097
rect 13174 20023 13230 20032
rect 13176 19168 13228 19174
rect 13174 19136 13176 19145
rect 13228 19136 13230 19145
rect 13174 19071 13230 19080
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14482 13216 14758
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13096 14074 13124 14418
rect 13280 14385 13308 24550
rect 13542 24440 13598 24449
rect 13542 24375 13598 24384
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13464 23322 13492 24006
rect 13452 23316 13504 23322
rect 13452 23258 13504 23264
rect 13452 23180 13504 23186
rect 13452 23122 13504 23128
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13372 21146 13400 21966
rect 13464 21894 13492 23122
rect 13556 22012 13584 24375
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13832 23866 13860 24210
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13832 23338 13860 23462
rect 13740 23310 13860 23338
rect 13740 22030 13768 23310
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13832 22778 13860 23054
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13728 22024 13780 22030
rect 13556 21984 13676 22012
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13648 21049 13676 21984
rect 13728 21966 13780 21972
rect 13740 21690 13768 21966
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13820 21344 13872 21350
rect 13740 21292 13820 21298
rect 13740 21286 13872 21292
rect 13740 21270 13860 21286
rect 13634 21040 13690 21049
rect 13634 20975 13690 20984
rect 13360 20528 13412 20534
rect 13360 20470 13412 20476
rect 13372 19922 13400 20470
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13740 18970 13768 21270
rect 13924 18970 13952 27520
rect 14372 25356 14424 25362
rect 14372 25298 14424 25304
rect 14384 24614 14412 25298
rect 14568 24970 14596 27520
rect 15304 25498 15332 27520
rect 15292 25492 15344 25498
rect 15292 25434 15344 25440
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14476 24942 14596 24970
rect 14476 24721 14504 24942
rect 14554 24848 14610 24857
rect 14554 24783 14610 24792
rect 15384 24812 15436 24818
rect 14462 24712 14518 24721
rect 14462 24647 14518 24656
rect 14568 24614 14596 24783
rect 15384 24754 15436 24760
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 14016 23526 14044 24142
rect 14280 23588 14332 23594
rect 14280 23530 14332 23536
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 14094 22128 14150 22137
rect 14094 22063 14150 22072
rect 14108 20913 14136 22063
rect 14094 20904 14150 20913
rect 14094 20839 14150 20848
rect 14094 20768 14150 20777
rect 14094 20703 14150 20712
rect 14108 18970 14136 20703
rect 14188 20256 14240 20262
rect 14186 20224 14188 20233
rect 14240 20224 14242 20233
rect 14186 20159 14242 20168
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14200 19378 14228 19858
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 13924 18426 13952 18906
rect 14108 18737 14136 18906
rect 14200 18766 14228 19110
rect 14188 18760 14240 18766
rect 14094 18728 14150 18737
rect 14188 18702 14240 18708
rect 14094 18663 14150 18672
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13358 18320 13414 18329
rect 13358 18255 13414 18264
rect 13372 18222 13400 18255
rect 14016 18222 14044 18566
rect 14108 18358 14136 18663
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 14200 18290 14228 18702
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 13372 17882 13400 18158
rect 13544 18080 13596 18086
rect 14292 18034 14320 23530
rect 13544 18022 13596 18028
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13358 16552 13414 16561
rect 13358 16487 13414 16496
rect 13266 14376 13322 14385
rect 13266 14311 13322 14320
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13280 13977 13308 14214
rect 13266 13968 13322 13977
rect 13266 13903 13322 13912
rect 13372 13818 13400 16487
rect 13556 16017 13584 18022
rect 13924 18006 14320 18034
rect 13542 16008 13598 16017
rect 13542 15943 13598 15952
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 15065 13768 15846
rect 13726 15056 13782 15065
rect 13726 14991 13782 15000
rect 13450 14784 13506 14793
rect 13450 14719 13506 14728
rect 13280 13790 13400 13818
rect 13082 13288 13138 13297
rect 13082 13223 13138 13232
rect 13096 12889 13124 13223
rect 13082 12880 13138 12889
rect 13082 12815 13138 12824
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12898 6352 12954 6361
rect 13096 6304 13124 12815
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13188 12442 13216 12582
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13188 9178 13216 9998
rect 13280 9926 13308 13790
rect 13358 12744 13414 12753
rect 13358 12679 13414 12688
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13372 7936 13400 12679
rect 13280 7908 13400 7936
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12898 6287 12954 6296
rect 13004 6276 13124 6304
rect 13004 3602 13032 6276
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13096 5574 13124 6054
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 5166 13124 5510
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13188 5098 13216 6598
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13188 4826 13216 5034
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13280 4146 13308 7908
rect 13464 7886 13492 14719
rect 13820 13864 13872 13870
rect 13740 13812 13820 13818
rect 13740 13806 13872 13812
rect 13740 13790 13860 13806
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13556 12322 13584 13398
rect 13740 12442 13768 13790
rect 13924 13530 13952 18006
rect 14002 17912 14058 17921
rect 14002 17847 14058 17856
rect 14016 17814 14044 17847
rect 14004 17808 14056 17814
rect 14280 17808 14332 17814
rect 14004 17750 14056 17756
rect 14278 17776 14280 17785
rect 14332 17776 14334 17785
rect 14016 16794 14044 17750
rect 14278 17711 14334 17720
rect 14292 16998 14320 17711
rect 14280 16992 14332 16998
rect 14278 16960 14280 16969
rect 14332 16960 14334 16969
rect 14278 16895 14334 16904
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14280 16516 14332 16522
rect 14280 16458 14332 16464
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14200 15201 14228 15846
rect 14292 15570 14320 16458
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14186 15192 14242 15201
rect 14292 15162 14320 15506
rect 14186 15127 14242 15136
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14094 14512 14150 14521
rect 14094 14447 14150 14456
rect 14002 13832 14058 13841
rect 14002 13767 14058 13776
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13924 12918 13952 13330
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13924 12617 13952 12650
rect 13910 12608 13966 12617
rect 13910 12543 13966 12552
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13912 12368 13964 12374
rect 13556 12294 13860 12322
rect 13912 12310 13964 12316
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11762 13584 12038
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13648 11354 13676 12174
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13544 10600 13596 10606
rect 13648 10577 13676 10746
rect 13544 10542 13596 10548
rect 13634 10568 13690 10577
rect 13556 10169 13584 10542
rect 13634 10503 13690 10512
rect 13740 10266 13768 11018
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13636 10192 13688 10198
rect 13542 10160 13598 10169
rect 13636 10134 13688 10140
rect 13542 10095 13598 10104
rect 13648 10033 13676 10134
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13634 10024 13690 10033
rect 13634 9959 13690 9968
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13648 8945 13676 9522
rect 13740 9382 13768 10066
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13634 8936 13690 8945
rect 13634 8871 13690 8880
rect 13832 8090 13860 12294
rect 13924 10810 13952 12310
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13924 9625 13952 10474
rect 13910 9616 13966 9625
rect 13910 9551 13966 9560
rect 13912 9376 13964 9382
rect 13910 9344 13912 9353
rect 13964 9344 13966 9353
rect 13910 9279 13966 9288
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7002 13492 7686
rect 13832 7546 13860 8026
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13924 7478 13952 7890
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13464 5914 13492 6938
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13556 6769 13584 6802
rect 13636 6792 13688 6798
rect 13542 6760 13598 6769
rect 13636 6734 13688 6740
rect 13542 6695 13598 6704
rect 13648 6322 13676 6734
rect 13728 6656 13780 6662
rect 13832 6644 13860 7142
rect 13780 6616 13860 6644
rect 13728 6598 13780 6604
rect 13832 6338 13860 6616
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13740 6310 13860 6338
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13450 5808 13506 5817
rect 13648 5778 13676 6258
rect 13740 6254 13768 6310
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13450 5743 13506 5752
rect 13636 5772 13688 5778
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13004 3194 13032 3538
rect 13464 3194 13492 5743
rect 13636 5714 13688 5720
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13556 4826 13584 5170
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13556 4010 13584 4762
rect 13924 4078 13952 5102
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13556 3738 13584 3946
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13924 3670 13952 4014
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 14016 3516 14044 13767
rect 14108 11234 14136 14447
rect 14278 14376 14334 14385
rect 14278 14311 14280 14320
rect 14332 14311 14334 14320
rect 14280 14282 14332 14288
rect 14186 13424 14242 13433
rect 14186 13359 14188 13368
rect 14240 13359 14242 13368
rect 14188 13330 14240 13336
rect 14280 13320 14332 13326
rect 14278 13288 14280 13297
rect 14332 13288 14334 13297
rect 14200 13246 14278 13274
rect 14200 12986 14228 13246
rect 14278 13223 14334 13232
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14200 12102 14228 12718
rect 14292 12442 14320 13126
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14292 11898 14320 12174
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14384 11778 14412 24550
rect 14464 24268 14516 24274
rect 14464 24210 14516 24216
rect 14476 23118 14504 24210
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14568 23905 14596 24074
rect 14554 23896 14610 23905
rect 14554 23831 14610 23840
rect 14464 23112 14516 23118
rect 14462 23080 14464 23089
rect 14516 23080 14518 23089
rect 14462 23015 14518 23024
rect 14568 22930 14596 23831
rect 14476 22902 14596 22930
rect 14476 13462 14504 22902
rect 14660 22794 14688 24686
rect 15028 24138 15056 24686
rect 15396 24585 15424 24754
rect 15580 24682 15608 25298
rect 15948 24857 15976 27520
rect 16592 25498 16620 27520
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 15934 24848 15990 24857
rect 16408 24818 16436 25094
rect 15934 24783 15990 24792
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 15568 24676 15620 24682
rect 15568 24618 15620 24624
rect 15476 24608 15528 24614
rect 15382 24576 15438 24585
rect 15476 24550 15528 24556
rect 15382 24511 15438 24520
rect 15396 24274 15424 24511
rect 15488 24410 15516 24550
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15384 24268 15436 24274
rect 15384 24210 15436 24216
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 15304 22982 15332 23462
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 15474 22944 15530 22953
rect 14568 22766 14688 22794
rect 14568 14006 14596 22766
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14660 19922 14688 20334
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 14660 18714 14688 19858
rect 14752 18902 14780 21286
rect 14844 21146 14872 22918
rect 14956 22876 15252 22896
rect 15474 22879 15530 22888
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14924 22432 14976 22438
rect 14924 22374 14976 22380
rect 15292 22432 15344 22438
rect 15384 22432 15436 22438
rect 15292 22374 15344 22380
rect 15382 22400 15384 22409
rect 15436 22400 15438 22409
rect 14936 22234 14964 22374
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 15304 22030 15332 22374
rect 15382 22335 15438 22344
rect 15488 22250 15516 22879
rect 15396 22222 15516 22250
rect 15292 22024 15344 22030
rect 15290 21992 15292 22001
rect 15344 21992 15346 22001
rect 15290 21927 15346 21936
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15200 21480 15252 21486
rect 15304 21468 15332 21927
rect 15252 21440 15332 21468
rect 15200 21422 15252 21428
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 15396 21078 15424 22222
rect 15384 21072 15436 21078
rect 15384 21014 15436 21020
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 14844 20330 14872 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14844 19174 14872 20266
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 15304 18970 15332 20742
rect 15396 20262 15424 21014
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14660 18686 14780 18714
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14660 18222 14688 18566
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14660 17746 14688 18158
rect 14752 18154 14780 18686
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15396 18329 15424 18566
rect 15382 18320 15438 18329
rect 15382 18255 15438 18264
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14752 17814 14780 18090
rect 14740 17808 14792 17814
rect 14740 17750 14792 17756
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14660 16726 14688 17682
rect 14752 17338 14780 17750
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14844 17066 14872 17614
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14844 16794 14872 17002
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 15304 16726 15332 17478
rect 15474 16960 15530 16969
rect 15580 16946 15608 24618
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 15672 24070 15700 24101
rect 15660 24064 15712 24070
rect 15658 24032 15660 24041
rect 15712 24032 15714 24041
rect 15658 23967 15714 23976
rect 15672 23730 15700 23967
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15672 23322 15700 23666
rect 16040 23526 16068 24210
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 16132 23866 16160 24142
rect 16316 23866 16344 24346
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16118 23760 16174 23769
rect 16118 23695 16174 23704
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15672 22642 15700 23258
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15856 22778 15884 23054
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15948 22030 15976 23190
rect 15660 22024 15712 22030
rect 15844 22024 15896 22030
rect 15712 21984 15792 22012
rect 15660 21966 15712 21972
rect 15764 21350 15792 21984
rect 15844 21966 15896 21972
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15856 21690 15884 21966
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 15672 20505 15700 20946
rect 15658 20496 15714 20505
rect 15658 20431 15714 20440
rect 15764 20346 15792 21286
rect 15856 20942 15884 21490
rect 15948 21146 15976 21966
rect 16040 21962 16068 23462
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 16026 21856 16082 21865
rect 16026 21791 16082 21800
rect 16040 21690 16068 21791
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15856 20602 15884 20878
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15672 20318 15792 20346
rect 15672 17746 15700 20318
rect 15750 20088 15806 20097
rect 15750 20023 15806 20032
rect 15764 19394 15792 20023
rect 15856 19990 15884 20538
rect 16040 20097 16068 21626
rect 16026 20088 16082 20097
rect 16026 20023 16082 20032
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15856 19514 15884 19926
rect 15934 19816 15990 19825
rect 15934 19751 15990 19760
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15764 19366 15884 19394
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15764 18426 15792 19178
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15672 17513 15700 17682
rect 15658 17504 15714 17513
rect 15658 17439 15714 17448
rect 15530 16918 15608 16946
rect 15474 16895 15530 16904
rect 14648 16720 14700 16726
rect 15292 16720 15344 16726
rect 14700 16668 14872 16674
rect 14648 16662 14872 16668
rect 15292 16662 15344 16668
rect 14660 16646 14872 16662
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14660 16046 14688 16526
rect 14752 16250 14780 16526
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14738 16144 14794 16153
rect 14844 16114 14872 16646
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16130 15332 16662
rect 15580 16561 15608 16918
rect 15672 16794 15700 17439
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15764 16590 15792 18362
rect 15856 16794 15884 19366
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15752 16584 15804 16590
rect 15566 16552 15622 16561
rect 15752 16526 15804 16532
rect 15566 16487 15622 16496
rect 15764 16250 15792 16526
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 14738 16079 14794 16088
rect 14832 16108 14884 16114
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14660 15706 14688 15982
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14660 14074 14688 14418
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14476 12782 14504 13126
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14660 11898 14688 13126
rect 14648 11892 14700 11898
rect 14292 11750 14412 11778
rect 14568 11852 14648 11880
rect 14108 11206 14228 11234
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14108 10198 14136 11086
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14200 7970 14228 11206
rect 14292 10266 14320 11750
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14476 10810 14504 11222
rect 14568 11150 14596 11852
rect 14648 11834 14700 11840
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14660 11354 14688 11562
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14660 10674 14688 11290
rect 14752 11286 14780 16079
rect 14832 16050 14884 16056
rect 15120 16102 15332 16130
rect 15120 15706 15148 16102
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 15745 15240 15846
rect 15198 15736 15254 15745
rect 15108 15700 15160 15706
rect 15198 15671 15254 15680
rect 15108 15642 15160 15648
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 15106 15464 15162 15473
rect 14844 15162 14872 15438
rect 15106 15399 15108 15408
rect 15160 15399 15162 15408
rect 15108 15370 15160 15376
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15212 14618 15240 14758
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15304 14550 15332 15302
rect 15764 15201 15792 15506
rect 15750 15192 15806 15201
rect 15750 15127 15752 15136
rect 15804 15127 15806 15136
rect 15752 15098 15804 15104
rect 15764 14793 15792 15098
rect 15750 14784 15806 14793
rect 15750 14719 15806 14728
rect 15474 14648 15530 14657
rect 15474 14583 15530 14592
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15488 13682 15516 14583
rect 15568 13864 15620 13870
rect 15566 13832 15568 13841
rect 15620 13832 15622 13841
rect 15566 13767 15622 13776
rect 15948 13734 15976 19751
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16040 18426 16068 18702
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16026 17368 16082 17377
rect 16026 17303 16082 17312
rect 16040 17134 16068 17303
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 16132 15978 16160 23695
rect 16302 23624 16358 23633
rect 16302 23559 16358 23568
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 16224 19174 16252 19858
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16316 18601 16344 23559
rect 16408 23254 16436 24754
rect 16684 24614 16712 25298
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16500 23338 16528 24142
rect 17038 23896 17094 23905
rect 17038 23831 17040 23840
rect 17092 23831 17094 23840
rect 17040 23802 17092 23808
rect 17038 23488 17094 23497
rect 17038 23423 17094 23432
rect 16500 23322 16620 23338
rect 16500 23316 16632 23322
rect 16500 23310 16580 23316
rect 16580 23258 16632 23264
rect 16396 23248 16448 23254
rect 16396 23190 16448 23196
rect 16408 22778 16436 23190
rect 17052 22778 17080 23423
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 16486 22672 16542 22681
rect 16486 22607 16542 22616
rect 16500 22250 16528 22607
rect 16500 22222 16620 22250
rect 16592 22012 16620 22222
rect 16672 22024 16724 22030
rect 16592 21984 16672 22012
rect 16396 21888 16448 21894
rect 16396 21830 16448 21836
rect 16408 21486 16436 21830
rect 16592 21554 16620 21984
rect 16672 21966 16724 21972
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16302 18592 16358 18601
rect 16302 18527 16358 18536
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16316 17338 16344 17614
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16408 17218 16436 21422
rect 16960 21146 16988 21830
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 17052 20806 17080 21286
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16580 20528 16632 20534
rect 16578 20496 16580 20505
rect 16632 20496 16634 20505
rect 16578 20431 16634 20440
rect 17052 20330 17080 20742
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16592 18222 16620 18566
rect 16684 18358 16712 18838
rect 16776 18426 16804 19654
rect 17144 19242 17172 24550
rect 17328 21690 17356 27520
rect 17972 25498 18000 27520
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18432 24750 18460 25230
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 17500 24676 17552 24682
rect 17500 24618 17552 24624
rect 17512 22778 17540 24618
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17788 23769 17816 24006
rect 17774 23760 17830 23769
rect 17774 23695 17830 23704
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17788 22778 17816 23258
rect 18064 22778 18092 24210
rect 18142 23624 18198 23633
rect 18142 23559 18198 23568
rect 18156 23322 18184 23559
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17776 22772 17828 22778
rect 17776 22714 17828 22720
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17512 22574 17540 22714
rect 18156 22642 18184 23258
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 18340 22574 18368 24550
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 18432 23594 18460 24142
rect 18420 23588 18472 23594
rect 18420 23530 18472 23536
rect 18616 23526 18644 24210
rect 18604 23520 18656 23526
rect 18708 23497 18736 27520
rect 19352 25514 19380 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19352 25486 19472 25514
rect 20088 25498 20116 27520
rect 19340 25356 19392 25362
rect 19340 25298 19392 25304
rect 18880 24948 18932 24954
rect 18880 24890 18932 24896
rect 18604 23462 18656 23468
rect 18694 23488 18750 23497
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 17500 22568 17552 22574
rect 17406 22536 17462 22545
rect 17500 22510 17552 22516
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 17406 22471 17462 22480
rect 17420 22234 17448 22471
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17420 21418 17448 22170
rect 17408 21412 17460 21418
rect 17408 21354 17460 21360
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16960 18766 16988 19110
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16580 18216 16632 18222
rect 16316 17190 16436 17218
rect 16500 18164 16580 18170
rect 16500 18158 16632 18164
rect 16500 18142 16620 18158
rect 16960 18154 16988 18702
rect 16948 18148 17000 18154
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16210 15600 16266 15609
rect 16210 15535 16266 15544
rect 16224 15502 16252 15535
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16224 14890 16252 15438
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16132 13870 16160 14554
rect 16224 14550 16252 14826
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 15936 13728 15988 13734
rect 15488 13654 15608 13682
rect 15936 13670 15988 13676
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14844 12714 14872 13466
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15488 12238 15516 12582
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11898 15332 12038
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15488 11393 15516 12038
rect 15474 11384 15530 11393
rect 15474 11319 15530 11328
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14568 10470 14596 10542
rect 14556 10464 14608 10470
rect 14554 10432 14556 10441
rect 14608 10432 14610 10441
rect 14554 10367 14610 10376
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14462 10160 14518 10169
rect 14280 10124 14332 10130
rect 14752 10130 14780 10950
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10266 15332 11154
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14462 10095 14518 10104
rect 14740 10124 14792 10130
rect 14280 10066 14332 10072
rect 14292 9178 14320 10066
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14108 7942 14228 7970
rect 14108 5273 14136 7942
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14200 7410 14228 7822
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14200 6662 14228 7346
rect 14188 6656 14240 6662
rect 14186 6624 14188 6633
rect 14240 6624 14242 6633
rect 14242 6582 14320 6610
rect 14186 6559 14242 6568
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14094 5264 14150 5273
rect 14094 5199 14150 5208
rect 14108 3738 14136 5199
rect 14200 5098 14228 6122
rect 14292 5370 14320 6582
rect 14476 6361 14504 10095
rect 14740 10066 14792 10072
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 8838 14780 9454
rect 14844 9432 14872 9862
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14924 9444 14976 9450
rect 14844 9404 14924 9432
rect 14924 9386 14976 9392
rect 14936 9178 14964 9386
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 8430 14780 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14752 8090 14780 8366
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14752 6458 14780 8026
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15108 7336 15160 7342
rect 15304 7324 15332 10066
rect 15396 9926 15424 11086
rect 15488 10577 15516 11319
rect 15474 10568 15530 10577
rect 15580 10554 15608 13654
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15856 12986 15884 13330
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15672 11898 15700 12174
rect 16040 12102 16068 13262
rect 16316 12986 16344 17190
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16408 15570 16436 15846
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16500 15450 16528 18142
rect 16948 18090 17000 18096
rect 16854 17776 16910 17785
rect 16854 17711 16910 17720
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16776 16153 16804 16526
rect 16762 16144 16818 16153
rect 16762 16079 16818 16088
rect 16776 16046 16804 16079
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16408 15422 16528 15450
rect 16408 15162 16436 15422
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16500 15042 16528 15302
rect 16500 15026 16620 15042
rect 16500 15020 16632 15026
rect 16500 15014 16580 15020
rect 16580 14962 16632 14968
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16408 13938 16436 14486
rect 16592 14074 16620 14758
rect 16868 14600 16896 17711
rect 16960 17678 16988 18090
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16960 16998 16988 17614
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16658 16988 16934
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 16960 15910 16988 16594
rect 17144 16182 17172 16594
rect 17236 16425 17264 18022
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17420 17134 17448 17750
rect 17408 17128 17460 17134
rect 17406 17096 17408 17105
rect 17460 17096 17462 17105
rect 17406 17031 17462 17040
rect 17222 16416 17278 16425
rect 17222 16351 17278 16360
rect 17132 16176 17184 16182
rect 17052 16136 17132 16164
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16960 15502 16988 15846
rect 17052 15706 17080 16136
rect 17132 16118 17184 16124
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16960 14822 16988 15438
rect 17420 14958 17448 15506
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16776 14572 16896 14600
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16408 13818 16436 13874
rect 16408 13790 16620 13818
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16224 12345 16252 12922
rect 16210 12336 16266 12345
rect 16210 12271 16266 12280
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15672 11082 15700 11834
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11354 15792 11494
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 16316 11082 16344 11698
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 15752 10600 15804 10606
rect 15580 10526 15700 10554
rect 15752 10542 15804 10548
rect 15842 10568 15898 10577
rect 15474 10503 15530 10512
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10198 15608 10406
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15566 9888 15622 9897
rect 15566 9823 15622 9832
rect 15580 7993 15608 9823
rect 15566 7984 15622 7993
rect 15566 7919 15622 7928
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15160 7296 15332 7324
rect 15108 7278 15160 7284
rect 15290 6760 15346 6769
rect 15290 6695 15346 6704
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14462 6352 14518 6361
rect 14462 6287 14518 6296
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14200 4826 14228 5034
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14476 4434 14504 6287
rect 14752 5166 14780 6394
rect 15304 5642 15332 6695
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14646 4856 14702 4865
rect 15120 4826 15148 5238
rect 14646 4791 14702 4800
rect 15108 4820 15160 4826
rect 14660 4593 14688 4791
rect 15108 4762 15160 4768
rect 14646 4584 14702 4593
rect 14646 4519 14702 4528
rect 14740 4480 14792 4486
rect 14476 4406 14688 4434
rect 14740 4422 14792 4428
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 13634 3496 13690 3505
rect 13634 3431 13636 3440
rect 13688 3431 13690 3440
rect 13832 3488 14044 3516
rect 13636 3402 13688 3408
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13464 2990 13492 3130
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13634 2952 13690 2961
rect 13634 2887 13690 2896
rect 13648 2854 13676 2887
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13082 2680 13138 2689
rect 13832 2666 13860 3488
rect 14108 3058 14136 3674
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14200 3194 14228 3538
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14568 3058 14596 3606
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14554 2816 14610 2825
rect 14554 2751 14610 2760
rect 13832 2638 13952 2666
rect 13082 2615 13084 2624
rect 13136 2615 13138 2624
rect 13084 2586 13136 2592
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13372 2009 13400 2246
rect 13358 2000 13414 2009
rect 13358 1935 13414 1944
rect 12808 604 12860 610
rect 12808 546 12860 552
rect 13176 604 13228 610
rect 13176 546 13228 552
rect 13188 480 13216 546
rect 13924 480 13952 2638
rect 14462 2408 14518 2417
rect 14462 2343 14464 2352
rect 14516 2343 14518 2352
rect 14464 2314 14516 2320
rect 14568 480 14596 2751
rect 14660 2514 14688 4406
rect 14752 4049 14780 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15396 4185 15424 6598
rect 15488 4690 15516 7482
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15580 6186 15608 6666
rect 15568 6180 15620 6186
rect 15568 6122 15620 6128
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15488 4282 15516 4626
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15382 4176 15438 4185
rect 15382 4111 15438 4120
rect 14738 4040 14794 4049
rect 14738 3975 14794 3984
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14844 3534 14872 3878
rect 15672 3602 15700 10526
rect 15764 9654 15792 10542
rect 15842 10503 15898 10512
rect 15856 9994 15884 10503
rect 16224 10266 16252 10610
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 16132 9738 16160 10134
rect 16224 10062 16252 10202
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 15948 9722 16160 9738
rect 16224 9722 16252 9998
rect 15936 9716 16160 9722
rect 15988 9710 16160 9716
rect 15936 9658 15988 9664
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15764 5760 15792 9454
rect 15844 7472 15896 7478
rect 15844 7414 15896 7420
rect 15856 6798 15884 7414
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 5914 15884 6734
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15844 5772 15896 5778
rect 15764 5732 15844 5760
rect 15844 5714 15896 5720
rect 15856 4486 15884 5714
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15948 5370 15976 5646
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 16040 4729 16068 9522
rect 16132 8922 16160 9710
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16224 9110 16252 9658
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16316 9042 16344 11018
rect 16408 9722 16436 13670
rect 16592 13462 16620 13790
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16684 12782 16712 13194
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 11880 16620 12582
rect 16500 11852 16620 11880
rect 16500 11694 16528 11852
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16500 9738 16528 10474
rect 16592 10266 16620 11154
rect 16684 11082 16712 11494
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16396 9716 16448 9722
rect 16500 9710 16620 9738
rect 16396 9658 16448 9664
rect 16592 9654 16620 9710
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16132 8894 16252 8922
rect 16224 6361 16252 8894
rect 16316 8294 16344 8978
rect 16580 8900 16632 8906
rect 16500 8860 16580 8888
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 8022 16344 8230
rect 16500 8090 16528 8860
rect 16580 8842 16632 8848
rect 16684 8090 16712 11018
rect 16776 10742 16804 14572
rect 16856 14476 16908 14482
rect 16960 14464 16988 14758
rect 17420 14618 17448 14894
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 16908 14436 16988 14464
rect 16856 14418 16908 14424
rect 16960 13870 16988 14436
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16960 11558 16988 13806
rect 17038 13288 17094 13297
rect 17038 13223 17094 13232
rect 17052 12442 17080 13223
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11150 16988 11494
rect 17052 11286 17080 12378
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17144 11898 17172 12242
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16960 10810 16988 11086
rect 17052 10810 17080 11222
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16764 10736 16816 10742
rect 16764 10678 16816 10684
rect 17512 10441 17540 22510
rect 18432 22234 18460 22646
rect 18420 22228 18472 22234
rect 18420 22170 18472 22176
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 18420 22024 18472 22030
rect 18524 22001 18552 22170
rect 18420 21966 18472 21972
rect 18510 21992 18566 22001
rect 17592 21888 17644 21894
rect 17592 21830 17644 21836
rect 17604 21078 17632 21830
rect 17696 21350 17724 21966
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17868 21412 17920 21418
rect 17868 21354 17920 21360
rect 17684 21344 17736 21350
rect 17684 21286 17736 21292
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17592 21072 17644 21078
rect 17592 21014 17644 21020
rect 17696 20058 17724 21082
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17696 18426 17724 18770
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17604 12102 17632 13398
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17788 12782 17816 13262
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17604 11801 17632 12038
rect 17590 11792 17646 11801
rect 17590 11727 17646 11736
rect 17498 10432 17554 10441
rect 17498 10367 17554 10376
rect 16762 10160 16818 10169
rect 16762 10095 16764 10104
rect 16816 10095 16818 10104
rect 17224 10124 17276 10130
rect 16764 10066 16816 10072
rect 17224 10066 17276 10072
rect 16776 9586 16804 10066
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16960 9382 16988 9998
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7410 16528 7686
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16500 7002 16528 7346
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16408 6746 16436 6870
rect 16408 6718 16620 6746
rect 16488 6656 16540 6662
rect 16486 6624 16488 6633
rect 16540 6624 16542 6633
rect 16486 6559 16542 6568
rect 16210 6352 16266 6361
rect 16210 6287 16266 6296
rect 16224 5846 16252 6287
rect 16500 6254 16528 6559
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 16224 5370 16252 5782
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16026 4720 16082 4729
rect 16026 4655 16082 4664
rect 16592 4486 16620 6718
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16684 5710 16712 6122
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16684 5030 16712 5646
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 15660 3596 15712 3602
rect 15712 3556 15792 3584
rect 15660 3538 15712 3544
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 14844 3398 14872 3470
rect 14832 3392 14884 3398
rect 15396 3369 15424 3470
rect 15476 3392 15528 3398
rect 14832 3334 14884 3340
rect 15382 3360 15438 3369
rect 14738 3224 14794 3233
rect 14738 3159 14794 3168
rect 14752 2650 14780 3159
rect 14844 2922 14872 3334
rect 14956 3292 15252 3312
rect 15476 3334 15528 3340
rect 15382 3295 15438 3304
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15488 3233 15516 3334
rect 15474 3224 15530 3233
rect 15474 3159 15530 3168
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14844 2582 14872 2858
rect 15764 2825 15792 3556
rect 15750 2816 15806 2825
rect 15750 2751 15806 2760
rect 15764 2582 15792 2751
rect 14832 2576 14884 2582
rect 14830 2544 14832 2553
rect 15752 2576 15804 2582
rect 14884 2544 14886 2553
rect 14648 2508 14700 2514
rect 15752 2518 15804 2524
rect 14830 2479 14886 2488
rect 14648 2450 14700 2456
rect 14844 2453 14872 2479
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15856 1465 15884 4422
rect 16040 4185 16068 4422
rect 16684 4298 16712 4966
rect 16776 4865 16804 9318
rect 17052 8974 17080 9005
rect 17040 8968 17092 8974
rect 17038 8936 17040 8945
rect 17092 8936 17094 8945
rect 17236 8906 17264 10066
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17420 9042 17448 9998
rect 17696 9738 17724 12038
rect 17788 11914 17816 12718
rect 17880 12102 17908 21354
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17972 17649 18000 21286
rect 18064 20466 18092 21490
rect 18432 21350 18460 21966
rect 18510 21927 18566 21936
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 18064 18086 18092 20402
rect 18432 20058 18460 20742
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18156 19310 18184 19654
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18512 19168 18564 19174
rect 18616 19145 18644 23462
rect 18694 23423 18750 23432
rect 18892 22234 18920 24890
rect 19352 24614 19380 25298
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 18972 24064 19024 24070
rect 18972 24006 19024 24012
rect 18984 23662 19012 24006
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 18984 23186 19012 23598
rect 18972 23180 19024 23186
rect 18972 23122 19024 23128
rect 18984 22438 19012 23122
rect 19154 22536 19210 22545
rect 19154 22471 19210 22480
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18880 22228 18932 22234
rect 18880 22170 18932 22176
rect 18892 21146 18920 22170
rect 18984 21690 19012 22374
rect 19168 21962 19196 22471
rect 19352 22114 19380 24550
rect 19444 23905 19472 25486
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20166 24848 20222 24857
rect 20166 24783 20222 24792
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19430 23896 19486 23905
rect 19430 23831 19486 23840
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 19444 23322 19472 23530
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19260 22086 19380 22114
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 18972 21684 19024 21690
rect 18972 21626 19024 21632
rect 18880 21140 18932 21146
rect 18880 21082 18932 21088
rect 19156 21004 19208 21010
rect 19156 20946 19208 20952
rect 18788 20800 18840 20806
rect 18786 20768 18788 20777
rect 18840 20768 18842 20777
rect 18786 20703 18842 20712
rect 18696 20324 18748 20330
rect 18696 20266 18748 20272
rect 18708 19417 18736 20266
rect 19168 20058 19196 20946
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18984 19446 19012 19858
rect 18972 19440 19024 19446
rect 18694 19408 18750 19417
rect 18972 19382 19024 19388
rect 18694 19343 18696 19352
rect 18748 19343 18750 19352
rect 18696 19314 18748 19320
rect 18512 19110 18564 19116
rect 18602 19136 18658 19145
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17958 17640 18014 17649
rect 17958 17575 18014 17584
rect 17972 13870 18000 17575
rect 18248 16697 18276 18022
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18234 16688 18290 16697
rect 18340 16658 18368 17478
rect 18234 16623 18290 16632
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 18248 15609 18276 16390
rect 18234 15600 18290 15609
rect 18234 15535 18290 15544
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18064 14074 18092 14350
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17972 13530 18000 13806
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18064 12170 18092 12718
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18144 12368 18196 12374
rect 18142 12336 18144 12345
rect 18196 12336 18198 12345
rect 18142 12271 18198 12280
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17788 11898 18000 11914
rect 17788 11892 18012 11898
rect 17788 11886 17960 11892
rect 17960 11834 18012 11840
rect 18248 11626 18276 12038
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18248 11393 18276 11562
rect 18234 11384 18290 11393
rect 18234 11319 18236 11328
rect 18288 11319 18290 11328
rect 18236 11290 18288 11296
rect 18050 11112 18106 11121
rect 18050 11047 18106 11056
rect 17774 10840 17830 10849
rect 17774 10775 17830 10784
rect 17788 10130 17816 10775
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17604 9710 17724 9738
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17038 8871 17094 8880
rect 17224 8900 17276 8906
rect 17052 8634 17080 8871
rect 17224 8842 17276 8848
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16868 6474 16896 7482
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16960 6633 16988 7346
rect 17052 7342 17080 8026
rect 17236 7886 17264 8230
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17236 6934 17264 7822
rect 17314 7304 17370 7313
rect 17314 7239 17370 7248
rect 17328 7002 17356 7239
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 16946 6624 17002 6633
rect 16946 6559 17002 6568
rect 16868 6446 16988 6474
rect 17328 6458 17356 6938
rect 16854 5264 16910 5273
rect 16854 5199 16910 5208
rect 16868 5166 16896 5199
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16762 4856 16818 4865
rect 16762 4791 16818 4800
rect 16592 4270 16712 4298
rect 16026 4176 16082 4185
rect 16592 4162 16620 4270
rect 16026 4111 16082 4120
rect 16500 4134 16620 4162
rect 16672 4140 16724 4146
rect 16212 4004 16264 4010
rect 16212 3946 16264 3952
rect 16118 3632 16174 3641
rect 16224 3618 16252 3946
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16174 3590 16252 3618
rect 16118 3567 16120 3576
rect 16172 3567 16174 3576
rect 16120 3538 16172 3544
rect 15934 3088 15990 3097
rect 15934 3023 15990 3032
rect 15290 1456 15346 1465
rect 15290 1391 15346 1400
rect 15842 1456 15898 1465
rect 15842 1391 15898 1400
rect 15304 480 15332 1391
rect 15948 480 15976 3023
rect 16118 2680 16174 2689
rect 16118 2615 16120 2624
rect 16172 2615 16174 2624
rect 16120 2586 16172 2592
rect 16316 2582 16344 3878
rect 16500 3602 16528 4134
rect 16672 4082 16724 4088
rect 16580 4072 16632 4078
rect 16578 4040 16580 4049
rect 16632 4040 16634 4049
rect 16578 3975 16634 3984
rect 16578 3768 16634 3777
rect 16578 3703 16634 3712
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16500 3194 16528 3538
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16500 3058 16528 3130
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16592 2938 16620 3703
rect 16684 3602 16712 4082
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16684 3126 16712 3538
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 16592 2910 16712 2938
rect 16684 2666 16712 2910
rect 16592 2638 16712 2666
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 16592 480 16620 2638
rect 16960 2145 16988 6446
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 17052 4321 17080 4966
rect 17512 4758 17540 9590
rect 17604 6934 17632 9710
rect 17880 9654 17908 10134
rect 17958 10024 18014 10033
rect 17958 9959 18014 9968
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17696 8090 17724 9522
rect 17774 9344 17830 9353
rect 17774 9279 17830 9288
rect 17788 9178 17816 9279
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17696 7206 17724 7890
rect 17788 7818 17816 8910
rect 17880 8634 17908 8978
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17880 7886 17908 8434
rect 17972 8090 18000 9959
rect 18064 9654 18092 11047
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18156 9450 18184 9862
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18248 9178 18276 9522
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18234 8664 18290 8673
rect 18340 8634 18368 12650
rect 18418 10704 18474 10713
rect 18418 10639 18474 10648
rect 18432 10266 18460 10639
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18524 9738 18552 19110
rect 18602 19071 18658 19080
rect 18616 18578 18644 19071
rect 18984 18970 19012 19382
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 19076 18902 19104 19926
rect 19260 19394 19288 22086
rect 19524 21888 19576 21894
rect 19524 21830 19576 21836
rect 19536 21486 19564 21830
rect 19524 21480 19576 21486
rect 19524 21422 19576 21428
rect 19536 21078 19564 21422
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19536 20602 19564 21014
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19536 19854 19564 20538
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19536 19514 19564 19790
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19168 19366 19288 19394
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 18616 18550 18828 18578
rect 18602 18456 18658 18465
rect 18602 18391 18604 18400
rect 18656 18391 18658 18400
rect 18604 18362 18656 18368
rect 18616 18222 18644 18362
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18696 15972 18748 15978
rect 18696 15914 18748 15920
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18616 14958 18644 15302
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18616 14618 18644 14894
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18616 13938 18644 14554
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18708 9761 18736 15914
rect 18800 10577 18828 18550
rect 19168 17626 19196 19366
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 18984 17598 19196 17626
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18892 12889 18920 13262
rect 18984 12918 19012 17598
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19062 17232 19118 17241
rect 19062 17167 19118 17176
rect 19076 17066 19104 17167
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 19076 16794 19104 17002
rect 19168 16998 19196 17478
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 19168 16250 19196 16934
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19168 16114 19196 16186
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19260 16046 19288 19246
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19430 18728 19486 18737
rect 19430 18663 19486 18672
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19352 17542 19380 18090
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19340 17060 19392 17066
rect 19340 17002 19392 17008
rect 19352 16969 19380 17002
rect 19338 16960 19394 16969
rect 19338 16895 19394 16904
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19062 14920 19118 14929
rect 19062 14855 19118 14864
rect 19076 14618 19104 14855
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 19168 14113 19196 15846
rect 19260 15706 19288 15982
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19444 15586 19472 18663
rect 19536 16794 19564 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19798 18864 19854 18873
rect 19798 18799 19800 18808
rect 19852 18799 19854 18808
rect 19800 18770 19852 18776
rect 19996 18714 20024 24686
rect 20180 24614 20208 24783
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 20732 24426 20760 27520
rect 21376 24857 21404 27520
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 22020 24886 22048 25298
rect 21456 24880 21508 24886
rect 21362 24848 21418 24857
rect 21180 24812 21232 24818
rect 21456 24822 21508 24828
rect 22008 24880 22060 24886
rect 22008 24822 22060 24828
rect 21362 24783 21418 24792
rect 21180 24754 21232 24760
rect 21088 24744 21140 24750
rect 21088 24686 21140 24692
rect 20640 24410 20760 24426
rect 20628 24404 20760 24410
rect 20680 24398 20760 24404
rect 20628 24346 20680 24352
rect 20904 24064 20956 24070
rect 20626 24032 20682 24041
rect 20904 24006 20956 24012
rect 20626 23967 20682 23976
rect 20534 23760 20590 23769
rect 20534 23695 20590 23704
rect 20260 22500 20312 22506
rect 20260 22442 20312 22448
rect 20074 22400 20130 22409
rect 20074 22335 20130 22344
rect 20088 18850 20116 22335
rect 20272 22234 20300 22442
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20272 21690 20300 22170
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20272 20942 20300 21626
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20272 20602 20300 20878
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20548 20754 20576 23695
rect 20640 23526 20668 23967
rect 20916 23633 20944 24006
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 20902 23624 20958 23633
rect 20902 23559 20958 23568
rect 20628 23520 20680 23526
rect 20680 23468 20852 23474
rect 20628 23462 20852 23468
rect 20640 23446 20852 23462
rect 20824 23118 20852 23446
rect 20812 23112 20864 23118
rect 20718 23080 20774 23089
rect 21008 23089 21036 23802
rect 20812 23054 20864 23060
rect 20994 23080 21050 23089
rect 20718 23015 20720 23024
rect 20772 23015 20774 23024
rect 20720 22986 20772 22992
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20732 21078 20760 22374
rect 20824 22234 20852 23054
rect 20994 23015 21050 23024
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 20904 21072 20956 21078
rect 20904 21014 20956 21020
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20456 20482 20484 20742
rect 20548 20726 20852 20754
rect 20456 20466 20760 20482
rect 20456 20460 20772 20466
rect 20456 20454 20720 20460
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20180 19174 20208 19654
rect 20272 19378 20300 19722
rect 20456 19417 20484 20454
rect 20720 20402 20772 20408
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20548 19990 20576 20198
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20640 19718 20668 20198
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 19417 20668 19654
rect 20442 19408 20498 19417
rect 20260 19372 20312 19378
rect 20442 19343 20498 19352
rect 20626 19408 20682 19417
rect 20626 19343 20682 19352
rect 20260 19314 20312 19320
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20088 18822 20208 18850
rect 19996 18686 20116 18714
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19996 18329 20024 18566
rect 19982 18320 20038 18329
rect 19982 18255 20038 18264
rect 20088 18034 20116 18686
rect 19996 18006 20116 18034
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19812 17649 19840 17682
rect 19798 17640 19854 17649
rect 19798 17575 19854 17584
rect 19996 17377 20024 18006
rect 20074 17912 20130 17921
rect 20074 17847 20076 17856
rect 20128 17847 20130 17856
rect 20076 17818 20128 17824
rect 20180 17785 20208 18822
rect 20166 17776 20222 17785
rect 20166 17711 20222 17720
rect 19982 17368 20038 17377
rect 19982 17303 20038 17312
rect 20272 17241 20300 19314
rect 20350 18864 20406 18873
rect 20350 18799 20406 18808
rect 20364 17882 20392 18799
rect 20456 18426 20484 19343
rect 20628 19168 20680 19174
rect 20680 19128 20760 19156
rect 20628 19110 20680 19116
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20732 17882 20760 19128
rect 20352 17876 20404 17882
rect 20352 17818 20404 17824
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20350 17640 20406 17649
rect 20350 17575 20406 17584
rect 20258 17232 20314 17241
rect 20258 17167 20314 17176
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20364 16794 20392 17575
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20534 16144 20590 16153
rect 20534 16079 20590 16088
rect 20548 15910 20576 16079
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19444 15558 19564 15586
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19444 14618 19472 15438
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19154 14104 19210 14113
rect 19154 14039 19210 14048
rect 19352 13938 19380 14282
rect 19444 14074 19472 14554
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 18972 12912 19024 12918
rect 18878 12880 18934 12889
rect 18972 12854 19024 12860
rect 18878 12815 18880 12824
rect 18932 12815 18934 12824
rect 18880 12786 18932 12792
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18984 11354 19012 11834
rect 19076 11694 19104 13806
rect 19352 13530 19380 13874
rect 19536 13530 19564 15558
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14346 20024 14758
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18786 10568 18842 10577
rect 18786 10503 18842 10512
rect 18892 10044 18920 10746
rect 18984 10588 19012 11290
rect 19064 10600 19116 10606
rect 18984 10560 19064 10588
rect 19064 10542 19116 10548
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 18972 10056 19024 10062
rect 18892 10016 18972 10044
rect 18432 9710 18552 9738
rect 18694 9752 18750 9761
rect 18234 8599 18290 8608
rect 18328 8628 18380 8634
rect 18248 8514 18276 8599
rect 18328 8570 18380 8576
rect 18248 8486 18368 8514
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17788 7546 17816 7754
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17880 7154 17908 7210
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17604 6458 17632 6870
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17604 5817 17632 6394
rect 17590 5808 17646 5817
rect 17590 5743 17646 5752
rect 17696 4758 17724 7142
rect 17880 7126 18000 7154
rect 17972 6730 18000 7126
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17774 6624 17830 6633
rect 17774 6559 17830 6568
rect 17788 5574 17816 6559
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17500 4752 17552 4758
rect 17420 4700 17500 4706
rect 17420 4694 17552 4700
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 17420 4678 17540 4694
rect 17038 4312 17094 4321
rect 17420 4282 17448 4678
rect 17788 4622 17816 5510
rect 17880 4826 17908 6054
rect 18156 4826 18184 8366
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18248 4826 18276 7278
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17776 4616 17828 4622
rect 18156 4604 18184 4762
rect 18156 4576 18276 4604
rect 17776 4558 17828 4564
rect 17038 4247 17094 4256
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 17144 2650 17172 3062
rect 17420 2854 17448 3334
rect 17512 3194 17540 4558
rect 18144 4208 18196 4214
rect 18064 4156 18144 4162
rect 18064 4150 18196 4156
rect 18064 4134 18184 4150
rect 18248 4146 18276 4576
rect 18236 4140 18288 4146
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17958 2952 18014 2961
rect 17958 2887 18014 2896
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17420 2446 17448 2790
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 16946 2136 17002 2145
rect 16946 2071 17002 2080
rect 17314 1592 17370 1601
rect 17314 1527 17370 1536
rect 17328 480 17356 1527
rect 17972 480 18000 2887
rect 18064 2582 18092 4134
rect 18236 4082 18288 4088
rect 18340 4078 18368 8486
rect 18432 8401 18460 9710
rect 18694 9687 18750 9696
rect 18510 9616 18566 9625
rect 18892 9586 18920 10016
rect 18972 9998 19024 10004
rect 18510 9551 18566 9560
rect 18880 9580 18932 9586
rect 18524 8430 18552 9551
rect 18880 9522 18932 9528
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8498 18736 8774
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18512 8424 18564 8430
rect 18418 8392 18474 8401
rect 18512 8366 18564 8372
rect 18418 8327 18420 8336
rect 18472 8327 18474 8336
rect 18420 8298 18472 8304
rect 18510 7984 18566 7993
rect 18510 7919 18512 7928
rect 18564 7919 18566 7928
rect 18512 7890 18564 7896
rect 18524 7546 18552 7890
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18616 7546 18644 7822
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18604 7540 18656 7546
rect 18656 7500 18736 7528
rect 18604 7482 18656 7488
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3058 18276 3878
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18052 2576 18104 2582
rect 18050 2544 18052 2553
rect 18104 2544 18106 2553
rect 18432 2514 18460 7142
rect 18616 6662 18644 7278
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18616 4593 18644 6598
rect 18602 4584 18658 4593
rect 18602 4519 18658 4528
rect 18708 4457 18736 7500
rect 18800 6798 18828 9386
rect 19076 9382 19104 10066
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 18892 6866 18920 9318
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18788 6792 18840 6798
rect 18892 6769 18920 6802
rect 19064 6792 19116 6798
rect 18788 6734 18840 6740
rect 18878 6760 18934 6769
rect 18800 6118 18828 6734
rect 19064 6734 19116 6740
rect 18878 6695 18934 6704
rect 18892 6458 18920 6695
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18694 4448 18750 4457
rect 18694 4383 18750 4392
rect 18694 4176 18750 4185
rect 18694 4111 18750 4120
rect 18050 2479 18106 2488
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18708 480 18736 4111
rect 18800 2553 18828 6054
rect 19076 5846 19104 6734
rect 19168 6225 19196 12582
rect 19248 12436 19300 12442
rect 19352 12424 19380 12786
rect 19536 12782 19564 13194
rect 19812 12986 19840 13262
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19812 12866 19840 12922
rect 19996 12866 20024 13670
rect 20088 13394 20116 15846
rect 20548 15706 20576 15846
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20732 15609 20760 17682
rect 20718 15600 20774 15609
rect 20718 15535 20774 15544
rect 20442 15192 20498 15201
rect 20442 15127 20498 15136
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20076 13388 20128 13394
rect 20076 13330 20128 13336
rect 20180 12986 20208 13466
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 19812 12838 20024 12866
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19300 12396 19380 12424
rect 19248 12378 19300 12384
rect 19246 10704 19302 10713
rect 19246 10639 19302 10648
rect 19260 10266 19288 10639
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19352 9081 19380 12396
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19444 11082 19472 12174
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19536 10266 19564 12242
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 9178 20024 12838
rect 20258 12336 20314 12345
rect 20258 12271 20314 12280
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20088 11558 20116 12174
rect 20076 11552 20128 11558
rect 20074 11520 20076 11529
rect 20128 11520 20130 11529
rect 20074 11455 20130 11464
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20180 10470 20208 10950
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20074 10296 20130 10305
rect 20074 10231 20130 10240
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19338 9072 19394 9081
rect 19338 9007 19394 9016
rect 19432 9036 19484 9042
rect 19352 8090 19380 9007
rect 19432 8978 19484 8984
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19352 7274 19380 8026
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19154 6216 19210 6225
rect 19154 6151 19210 6160
rect 19064 5840 19116 5846
rect 19062 5808 19064 5817
rect 19116 5808 19118 5817
rect 19062 5743 19118 5752
rect 18892 5302 18920 5333
rect 18880 5296 18932 5302
rect 18878 5264 18880 5273
rect 18932 5264 18934 5273
rect 18878 5199 18934 5208
rect 18892 5030 18920 5199
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18892 3738 18920 4762
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 2689 18920 3334
rect 18878 2680 18934 2689
rect 18878 2615 18934 2624
rect 18786 2544 18842 2553
rect 18786 2479 18842 2488
rect 18984 2446 19012 5034
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19076 4214 19104 4558
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 19168 4078 19196 4626
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19156 4072 19208 4078
rect 19154 4040 19156 4049
rect 19208 4040 19210 4049
rect 19154 3975 19210 3984
rect 19260 3738 19288 4490
rect 19338 4312 19394 4321
rect 19338 4247 19394 4256
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19156 3528 19208 3534
rect 19154 3496 19156 3505
rect 19208 3496 19210 3505
rect 19064 3460 19116 3466
rect 19154 3431 19210 3440
rect 19064 3402 19116 3408
rect 19076 2650 19104 3402
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 19352 480 19380 4247
rect 19444 2990 19472 8978
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19536 7857 19564 8910
rect 19996 8430 20024 9114
rect 20088 8673 20116 10231
rect 20180 9722 20208 10406
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20272 9636 20300 12271
rect 20456 10849 20484 15127
rect 20732 13705 20760 15535
rect 20824 15162 20852 20726
rect 20916 19922 20944 21014
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20916 19514 20944 19858
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20916 17746 20944 19314
rect 21008 17882 21036 23015
rect 21100 22953 21128 24686
rect 21192 24206 21220 24754
rect 21270 24712 21326 24721
rect 21270 24647 21326 24656
rect 21284 24614 21312 24647
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21272 24268 21324 24274
rect 21272 24210 21324 24216
rect 21180 24200 21232 24206
rect 21180 24142 21232 24148
rect 21192 23526 21220 24142
rect 21284 23866 21312 24210
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 21086 22944 21142 22953
rect 21086 22879 21142 22888
rect 21192 22080 21220 23462
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21284 22642 21312 23122
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21284 22522 21312 22578
rect 21284 22494 21404 22522
rect 21192 22052 21312 22080
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 21100 21332 21128 21898
rect 21180 21344 21232 21350
rect 21100 21304 21180 21332
rect 21180 21286 21232 21292
rect 21088 19984 21140 19990
rect 21088 19926 21140 19932
rect 21100 18698 21128 19926
rect 21192 19446 21220 21286
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21284 19258 21312 22052
rect 21376 20262 21404 22494
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21192 18970 21220 19246
rect 21284 19230 21404 19258
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 21192 18306 21220 18702
rect 21284 18465 21312 19110
rect 21270 18456 21326 18465
rect 21270 18391 21326 18400
rect 21192 18278 21312 18306
rect 21284 18086 21312 18278
rect 21376 18154 21404 19230
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 20916 16658 20944 17070
rect 21008 16794 21036 17818
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21100 16726 21128 17478
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20916 16250 20944 16594
rect 21100 16454 21128 16662
rect 21088 16448 21140 16454
rect 20994 16416 21050 16425
rect 21088 16390 21140 16396
rect 20994 16351 21050 16360
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20824 14958 20852 15098
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20916 14482 20944 14758
rect 21008 14550 21036 16351
rect 21100 16114 21128 16390
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 21192 16046 21220 16934
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21192 15706 21220 15982
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21284 15201 21312 18022
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21376 17066 21404 17682
rect 21364 17060 21416 17066
rect 21364 17002 21416 17008
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21270 15192 21326 15201
rect 21270 15127 21326 15136
rect 21376 14929 21404 15506
rect 21362 14920 21418 14929
rect 21362 14855 21364 14864
rect 21416 14855 21418 14864
rect 21364 14826 21416 14832
rect 20996 14544 21048 14550
rect 20996 14486 21048 14492
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20916 14074 20944 14418
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 21100 13841 21128 14214
rect 21086 13832 21142 13841
rect 21086 13767 21142 13776
rect 20996 13728 21048 13734
rect 20718 13696 20774 13705
rect 20996 13670 21048 13676
rect 20718 13631 20774 13640
rect 21008 13258 21036 13670
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20732 12782 20760 13126
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20810 12744 20866 12753
rect 20916 12714 20944 13126
rect 21100 12782 21128 13330
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21376 12986 21404 13262
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20810 12679 20866 12688
rect 20904 12708 20956 12714
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 12306 20576 12582
rect 20824 12442 20852 12679
rect 20904 12650 20956 12656
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20628 11620 20680 11626
rect 20548 11580 20628 11608
rect 20548 11150 20576 11580
rect 20628 11562 20680 11568
rect 20732 11558 20760 12174
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20548 11014 20576 11086
rect 20732 11082 20760 11494
rect 21008 11354 21036 12582
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20536 11008 20588 11014
rect 20536 10950 20588 10956
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20442 10840 20498 10849
rect 20442 10775 20498 10784
rect 20810 10568 20866 10577
rect 20810 10503 20812 10512
rect 20864 10503 20866 10512
rect 20812 10474 20864 10480
rect 20916 10266 20944 10950
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20272 9608 20392 9636
rect 20074 8664 20130 8673
rect 20074 8599 20130 8608
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 20074 8392 20130 8401
rect 20074 8327 20130 8336
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19996 8072 20024 8230
rect 19904 8044 20024 8072
rect 19522 7848 19578 7857
rect 19904 7818 19932 8044
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19522 7783 19578 7792
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19536 6254 19564 7278
rect 19904 7274 19932 7754
rect 19892 7268 19944 7274
rect 19892 7210 19944 7216
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19536 5914 19564 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19536 5030 19564 5170
rect 19996 5166 20024 7822
rect 20088 6866 20116 8327
rect 20166 7848 20222 7857
rect 20166 7783 20222 7792
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20088 5778 20116 6802
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 20180 5370 20208 7783
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19536 4486 19564 4966
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4826 20024 5102
rect 20180 5098 20208 5306
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 20074 4856 20130 4865
rect 19984 4820 20036 4826
rect 20074 4791 20130 4800
rect 19984 4762 20036 4768
rect 20088 4758 20116 4791
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19536 3738 19564 4082
rect 19628 4078 19656 4558
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 19996 4010 20024 4422
rect 19984 4004 20036 4010
rect 19984 3946 20036 3952
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19522 3360 19578 3369
rect 19522 3295 19578 3304
rect 19432 2984 19484 2990
rect 19536 2961 19564 3295
rect 19432 2926 19484 2932
rect 19522 2952 19578 2961
rect 19522 2887 19578 2896
rect 19628 2836 19656 3470
rect 19996 3058 20024 3946
rect 20272 3097 20300 5510
rect 20364 5273 20392 9608
rect 21100 9518 21128 12718
rect 21192 9518 21220 12922
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21284 12442 21312 12582
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21284 10266 21312 11154
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21376 10146 21404 12038
rect 21468 11354 21496 24822
rect 21732 24744 21784 24750
rect 21732 24686 21784 24692
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21560 18970 21588 23462
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21652 22234 21680 23258
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 21652 20398 21680 22170
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21744 20210 21772 24686
rect 21824 24676 21876 24682
rect 21824 24618 21876 24624
rect 21836 24206 21864 24618
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21836 23526 21864 24142
rect 21824 23520 21876 23526
rect 22112 23508 22140 27520
rect 22756 25498 22784 27520
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22650 24168 22706 24177
rect 22650 24103 22706 24112
rect 22664 23866 22692 24103
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 21824 23462 21876 23468
rect 21928 23480 22140 23508
rect 23112 23520 23164 23526
rect 21836 22778 21864 23462
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 21928 21962 21956 23480
rect 23112 23462 23164 23468
rect 22742 23352 22798 23361
rect 22742 23287 22798 23296
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22100 22092 22152 22098
rect 22100 22034 22152 22040
rect 21916 21956 21968 21962
rect 21916 21898 21968 21904
rect 22112 21690 22140 22034
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 22112 21146 22140 21626
rect 22388 21486 22416 21966
rect 22480 21554 22508 22918
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22558 21312 22614 21321
rect 22558 21247 22614 21256
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 21836 20602 21864 20946
rect 21914 20768 21970 20777
rect 21914 20703 21970 20712
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21652 20182 21772 20210
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 21560 18222 21588 18906
rect 21652 18766 21680 20182
rect 21822 19680 21878 19689
rect 21822 19615 21878 19624
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21744 18970 21772 19110
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21744 18426 21772 18906
rect 21732 18420 21784 18426
rect 21732 18362 21784 18368
rect 21548 18216 21600 18222
rect 21548 18158 21600 18164
rect 21836 18034 21864 19615
rect 21560 18006 21864 18034
rect 21560 15586 21588 18006
rect 21638 17504 21694 17513
rect 21638 17439 21694 17448
rect 21652 16998 21680 17439
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21836 16454 21864 17138
rect 21928 16640 21956 20703
rect 22112 20602 22140 20946
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22112 20058 22140 20538
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 22020 19310 22048 19654
rect 22112 19514 22140 19994
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22572 19394 22600 21247
rect 22480 19366 22600 19394
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22296 18834 22324 19110
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22296 18290 22324 18770
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22112 18193 22140 18226
rect 22098 18184 22154 18193
rect 22098 18119 22154 18128
rect 22112 17542 22140 18119
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 21928 16612 22048 16640
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21836 15706 21864 16050
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 21560 15558 21864 15586
rect 21928 15570 21956 16186
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21560 13433 21588 15302
rect 21546 13424 21602 13433
rect 21546 13359 21602 13368
rect 21548 13252 21600 13258
rect 21548 13194 21600 13200
rect 21560 12646 21588 13194
rect 21732 12844 21784 12850
rect 21732 12786 21784 12792
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21744 12374 21772 12786
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21744 11898 21772 12310
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21744 11558 21772 11834
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21284 10118 21404 10146
rect 21560 10130 21588 10406
rect 21548 10124 21600 10130
rect 21088 9512 21140 9518
rect 21086 9480 21088 9489
rect 21180 9512 21232 9518
rect 21140 9480 21142 9489
rect 21180 9454 21232 9460
rect 21086 9415 21142 9424
rect 21192 9353 21220 9454
rect 21178 9344 21234 9353
rect 21178 9279 21234 9288
rect 20994 9072 21050 9081
rect 20994 9007 21050 9016
rect 21178 9072 21234 9081
rect 21178 9007 21234 9016
rect 21008 8634 21036 9007
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 21100 8090 21128 8910
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 6254 20852 7142
rect 21192 6730 21220 9007
rect 21284 7177 21312 10118
rect 21548 10066 21600 10072
rect 21744 10062 21772 11494
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21376 9722 21404 9998
rect 21546 9752 21602 9761
rect 21364 9716 21416 9722
rect 21546 9687 21602 9696
rect 21364 9658 21416 9664
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21468 7546 21496 7890
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21468 7274 21496 7482
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 21270 7168 21326 7177
rect 21560 7154 21588 9687
rect 21744 9654 21772 9998
rect 21732 9648 21784 9654
rect 21732 9590 21784 9596
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21744 8566 21772 9046
rect 21732 8560 21784 8566
rect 21730 8528 21732 8537
rect 21784 8528 21786 8537
rect 21730 8463 21786 8472
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21270 7103 21326 7112
rect 21468 7126 21588 7154
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 21086 6352 21142 6361
rect 21086 6287 21142 6296
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20824 5710 20852 6190
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20916 5817 20944 6054
rect 21100 5817 21128 6287
rect 21362 6216 21418 6225
rect 21362 6151 21418 6160
rect 21376 5846 21404 6151
rect 21364 5840 21416 5846
rect 20902 5808 20958 5817
rect 20902 5743 20958 5752
rect 21086 5808 21142 5817
rect 21364 5782 21416 5788
rect 21086 5743 21142 5752
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 20812 5704 20864 5710
rect 21284 5681 21312 5714
rect 20812 5646 20864 5652
rect 21270 5672 21326 5681
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20350 5264 20406 5273
rect 20456 5234 20484 5510
rect 20824 5370 20852 5646
rect 21270 5607 21326 5616
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20720 5296 20772 5302
rect 20720 5238 20772 5244
rect 20350 5199 20406 5208
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20364 3194 20392 3334
rect 20442 3224 20498 3233
rect 20352 3188 20404 3194
rect 20442 3159 20498 3168
rect 20352 3130 20404 3136
rect 20258 3088 20314 3097
rect 19984 3052 20036 3058
rect 20258 3023 20314 3032
rect 19984 2994 20036 3000
rect 19536 2808 19656 2836
rect 19536 2650 19564 2808
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20364 2650 20392 3130
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 19892 2372 19944 2378
rect 19892 2314 19944 2320
rect 19904 1170 19932 2314
rect 19904 1142 20116 1170
rect 20088 480 20116 1142
rect 20456 610 20484 3159
rect 20548 2514 20576 4218
rect 20732 3738 20760 5238
rect 20916 4729 20944 5510
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 20902 4720 20958 4729
rect 21008 4690 21036 5170
rect 21284 4826 21312 5607
rect 21376 5370 21404 5782
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 20902 4655 20958 4664
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20902 4584 20958 4593
rect 20824 4214 20852 4558
rect 20902 4519 20958 4528
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20916 3466 20944 4519
rect 21008 4282 21036 4626
rect 21178 4448 21234 4457
rect 21100 4406 21178 4434
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 21100 2990 21128 4406
rect 21178 4383 21234 4392
rect 21468 3670 21496 7126
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21560 6118 21588 6734
rect 21652 6662 21680 7958
rect 21836 7800 21864 15558
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21928 15162 21956 15506
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21928 14822 21956 15098
rect 21916 14816 21968 14822
rect 21916 14758 21968 14764
rect 22020 12345 22048 16612
rect 22006 12336 22062 12345
rect 22006 12271 22062 12280
rect 22112 12102 22140 17478
rect 22282 17232 22338 17241
rect 22282 17167 22338 17176
rect 22296 16794 22324 17167
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22296 16114 22324 16730
rect 22284 16108 22336 16114
rect 22284 16050 22336 16056
rect 22192 15564 22244 15570
rect 22192 15506 22244 15512
rect 22204 15162 22232 15506
rect 22192 15156 22244 15162
rect 22244 15116 22324 15144
rect 22192 15098 22244 15104
rect 22190 14104 22246 14113
rect 22190 14039 22246 14048
rect 22204 13530 22232 14039
rect 22296 14006 22324 15116
rect 22480 14498 22508 19366
rect 22560 18148 22612 18154
rect 22560 18090 22612 18096
rect 22572 17338 22600 18090
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22572 17066 22600 17274
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22756 15162 22784 23287
rect 22926 23216 22982 23225
rect 22926 23151 22982 23160
rect 22940 23118 22968 23151
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 22940 22778 22968 23054
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 23124 22522 23152 23462
rect 23216 22642 23244 27639
rect 23478 27520 23534 28000
rect 24122 27520 24178 28000
rect 24766 27520 24822 28000
rect 25502 27520 25558 28000
rect 26146 27520 26202 28000
rect 26882 27520 26938 28000
rect 27526 27520 27582 28000
rect 23294 26616 23350 26625
rect 23294 26551 23350 26560
rect 23308 23322 23336 26551
rect 23492 24721 23520 27520
rect 23662 25936 23718 25945
rect 23662 25871 23718 25880
rect 23676 24886 23704 25871
rect 23664 24880 23716 24886
rect 23664 24822 23716 24828
rect 23754 24848 23810 24857
rect 23754 24783 23810 24792
rect 23478 24712 23534 24721
rect 23478 24647 23534 24656
rect 23662 24576 23718 24585
rect 23662 24511 23718 24520
rect 23676 24410 23704 24511
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23584 23322 23612 24142
rect 23662 23624 23718 23633
rect 23662 23559 23718 23568
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23308 22710 23336 23258
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23124 22494 23336 22522
rect 23308 22438 23336 22494
rect 23296 22432 23348 22438
rect 23294 22400 23296 22409
rect 23348 22400 23350 22409
rect 23294 22335 23350 22344
rect 23400 22234 23428 22578
rect 23676 22522 23704 23559
rect 23492 22494 23704 22522
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 23400 22098 23428 22170
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23124 21350 23152 21966
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23124 21078 23152 21286
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 22928 18692 22980 18698
rect 22928 18634 22980 18640
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22480 14470 22692 14498
rect 22284 14000 22336 14006
rect 22284 13942 22336 13948
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22572 13530 22600 13670
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22204 12782 22232 13466
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 21914 11384 21970 11393
rect 21914 11319 21970 11328
rect 21928 10606 21956 11319
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22020 10674 22048 11086
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 22204 10470 22232 11018
rect 22192 10464 22244 10470
rect 21914 10432 21970 10441
rect 22192 10406 22244 10412
rect 21914 10367 21970 10376
rect 21928 7886 21956 10367
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 22112 9586 22140 10066
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 22020 8974 22048 9318
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 22020 8634 22048 8910
rect 22296 8906 22324 10202
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21744 7772 21864 7800
rect 21744 7546 21772 7772
rect 22112 7750 22140 8366
rect 22100 7744 22152 7750
rect 21836 7704 22100 7732
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21744 6798 21772 7346
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21652 6458 21680 6598
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21548 6112 21600 6118
rect 21546 6080 21548 6089
rect 21600 6080 21602 6089
rect 21546 6015 21602 6024
rect 21744 5914 21772 6734
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21836 5370 21864 7704
rect 22100 7686 22152 7692
rect 22204 7410 22232 8774
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 22296 7478 22324 7958
rect 22388 7478 22416 8774
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22098 7168 22154 7177
rect 21916 6996 21968 7002
rect 21916 6938 21968 6944
rect 21928 6458 21956 6938
rect 22020 6905 22048 7142
rect 22098 7103 22154 7112
rect 22006 6896 22062 6905
rect 22006 6831 22062 6840
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 22020 5574 22048 6734
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 21638 5264 21694 5273
rect 21638 5199 21694 5208
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21376 3126 21404 3470
rect 21454 3224 21510 3233
rect 21454 3159 21510 3168
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 20824 2650 20852 2926
rect 21468 2922 21496 3159
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 21652 2514 21680 5199
rect 22020 4729 22048 5510
rect 22112 5250 22140 7103
rect 22204 7002 22232 7346
rect 22388 7342 22416 7414
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22192 6996 22244 7002
rect 22192 6938 22244 6944
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22204 6497 22232 6598
rect 22190 6488 22246 6497
rect 22190 6423 22246 6432
rect 22204 6322 22232 6423
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22480 5778 22508 12786
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22572 8401 22600 8502
rect 22558 8392 22614 8401
rect 22558 8327 22614 8336
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 22572 7818 22600 8230
rect 22664 7834 22692 14470
rect 22756 14414 22784 14758
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22756 14074 22784 14350
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22756 13870 22784 14010
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22940 13569 22968 18634
rect 23202 18592 23258 18601
rect 23202 18527 23258 18536
rect 23216 18426 23244 18527
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23308 17814 23336 21830
rect 23400 21146 23428 22034
rect 23492 21865 23520 22494
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23676 22166 23704 22374
rect 23664 22160 23716 22166
rect 23664 22102 23716 22108
rect 23478 21856 23534 21865
rect 23478 21791 23534 21800
rect 23768 21706 23796 24783
rect 24136 24614 24164 27520
rect 24214 27160 24270 27169
rect 24214 27095 24270 27104
rect 24124 24608 24176 24614
rect 24124 24550 24176 24556
rect 23938 24304 23994 24313
rect 23848 24268 23900 24274
rect 23938 24239 23994 24248
rect 24124 24268 24176 24274
rect 23848 24210 23900 24216
rect 23860 23526 23888 24210
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 23860 23361 23888 23462
rect 23846 23352 23902 23361
rect 23846 23287 23902 23296
rect 23848 23248 23900 23254
rect 23848 23190 23900 23196
rect 23860 22574 23888 23190
rect 23848 22568 23900 22574
rect 23952 22545 23980 24239
rect 24124 24210 24176 24216
rect 24136 23730 24164 24210
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 23848 22510 23900 22516
rect 23938 22536 23994 22545
rect 23938 22471 23994 22480
rect 23676 21678 23796 21706
rect 23388 21140 23440 21146
rect 23388 21082 23440 21088
rect 23572 21072 23624 21078
rect 23572 21014 23624 21020
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23492 20602 23520 20946
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23400 18034 23428 18702
rect 23492 18698 23520 20198
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23584 18154 23612 21014
rect 23676 19530 23704 21678
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23768 21146 23796 21490
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23860 19854 23888 21286
rect 24044 21078 24072 23462
rect 24032 21072 24084 21078
rect 24032 21014 24084 21020
rect 24136 20890 24164 23666
rect 24228 23202 24256 27095
rect 24780 25514 24808 27520
rect 24688 25486 24808 25514
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24688 24177 24716 25486
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24780 24954 24808 25327
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 25516 24585 25544 27520
rect 25502 24576 25558 24585
rect 25502 24511 25558 24520
rect 24766 24440 24822 24449
rect 24766 24375 24768 24384
rect 24820 24375 24822 24384
rect 24768 24346 24820 24352
rect 24674 24168 24730 24177
rect 24674 24103 24730 24112
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24766 23896 24822 23905
rect 24766 23831 24768 23840
rect 24820 23831 24822 23840
rect 24768 23802 24820 23808
rect 26160 23497 26188 27520
rect 26896 24449 26924 27520
rect 26882 24440 26938 24449
rect 26882 24375 26938 24384
rect 27540 23905 27568 27520
rect 27526 23896 27582 23905
rect 27526 23831 27582 23840
rect 24674 23488 24730 23497
rect 24674 23423 24730 23432
rect 26146 23488 26202 23497
rect 26146 23423 26202 23432
rect 24688 23322 24716 23423
rect 24676 23316 24728 23322
rect 24676 23258 24728 23264
rect 24228 23174 24716 23202
rect 24228 23089 24256 23174
rect 24214 23080 24270 23089
rect 24214 23015 24270 23024
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 24228 22642 24256 22918
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24228 21486 24256 21830
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24216 21480 24268 21486
rect 24216 21422 24268 21428
rect 24214 21040 24270 21049
rect 24688 21010 24716 23174
rect 24768 23180 24820 23186
rect 24768 23122 24820 23128
rect 24780 22438 24808 23122
rect 25410 23080 25466 23089
rect 25410 23015 25466 23024
rect 25424 22778 25452 23015
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24780 21944 24808 22374
rect 24780 21916 24900 21944
rect 24766 21856 24822 21865
rect 24766 21791 24822 21800
rect 24214 20975 24270 20984
rect 24676 21004 24728 21010
rect 24228 20942 24256 20975
rect 24676 20946 24728 20952
rect 23952 20862 24164 20890
rect 24216 20936 24268 20942
rect 24780 20890 24808 21791
rect 24216 20878 24268 20884
rect 24688 20862 24808 20890
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23676 19502 23796 19530
rect 23662 19408 23718 19417
rect 23662 19343 23718 19352
rect 23676 18970 23704 19343
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23676 18222 23704 18906
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23572 18148 23624 18154
rect 23572 18090 23624 18096
rect 23664 18080 23716 18086
rect 23400 18006 23520 18034
rect 23664 18022 23716 18028
rect 23296 17808 23348 17814
rect 23296 17750 23348 17756
rect 23296 17672 23348 17678
rect 23202 17640 23258 17649
rect 23296 17614 23348 17620
rect 23202 17575 23204 17584
rect 23256 17575 23258 17584
rect 23204 17546 23256 17552
rect 23308 17338 23336 17614
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23202 17096 23258 17105
rect 23308 17082 23336 17274
rect 23258 17054 23336 17082
rect 23202 17031 23258 17040
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 23032 16454 23060 16934
rect 23216 16726 23244 17031
rect 23204 16720 23256 16726
rect 23204 16662 23256 16668
rect 23492 16658 23520 18006
rect 23676 17882 23704 18022
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23584 16794 23612 17682
rect 23664 17264 23716 17270
rect 23768 17252 23796 19502
rect 23860 19242 23888 19790
rect 23952 19310 23980 20862
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24136 20398 24164 20742
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 24136 20058 24164 20198
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24030 19408 24086 19417
rect 24030 19343 24086 19352
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 23848 19236 23900 19242
rect 23848 19178 23900 19184
rect 23860 18766 23888 19178
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23952 18873 23980 19110
rect 23938 18864 23994 18873
rect 23938 18799 23994 18808
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23860 18426 23888 18702
rect 23848 18420 23900 18426
rect 23848 18362 23900 18368
rect 23848 18148 23900 18154
rect 23848 18090 23900 18096
rect 23716 17224 23796 17252
rect 23664 17206 23716 17212
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23676 16590 23704 16730
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 23032 15706 23060 16390
rect 23676 15910 23704 16526
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23570 15192 23626 15201
rect 23570 15127 23626 15136
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23124 14074 23152 14758
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23308 13802 23336 14418
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 23110 13696 23166 13705
rect 23110 13631 23166 13640
rect 22926 13560 22982 13569
rect 23124 13530 23152 13631
rect 22926 13495 22982 13504
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23032 12986 23060 13466
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23124 12850 23152 13466
rect 23308 13326 23336 13738
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23112 12844 23164 12850
rect 23112 12786 23164 12792
rect 23308 12646 23336 13262
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23204 12640 23256 12646
rect 23204 12582 23256 12588
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 23216 12481 23244 12582
rect 23202 12472 23258 12481
rect 23202 12407 23258 12416
rect 23492 12374 23520 12854
rect 23584 12594 23612 15127
rect 23676 12753 23704 15846
rect 23860 15201 23888 18090
rect 24044 16674 24072 19343
rect 24136 19310 24164 19994
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24228 19242 24256 20742
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20369 24716 20862
rect 24766 20768 24822 20777
rect 24766 20703 24822 20712
rect 24674 20360 24730 20369
rect 24674 20295 24730 20304
rect 24780 19961 24808 20703
rect 24872 20330 24900 21916
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25516 20942 25544 21286
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24860 20324 24912 20330
rect 24860 20266 24912 20272
rect 24964 20262 24992 20742
rect 25516 20602 25544 20878
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 24766 19952 24822 19961
rect 24766 19887 24822 19896
rect 24964 19802 24992 20198
rect 25056 19990 25084 20402
rect 25044 19984 25096 19990
rect 25044 19926 25096 19932
rect 24780 19774 24992 19802
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24216 19236 24268 19242
rect 24216 19178 24268 19184
rect 24124 19168 24176 19174
rect 24124 19110 24176 19116
rect 24136 16794 24164 19110
rect 24596 18902 24624 19314
rect 24674 19000 24730 19009
rect 24674 18935 24730 18944
rect 24216 18896 24268 18902
rect 24216 18838 24268 18844
rect 24584 18896 24636 18902
rect 24584 18838 24636 18844
rect 24228 17882 24256 18838
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24044 16646 24164 16674
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 24044 16250 24072 16526
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23846 15192 23902 15201
rect 23846 15127 23902 15136
rect 24136 14362 24164 16646
rect 24216 16652 24268 16658
rect 24216 16594 24268 16600
rect 24228 16250 24256 16594
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 24584 16040 24636 16046
rect 24582 16008 24584 16017
rect 24636 16008 24638 16017
rect 24582 15943 24638 15952
rect 24584 15564 24636 15570
rect 24688 15552 24716 18935
rect 24780 18408 24808 19774
rect 25056 19514 25084 19926
rect 25320 19712 25372 19718
rect 25320 19654 25372 19660
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 25332 19378 25360 19654
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25504 19304 25556 19310
rect 25504 19246 25556 19252
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25240 18426 25268 18566
rect 25228 18420 25280 18426
rect 24780 18380 24900 18408
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24780 17134 24808 18226
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24780 16794 24808 17070
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24766 16008 24822 16017
rect 24766 15943 24822 15952
rect 24780 15910 24808 15943
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24872 15722 24900 18380
rect 25228 18362 25280 18368
rect 25226 18320 25282 18329
rect 25226 18255 25282 18264
rect 25240 18222 25268 18255
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25412 18080 25464 18086
rect 25412 18022 25464 18028
rect 25424 17785 25452 18022
rect 25516 17921 25544 19246
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25700 18465 25728 19110
rect 25686 18456 25742 18465
rect 25686 18391 25742 18400
rect 25502 17912 25558 17921
rect 25502 17847 25558 17856
rect 25410 17776 25466 17785
rect 25410 17711 25466 17720
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24964 17241 24992 17478
rect 25608 17338 25636 17682
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 24950 17232 25006 17241
rect 24950 17167 25006 17176
rect 25228 16788 25280 16794
rect 25228 16730 25280 16736
rect 25240 16697 25268 16730
rect 25042 16688 25098 16697
rect 25042 16623 25044 16632
rect 25096 16623 25098 16632
rect 25226 16688 25282 16697
rect 25226 16623 25282 16632
rect 25044 16594 25096 16600
rect 25056 16250 25084 16594
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 24872 15694 24992 15722
rect 24688 15524 24900 15552
rect 24584 15506 24636 15512
rect 24596 15473 24624 15506
rect 24582 15464 24638 15473
rect 24766 15464 24822 15473
rect 24638 15422 24716 15450
rect 24582 15399 24638 15408
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15162 24716 15422
rect 24766 15399 24768 15408
rect 24820 15399 24822 15408
rect 24768 15370 24820 15376
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24582 15056 24638 15065
rect 24582 14991 24638 15000
rect 24596 14958 24624 14991
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24766 14920 24822 14929
rect 24766 14855 24822 14864
rect 24780 14822 24808 14855
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24872 14618 24900 15524
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24136 14334 24256 14362
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24136 14006 24164 14214
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24124 13728 24176 13734
rect 24124 13670 24176 13676
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23756 12776 23808 12782
rect 23662 12744 23718 12753
rect 23756 12718 23808 12724
rect 23662 12679 23718 12688
rect 23584 12566 23704 12594
rect 23480 12368 23532 12374
rect 23480 12310 23532 12316
rect 23570 12336 23626 12345
rect 23570 12271 23572 12280
rect 23624 12271 23626 12280
rect 23572 12242 23624 12248
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22744 11552 22796 11558
rect 22848 11529 22876 12038
rect 23676 11898 23704 12566
rect 23768 12442 23796 12718
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23480 11552 23532 11558
rect 22744 11494 22796 11500
rect 22834 11520 22890 11529
rect 22756 10266 22784 11494
rect 23480 11494 23532 11500
rect 22834 11455 22890 11464
rect 22848 11218 22876 11455
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22848 10810 22876 11154
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 23492 10282 23520 11494
rect 23860 11098 23888 13466
rect 24044 13258 24072 13670
rect 24136 13530 24164 13670
rect 24228 13530 24256 14334
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24766 13832 24822 13841
rect 24766 13767 24822 13776
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24582 13424 24638 13433
rect 24582 13359 24584 13368
rect 24636 13359 24638 13368
rect 24584 13330 24636 13336
rect 24596 13274 24624 13330
rect 24032 13252 24084 13258
rect 24596 13246 24716 13274
rect 24032 13194 24084 13200
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12986 24716 13246
rect 24780 13161 24808 13767
rect 24766 13152 24822 13161
rect 24766 13087 24822 13096
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24032 12640 24084 12646
rect 24768 12640 24820 12646
rect 24032 12582 24084 12588
rect 24766 12608 24768 12617
rect 24820 12608 24822 12617
rect 23572 11076 23624 11082
rect 23860 11070 23980 11098
rect 23572 11018 23624 11024
rect 23400 10266 23520 10282
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23388 10260 23520 10266
rect 23440 10254 23520 10260
rect 23388 10202 23440 10208
rect 23032 9110 23060 10202
rect 23480 10192 23532 10198
rect 23480 10134 23532 10140
rect 23492 9450 23520 10134
rect 23584 9897 23612 11018
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23860 10538 23888 10950
rect 23848 10532 23900 10538
rect 23848 10474 23900 10480
rect 23664 10464 23716 10470
rect 23860 10441 23888 10474
rect 23664 10406 23716 10412
rect 23846 10432 23902 10441
rect 23676 9926 23704 10406
rect 23846 10367 23902 10376
rect 23664 9920 23716 9926
rect 23570 9888 23626 9897
rect 23664 9862 23716 9868
rect 23570 9823 23626 9832
rect 23676 9738 23704 9862
rect 23584 9710 23704 9738
rect 23480 9444 23532 9450
rect 23480 9386 23532 9392
rect 23584 9382 23612 9710
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 23020 9104 23072 9110
rect 23020 9046 23072 9052
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22940 8634 22968 8910
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23400 8430 23428 9318
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 22928 7948 22980 7954
rect 22928 7890 22980 7896
rect 22560 7812 22612 7818
rect 22664 7806 22784 7834
rect 22560 7754 22612 7760
rect 22572 7342 22600 7754
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 7546 22692 7686
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22664 7410 22692 7482
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22572 6866 22600 7278
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 22572 6458 22600 6802
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22480 5370 22508 5714
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22112 5222 22232 5250
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 22006 4720 22062 4729
rect 22006 4655 22062 4664
rect 22112 3738 22140 5102
rect 22204 4078 22232 5222
rect 22756 5137 22784 7806
rect 22940 7002 22968 7890
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 22940 6322 22968 6938
rect 23020 6860 23072 6866
rect 23020 6802 23072 6808
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 22940 5914 22968 6258
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 23032 5556 23060 6802
rect 23676 6322 23704 9590
rect 23846 9480 23902 9489
rect 23846 9415 23902 9424
rect 23754 9344 23810 9353
rect 23754 9279 23810 9288
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23400 6186 23704 6202
rect 23388 6180 23704 6186
rect 23440 6174 23704 6180
rect 23388 6122 23440 6128
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 23112 5568 23164 5574
rect 23032 5528 23112 5556
rect 23112 5510 23164 5516
rect 23296 5568 23348 5574
rect 23296 5510 23348 5516
rect 23124 5370 23152 5510
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23308 5166 23336 5510
rect 23296 5160 23348 5166
rect 22742 5128 22798 5137
rect 23296 5102 23348 5108
rect 22742 5063 22798 5072
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22388 3777 22416 3878
rect 22374 3768 22430 3777
rect 22100 3732 22152 3738
rect 22480 3738 22508 4966
rect 23124 4486 23152 4966
rect 23296 4820 23348 4826
rect 23296 4762 23348 4768
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 23124 4214 23152 4422
rect 23112 4208 23164 4214
rect 22558 4176 22614 4185
rect 23112 4150 23164 4156
rect 22558 4111 22614 4120
rect 22374 3703 22430 3712
rect 22468 3732 22520 3738
rect 22100 3674 22152 3680
rect 22468 3674 22520 3680
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21744 3194 21772 3470
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 22572 2990 22600 4111
rect 23216 3670 23244 4626
rect 23308 3738 23336 4762
rect 23400 4026 23428 5578
rect 23492 4826 23520 5646
rect 23584 5234 23612 6054
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 23400 3998 23520 4026
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 22744 3664 22796 3670
rect 22742 3632 22744 3641
rect 23204 3664 23256 3670
rect 22796 3632 22798 3641
rect 23204 3606 23256 3612
rect 22742 3567 22798 3576
rect 23296 3460 23348 3466
rect 23296 3402 23348 3408
rect 23308 3194 23336 3402
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 22742 3088 22798 3097
rect 22742 3023 22798 3032
rect 22560 2984 22612 2990
rect 22480 2932 22560 2938
rect 22480 2926 22612 2932
rect 22480 2910 22600 2926
rect 22480 2650 22508 2910
rect 22652 2848 22704 2854
rect 22650 2816 22652 2825
rect 22704 2816 22706 2825
rect 22650 2751 22706 2760
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 22098 2408 22154 2417
rect 22098 2343 22154 2352
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 20718 2000 20774 2009
rect 20718 1935 20774 1944
rect 20444 604 20496 610
rect 20444 546 20496 552
rect 20732 480 20760 1935
rect 21928 1465 21956 2246
rect 21914 1456 21970 1465
rect 21914 1391 21970 1400
rect 21364 604 21416 610
rect 21364 546 21416 552
rect 21376 480 21404 546
rect 22112 480 22140 2343
rect 22756 480 22784 3023
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22848 2145 22876 2450
rect 22834 2136 22890 2145
rect 22834 2071 22890 2080
rect 23492 480 23520 3998
rect 23676 3913 23704 6174
rect 23662 3904 23718 3913
rect 23662 3839 23718 3848
rect 23768 3641 23796 9279
rect 23860 7313 23888 9415
rect 23952 9178 23980 11070
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 24044 8906 24072 12582
rect 24766 12543 24822 12552
rect 24964 12442 24992 15694
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25792 14074 25820 14418
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25412 14000 25464 14006
rect 25042 13968 25098 13977
rect 25412 13942 25464 13948
rect 25042 13903 25044 13912
rect 25096 13903 25098 13912
rect 25044 13874 25096 13880
rect 25424 13705 25452 13942
rect 25410 13696 25466 13705
rect 25410 13631 25466 13640
rect 25410 12472 25466 12481
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24952 12436 25004 12442
rect 25410 12407 25466 12416
rect 24952 12378 25004 12384
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 24136 11626 24164 12038
rect 24124 11620 24176 11626
rect 24124 11562 24176 11568
rect 24136 10198 24164 11562
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24124 9648 24176 9654
rect 24228 9636 24256 12378
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12242
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24780 11937 24808 12038
rect 24766 11928 24822 11937
rect 24676 11892 24728 11898
rect 24766 11863 24822 11872
rect 24676 11834 24728 11840
rect 25226 11384 25282 11393
rect 25226 11319 25228 11328
rect 25280 11319 25282 11328
rect 25228 11290 25280 11296
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 25056 10198 25084 10406
rect 25240 10266 25268 11290
rect 25424 11150 25452 12407
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25412 11144 25464 11150
rect 25412 11086 25464 11092
rect 25424 10810 25452 11086
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 25608 10470 25636 11154
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25608 10305 25636 10406
rect 25594 10296 25650 10305
rect 25228 10260 25280 10266
rect 25594 10231 25650 10240
rect 25228 10202 25280 10208
rect 25044 10192 25096 10198
rect 25044 10134 25096 10140
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24176 9608 24256 9636
rect 24872 9602 24900 9862
rect 24124 9590 24176 9596
rect 24780 9574 24900 9602
rect 24780 9518 24808 9574
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24780 9110 24808 9454
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24768 9104 24820 9110
rect 24674 9072 24730 9081
rect 24584 9036 24636 9042
rect 24768 9046 24820 9052
rect 24674 9007 24676 9016
rect 24584 8978 24636 8984
rect 24728 9007 24730 9016
rect 24676 8978 24728 8984
rect 24596 8922 24624 8978
rect 24766 8936 24822 8945
rect 24032 8900 24084 8906
rect 24596 8894 24716 8922
rect 24032 8842 24084 8848
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24688 8537 24716 8894
rect 24766 8871 24822 8880
rect 24674 8528 24730 8537
rect 24674 8463 24730 8472
rect 24688 8430 24716 8463
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24032 8356 24084 8362
rect 24032 8298 24084 8304
rect 24400 8356 24452 8362
rect 24400 8298 24452 8304
rect 23846 7304 23902 7313
rect 23846 7239 23902 7248
rect 24044 6458 24072 8298
rect 24412 8022 24440 8298
rect 24400 8016 24452 8022
rect 24780 7993 24808 8871
rect 24872 8362 24900 9318
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24964 8294 24992 8842
rect 24952 8288 25004 8294
rect 24952 8230 25004 8236
rect 24964 8090 24992 8230
rect 24952 8084 25004 8090
rect 24952 8026 25004 8032
rect 24400 7958 24452 7964
rect 24766 7984 24822 7993
rect 24766 7919 24822 7928
rect 24122 7848 24178 7857
rect 24122 7783 24178 7792
rect 24136 7410 24164 7783
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24320 7002 24348 7346
rect 24308 6996 24360 7002
rect 24308 6938 24360 6944
rect 25226 6896 25282 6905
rect 25226 6831 25228 6840
rect 25280 6831 25282 6840
rect 25228 6802 25280 6808
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 25240 6458 25268 6802
rect 25412 6656 25464 6662
rect 25412 6598 25464 6604
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 23848 4752 23900 4758
rect 23846 4720 23848 4729
rect 23900 4720 23902 4729
rect 23846 4655 23902 4664
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23754 3632 23810 3641
rect 23754 3567 23810 3576
rect 23860 3534 23888 3946
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23848 3528 23900 3534
rect 23952 3505 23980 6258
rect 24674 6080 24730 6089
rect 24674 6015 24730 6024
rect 24032 5636 24084 5642
rect 24032 5578 24084 5584
rect 24044 5098 24072 5578
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24032 5092 24084 5098
rect 24032 5034 24084 5040
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24030 4040 24086 4049
rect 24030 3975 24086 3984
rect 23848 3470 23900 3476
rect 23938 3496 23994 3505
rect 23768 3369 23796 3470
rect 23754 3360 23810 3369
rect 23754 3295 23810 3304
rect 23570 3224 23626 3233
rect 23768 3194 23796 3295
rect 23570 3159 23626 3168
rect 23756 3188 23808 3194
rect 23584 921 23612 3159
rect 23756 3130 23808 3136
rect 23860 2650 23888 3470
rect 23938 3431 23994 3440
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23952 2514 23980 3431
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 24044 1601 24072 3975
rect 24122 3768 24178 3777
rect 24122 3703 24178 3712
rect 24030 1592 24086 1601
rect 24030 1527 24086 1536
rect 23570 912 23626 921
rect 23570 847 23626 856
rect 24136 480 24164 3703
rect 24688 3346 24716 6015
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24872 5370 24900 5714
rect 25056 5574 25084 6258
rect 25136 6180 25188 6186
rect 25136 6122 25188 6128
rect 25148 5914 25176 6122
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24780 3466 24808 4422
rect 24872 3738 24900 5306
rect 24952 4752 25004 4758
rect 24952 4694 25004 4700
rect 24964 4457 24992 4694
rect 24950 4448 25006 4457
rect 24950 4383 25006 4392
rect 24964 3738 24992 4383
rect 25056 4282 25084 5510
rect 25044 4276 25096 4282
rect 25044 4218 25096 4224
rect 25424 4185 25452 6598
rect 25410 4176 25466 4185
rect 25410 4111 25466 4120
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 24872 3346 24900 3470
rect 24688 3318 24900 3346
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24872 3194 24900 3318
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24766 2952 24822 2961
rect 24766 2887 24822 2896
rect 24780 2854 24808 2887
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 24872 2666 24900 3130
rect 24964 3058 24992 3674
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25516 3194 25544 3470
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 24952 3052 25004 3058
rect 24952 2994 25004 3000
rect 27526 2952 27582 2961
rect 27526 2887 27582 2896
rect 25502 2816 25558 2825
rect 25502 2751 25558 2760
rect 24780 2638 24900 2666
rect 24676 2372 24728 2378
rect 24676 2314 24728 2320
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24582 1320 24638 1329
rect 24582 1255 24638 1264
rect 294 0 350 480
rect 938 0 994 480
rect 1582 0 1638 480
rect 2318 0 2374 480
rect 2962 0 3018 480
rect 3698 0 3754 480
rect 4342 0 4398 480
rect 4986 0 5042 480
rect 5722 0 5778 480
rect 6366 0 6422 480
rect 7102 0 7158 480
rect 7746 0 7802 480
rect 8390 0 8446 480
rect 9126 0 9182 480
rect 9770 0 9826 480
rect 10506 0 10562 480
rect 11150 0 11206 480
rect 11886 0 11942 480
rect 12530 0 12586 480
rect 13174 0 13230 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15290 0 15346 480
rect 15934 0 15990 480
rect 16578 0 16634 480
rect 17314 0 17370 480
rect 17958 0 18014 480
rect 18694 0 18750 480
rect 19338 0 19394 480
rect 20074 0 20130 480
rect 20718 0 20774 480
rect 21362 0 21418 480
rect 22098 0 22154 480
rect 22742 0 22798 480
rect 23478 0 23534 480
rect 24122 0 24178 480
rect 24596 377 24624 1255
rect 24688 1170 24716 2314
rect 24780 1329 24808 2638
rect 24766 1320 24822 1329
rect 24766 1255 24822 1264
rect 24688 1142 24808 1170
rect 24780 480 24808 1142
rect 25516 480 25544 2751
rect 26148 2372 26200 2378
rect 26148 2314 26200 2320
rect 26160 480 26188 2314
rect 26790 1456 26846 1465
rect 26846 1414 26924 1442
rect 26790 1391 26846 1400
rect 26896 480 26924 1414
rect 27540 480 27568 2887
rect 24582 368 24638 377
rect 24582 303 24638 312
rect 24766 0 24822 480
rect 25502 0 25558 480
rect 26146 0 26202 480
rect 26882 0 26938 480
rect 27526 0 27582 480
<< via2 >>
rect 23202 27648 23258 27704
rect 1582 24656 1638 24712
rect 1490 22616 1546 22672
rect 1582 20868 1638 20904
rect 1582 20848 1584 20868
rect 1584 20848 1636 20868
rect 1636 20848 1638 20868
rect 1582 20304 1638 20360
rect 938 3440 994 3496
rect 294 1672 350 1728
rect 1674 13912 1730 13968
rect 1490 9696 1546 9752
rect 2962 24792 3018 24848
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4986 24112 5042 24168
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 4342 23704 4398 23760
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 3698 22480 3754 22536
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6366 23840 6422 23896
rect 5998 21664 6054 21720
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 7102 19216 7158 19272
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 9126 20712 9182 20768
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10690 23160 10746 23216
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 9954 22208 10010 22264
rect 9770 20984 9826 21040
rect 11058 21684 11114 21720
rect 11058 21664 11060 21684
rect 11060 21664 11112 21684
rect 11112 21664 11114 21684
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10322 20460 10378 20496
rect 10322 20440 10324 20460
rect 10324 20440 10376 20460
rect 10376 20440 10378 20460
rect 12346 24792 12402 24848
rect 11886 24384 11942 24440
rect 11518 24112 11574 24168
rect 11426 23840 11482 23896
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9954 19760 10010 19816
rect 10782 19216 10838 19272
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 7746 17720 7802 17776
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 9586 16088 9642 16144
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 2318 13232 2374 13288
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 4986 11600 5042 11656
rect 4342 10104 4398 10160
rect 2870 9696 2926 9752
rect 2778 9560 2834 9616
rect 2870 9288 2926 9344
rect 2318 6296 2374 6352
rect 1950 3440 2006 3496
rect 3698 7928 3754 7984
rect 2962 5072 3018 5128
rect 2870 4664 2926 4720
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 9494 15136 9550 15192
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10874 17176 10930 17232
rect 10782 14592 10838 14648
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10874 10684 10876 10704
rect 10876 10684 10928 10704
rect 10928 10684 10930 10704
rect 10874 10648 10930 10684
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6918 7520 6974 7576
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 11242 17856 11298 17912
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10138 9560 10194 9616
rect 10966 9560 11022 9616
rect 9678 9324 9680 9344
rect 9680 9324 9732 9344
rect 9732 9324 9734 9344
rect 9678 9288 9734 9324
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 9126 8880 9182 8936
rect 8298 4664 8354 4720
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5722 2488 5778 2544
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7102 3984 7158 4040
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10782 4936 10838 4992
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 9770 4528 9826 4584
rect 10690 4120 10746 4176
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3188 10194 3224
rect 10138 3168 10140 3188
rect 10140 3168 10192 3188
rect 10192 3168 10194 3188
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11058 8472 11114 8528
rect 11058 3984 11114 4040
rect 10966 1400 11022 1456
rect 12990 24656 13046 24712
rect 13174 23704 13230 23760
rect 12530 23568 12586 23624
rect 12530 23160 12586 23216
rect 11702 20984 11758 21040
rect 12070 19896 12126 19952
rect 11702 18128 11758 18184
rect 11610 14456 11666 14512
rect 11610 14320 11666 14376
rect 11426 3068 11428 3088
rect 11428 3068 11480 3088
rect 11480 3068 11482 3088
rect 11426 3032 11482 3068
rect 11610 2760 11666 2816
rect 11886 5616 11942 5672
rect 12438 19216 12494 19272
rect 12714 20168 12770 20224
rect 12346 12552 12402 12608
rect 12070 11736 12126 11792
rect 12346 11600 12402 11656
rect 12530 11092 12532 11112
rect 12532 11092 12584 11112
rect 12584 11092 12586 11112
rect 12530 11056 12586 11092
rect 12438 10648 12494 10704
rect 12254 8880 12310 8936
rect 12254 7656 12310 7712
rect 12806 19216 12862 19272
rect 12714 9016 12770 9072
rect 12530 7928 12586 7984
rect 12438 7520 12494 7576
rect 12254 6568 12310 6624
rect 11702 2488 11758 2544
rect 11610 1536 11666 1592
rect 12438 3576 12494 3632
rect 12714 3732 12770 3768
rect 12714 3712 12716 3732
rect 12716 3712 12768 3732
rect 12768 3712 12770 3732
rect 12622 1672 12678 1728
rect 13174 20032 13230 20088
rect 13174 19116 13176 19136
rect 13176 19116 13228 19136
rect 13228 19116 13230 19136
rect 13174 19080 13230 19116
rect 13542 24384 13598 24440
rect 13634 20984 13690 21040
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14554 24792 14610 24848
rect 14462 24656 14518 24712
rect 14094 22072 14150 22128
rect 14094 20848 14150 20904
rect 14094 20712 14150 20768
rect 14186 20204 14188 20224
rect 14188 20204 14240 20224
rect 14240 20204 14242 20224
rect 14186 20168 14242 20204
rect 14094 18672 14150 18728
rect 13358 18264 13414 18320
rect 13358 16496 13414 16552
rect 13266 14320 13322 14376
rect 13266 13912 13322 13968
rect 13542 15952 13598 16008
rect 13726 15000 13782 15056
rect 13450 14728 13506 14784
rect 13082 13232 13138 13288
rect 13082 12824 13138 12880
rect 12898 6296 12954 6352
rect 13358 12688 13414 12744
rect 14002 17856 14058 17912
rect 14278 17756 14280 17776
rect 14280 17756 14332 17776
rect 14332 17756 14334 17776
rect 14278 17720 14334 17756
rect 14278 16940 14280 16960
rect 14280 16940 14332 16960
rect 14332 16940 14334 16960
rect 14278 16904 14334 16940
rect 14186 15136 14242 15192
rect 14094 14456 14150 14512
rect 14002 13776 14058 13832
rect 13910 12552 13966 12608
rect 13634 10512 13690 10568
rect 13542 10104 13598 10160
rect 13634 9968 13690 10024
rect 13634 8880 13690 8936
rect 13910 9560 13966 9616
rect 13910 9324 13912 9344
rect 13912 9324 13964 9344
rect 13964 9324 13966 9344
rect 13910 9288 13966 9324
rect 13542 6704 13598 6760
rect 13450 5752 13506 5808
rect 14278 14340 14334 14376
rect 14278 14320 14280 14340
rect 14280 14320 14332 14340
rect 14332 14320 14334 14340
rect 14186 13388 14242 13424
rect 14186 13368 14188 13388
rect 14188 13368 14240 13388
rect 14240 13368 14242 13388
rect 14278 13268 14280 13288
rect 14280 13268 14332 13288
rect 14332 13268 14334 13288
rect 14278 13232 14334 13268
rect 14554 23840 14610 23896
rect 14462 23060 14464 23080
rect 14464 23060 14516 23080
rect 14516 23060 14518 23080
rect 14462 23024 14518 23060
rect 15934 24792 15990 24848
rect 15382 24520 15438 24576
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15474 22888 15530 22944
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15382 22380 15384 22400
rect 15384 22380 15436 22400
rect 15436 22380 15438 22400
rect 15382 22344 15438 22380
rect 15290 21972 15292 21992
rect 15292 21972 15344 21992
rect 15344 21972 15346 21992
rect 15290 21936 15346 21972
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15382 18264 15438 18320
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15474 16904 15530 16960
rect 15658 24012 15660 24032
rect 15660 24012 15712 24032
rect 15712 24012 15714 24032
rect 15658 23976 15714 24012
rect 16118 23704 16174 23760
rect 15658 20440 15714 20496
rect 16026 21800 16082 21856
rect 15750 20032 15806 20088
rect 16026 20032 16082 20088
rect 15934 19760 15990 19816
rect 15658 17448 15714 17504
rect 14738 16088 14794 16144
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15566 16496 15622 16552
rect 15198 15680 15254 15736
rect 15106 15428 15162 15464
rect 15106 15408 15108 15428
rect 15108 15408 15160 15428
rect 15160 15408 15162 15428
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15750 15156 15806 15192
rect 15750 15136 15752 15156
rect 15752 15136 15804 15156
rect 15804 15136 15806 15156
rect 15750 14728 15806 14784
rect 15474 14592 15530 14648
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15566 13812 15568 13832
rect 15568 13812 15620 13832
rect 15620 13812 15622 13832
rect 15566 13776 15622 13812
rect 16026 17312 16082 17368
rect 16302 23568 16358 23624
rect 17038 23860 17094 23896
rect 17038 23840 17040 23860
rect 17040 23840 17092 23860
rect 17092 23840 17094 23860
rect 17038 23432 17094 23488
rect 16486 22616 16542 22672
rect 16302 18536 16358 18592
rect 16578 20476 16580 20496
rect 16580 20476 16632 20496
rect 16632 20476 16634 20496
rect 16578 20440 16634 20476
rect 17774 23704 17830 23760
rect 18142 23568 18198 23624
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 17406 22480 17462 22536
rect 16210 15544 16266 15600
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15474 11328 15530 11384
rect 14554 10412 14556 10432
rect 14556 10412 14608 10432
rect 14608 10412 14610 10432
rect 14554 10376 14610 10412
rect 14462 10104 14518 10160
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14186 6604 14188 6624
rect 14188 6604 14240 6624
rect 14240 6604 14242 6624
rect 14186 6568 14242 6604
rect 14094 5208 14150 5264
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15474 10512 15530 10568
rect 16854 17720 16910 17776
rect 16762 16088 16818 16144
rect 17406 17076 17408 17096
rect 17408 17076 17460 17096
rect 17460 17076 17462 17096
rect 17406 17040 17462 17076
rect 17222 16360 17278 16416
rect 16210 12280 16266 12336
rect 15566 9832 15622 9888
rect 15566 7928 15622 7984
rect 15290 6704 15346 6760
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14462 6296 14518 6352
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14646 4800 14702 4856
rect 14646 4528 14702 4584
rect 13634 3460 13690 3496
rect 13634 3440 13636 3460
rect 13636 3440 13688 3460
rect 13688 3440 13690 3460
rect 13634 2896 13690 2952
rect 13082 2644 13138 2680
rect 13082 2624 13084 2644
rect 13084 2624 13136 2644
rect 13136 2624 13138 2644
rect 14554 2760 14610 2816
rect 13358 1944 13414 2000
rect 14462 2372 14518 2408
rect 14462 2352 14464 2372
rect 14464 2352 14516 2372
rect 14516 2352 14518 2372
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15382 4120 15438 4176
rect 14738 3984 14794 4040
rect 15842 10512 15898 10568
rect 17038 13232 17094 13288
rect 17590 11736 17646 11792
rect 17498 10376 17554 10432
rect 16762 10124 16818 10160
rect 16762 10104 16764 10124
rect 16764 10104 16816 10124
rect 16816 10104 16818 10124
rect 16486 6604 16488 6624
rect 16488 6604 16540 6624
rect 16540 6604 16542 6624
rect 16486 6568 16542 6604
rect 16210 6296 16266 6352
rect 16026 4664 16082 4720
rect 14738 3168 14794 3224
rect 15382 3304 15438 3360
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15474 3168 15530 3224
rect 15750 2760 15806 2816
rect 14830 2524 14832 2544
rect 14832 2524 14884 2544
rect 14884 2524 14886 2544
rect 14830 2488 14886 2524
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17038 8916 17040 8936
rect 17040 8916 17092 8936
rect 17092 8916 17094 8936
rect 17038 8880 17094 8916
rect 18510 21936 18566 21992
rect 18694 23432 18750 23488
rect 19154 22480 19210 22536
rect 20166 24792 20222 24848
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19430 23840 19486 23896
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 18786 20748 18788 20768
rect 18788 20748 18840 20768
rect 18840 20748 18842 20768
rect 18786 20712 18842 20748
rect 18694 19372 18750 19408
rect 18694 19352 18696 19372
rect 18696 19352 18748 19372
rect 18748 19352 18750 19372
rect 17958 17584 18014 17640
rect 18234 16632 18290 16688
rect 18234 15544 18290 15600
rect 18142 12316 18144 12336
rect 18144 12316 18196 12336
rect 18196 12316 18198 12336
rect 18142 12280 18198 12316
rect 18234 11348 18290 11384
rect 18234 11328 18236 11348
rect 18236 11328 18288 11348
rect 18288 11328 18290 11348
rect 18050 11056 18106 11112
rect 17774 10784 17830 10840
rect 17314 7248 17370 7304
rect 16946 6568 17002 6624
rect 16854 5208 16910 5264
rect 16762 4800 16818 4856
rect 16026 4120 16082 4176
rect 16118 3596 16174 3632
rect 16118 3576 16120 3596
rect 16120 3576 16172 3596
rect 16172 3576 16174 3596
rect 15934 3032 15990 3088
rect 15290 1400 15346 1456
rect 15842 1400 15898 1456
rect 16118 2644 16174 2680
rect 16118 2624 16120 2644
rect 16120 2624 16172 2644
rect 16172 2624 16174 2644
rect 16578 4020 16580 4040
rect 16580 4020 16632 4040
rect 16632 4020 16634 4040
rect 16578 3984 16634 4020
rect 16578 3712 16634 3768
rect 17958 9968 18014 10024
rect 17774 9288 17830 9344
rect 18234 8608 18290 8664
rect 18418 10648 18474 10704
rect 18602 19080 18658 19136
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 18602 18420 18658 18456
rect 18602 18400 18604 18420
rect 18604 18400 18656 18420
rect 18656 18400 18658 18420
rect 19062 17176 19118 17232
rect 19430 18672 19486 18728
rect 19338 16904 19394 16960
rect 19062 14864 19118 14920
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19798 18828 19854 18864
rect 19798 18808 19800 18828
rect 19800 18808 19852 18828
rect 19852 18808 19854 18828
rect 21362 24792 21418 24848
rect 20626 23976 20682 24032
rect 20534 23704 20590 23760
rect 20074 22344 20130 22400
rect 20902 23568 20958 23624
rect 20718 23044 20774 23080
rect 20718 23024 20720 23044
rect 20720 23024 20772 23044
rect 20772 23024 20774 23044
rect 20994 23024 21050 23080
rect 20442 19352 20498 19408
rect 20626 19352 20682 19408
rect 19982 18264 20038 18320
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19798 17584 19854 17640
rect 20074 17876 20130 17912
rect 20074 17856 20076 17876
rect 20076 17856 20128 17876
rect 20128 17856 20130 17876
rect 20166 17720 20222 17776
rect 19982 17312 20038 17368
rect 20350 18808 20406 18864
rect 20350 17584 20406 17640
rect 20258 17176 20314 17232
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20534 16088 20590 16144
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19154 14048 19210 14104
rect 18878 12844 18934 12880
rect 18878 12824 18880 12844
rect 18880 12824 18932 12844
rect 18932 12824 18934 12844
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 18786 10512 18842 10568
rect 17590 5752 17646 5808
rect 17774 6568 17830 6624
rect 17038 4256 17094 4312
rect 17958 2896 18014 2952
rect 16946 2080 17002 2136
rect 17314 1536 17370 1592
rect 18694 9696 18750 9752
rect 18510 9560 18566 9616
rect 18418 8356 18474 8392
rect 18418 8336 18420 8356
rect 18420 8336 18472 8356
rect 18472 8336 18474 8356
rect 18510 7948 18566 7984
rect 18510 7928 18512 7948
rect 18512 7928 18564 7948
rect 18564 7928 18566 7948
rect 18050 2524 18052 2544
rect 18052 2524 18104 2544
rect 18104 2524 18106 2544
rect 18050 2488 18106 2524
rect 18602 4528 18658 4584
rect 18878 6704 18934 6760
rect 18694 4392 18750 4448
rect 18694 4120 18750 4176
rect 20718 15544 20774 15600
rect 20442 15136 20498 15192
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19246 10648 19302 10704
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 20258 12280 20314 12336
rect 20074 11500 20076 11520
rect 20076 11500 20128 11520
rect 20128 11500 20130 11520
rect 20074 11464 20130 11500
rect 20074 10240 20130 10296
rect 19338 9016 19394 9072
rect 19154 6160 19210 6216
rect 19062 5788 19064 5808
rect 19064 5788 19116 5808
rect 19116 5788 19118 5808
rect 19062 5752 19118 5788
rect 18878 5244 18880 5264
rect 18880 5244 18932 5264
rect 18932 5244 18934 5264
rect 18878 5208 18934 5244
rect 18878 2624 18934 2680
rect 18786 2488 18842 2544
rect 19154 4020 19156 4040
rect 19156 4020 19208 4040
rect 19208 4020 19210 4040
rect 19154 3984 19210 4020
rect 19338 4256 19394 4312
rect 19154 3476 19156 3496
rect 19156 3476 19208 3496
rect 19208 3476 19210 3496
rect 19154 3440 19210 3476
rect 21270 24656 21326 24712
rect 21086 22888 21142 22944
rect 21270 18400 21326 18456
rect 20994 16360 21050 16416
rect 21270 15136 21326 15192
rect 21362 14884 21418 14920
rect 21362 14864 21364 14884
rect 21364 14864 21416 14884
rect 21416 14864 21418 14884
rect 21086 13776 21142 13832
rect 20718 13640 20774 13696
rect 20810 12688 20866 12744
rect 20442 10784 20498 10840
rect 20810 10532 20866 10568
rect 20810 10512 20812 10532
rect 20812 10512 20864 10532
rect 20864 10512 20866 10532
rect 20074 8608 20130 8664
rect 20074 8336 20130 8392
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19522 7792 19578 7848
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 20166 7792 20222 7848
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 20074 4800 20130 4856
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19522 3304 19578 3360
rect 19522 2896 19578 2952
rect 22650 24112 22706 24168
rect 22742 23296 22798 23352
rect 22558 21256 22614 21312
rect 21914 20712 21970 20768
rect 21822 19624 21878 19680
rect 21638 17448 21694 17504
rect 22098 18128 22154 18184
rect 21546 13368 21602 13424
rect 21086 9460 21088 9480
rect 21088 9460 21140 9480
rect 21140 9460 21142 9480
rect 21086 9424 21142 9460
rect 21178 9288 21234 9344
rect 20994 9016 21050 9072
rect 21178 9016 21234 9072
rect 21546 9696 21602 9752
rect 21270 7112 21326 7168
rect 21730 8508 21732 8528
rect 21732 8508 21784 8528
rect 21784 8508 21786 8528
rect 21730 8472 21786 8508
rect 21086 6296 21142 6352
rect 21362 6160 21418 6216
rect 20902 5752 20958 5808
rect 21086 5752 21142 5808
rect 20350 5208 20406 5264
rect 21270 5616 21326 5672
rect 20442 3168 20498 3224
rect 20258 3032 20314 3088
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20902 4664 20958 4720
rect 20902 4528 20958 4584
rect 21178 4392 21234 4448
rect 22006 12280 22062 12336
rect 22282 17176 22338 17232
rect 22190 14048 22246 14104
rect 22926 23160 22982 23216
rect 23294 26560 23350 26616
rect 23662 25880 23718 25936
rect 23754 24792 23810 24848
rect 23478 24656 23534 24712
rect 23662 24520 23718 24576
rect 23662 23568 23718 23624
rect 23294 22380 23296 22400
rect 23296 22380 23348 22400
rect 23348 22380 23350 22400
rect 23294 22344 23350 22380
rect 21914 11328 21970 11384
rect 21914 10376 21970 10432
rect 21546 6060 21548 6080
rect 21548 6060 21600 6080
rect 21600 6060 21602 6080
rect 21546 6024 21602 6060
rect 22098 7112 22154 7168
rect 22006 6840 22062 6896
rect 21638 5208 21694 5264
rect 21454 3168 21510 3224
rect 22190 6432 22246 6488
rect 22558 8336 22614 8392
rect 23202 18536 23258 18592
rect 23478 21800 23534 21856
rect 24214 27104 24270 27160
rect 23938 24248 23994 24304
rect 23846 23296 23902 23352
rect 23938 22480 23994 22536
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 25336 24822 25392
rect 25502 24520 25558 24576
rect 24766 24404 24822 24440
rect 24766 24384 24768 24404
rect 24768 24384 24820 24404
rect 24820 24384 24822 24404
rect 24674 24112 24730 24168
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 23860 24822 23896
rect 24766 23840 24768 23860
rect 24768 23840 24820 23860
rect 24820 23840 24822 23860
rect 26882 24384 26938 24440
rect 27526 23840 27582 23896
rect 24674 23432 24730 23488
rect 26146 23432 26202 23488
rect 24214 23024 24270 23080
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24214 20984 24270 21040
rect 25410 23024 25466 23080
rect 24766 21800 24822 21856
rect 23662 19352 23718 19408
rect 23202 17604 23258 17640
rect 23202 17584 23204 17604
rect 23204 17584 23256 17604
rect 23256 17584 23258 17604
rect 23202 17040 23258 17096
rect 24030 19352 24086 19408
rect 23938 18808 23994 18864
rect 23570 15136 23626 15192
rect 23110 13640 23166 13696
rect 22926 13504 22982 13560
rect 23202 12416 23258 12472
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 20712 24822 20768
rect 24674 20304 24730 20360
rect 24766 19896 24822 19952
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24674 18944 24730 19000
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 23846 15136 23902 15192
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24582 15988 24584 16008
rect 24584 15988 24636 16008
rect 24636 15988 24638 16008
rect 24582 15952 24638 15988
rect 24766 15952 24822 16008
rect 25226 18264 25282 18320
rect 25686 18400 25742 18456
rect 25502 17856 25558 17912
rect 25410 17720 25466 17776
rect 24950 17176 25006 17232
rect 25042 16652 25098 16688
rect 25042 16632 25044 16652
rect 25044 16632 25096 16652
rect 25096 16632 25098 16652
rect 25226 16632 25282 16688
rect 24582 15408 24638 15464
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24766 15428 24822 15464
rect 24766 15408 24768 15428
rect 24768 15408 24820 15428
rect 24820 15408 24822 15428
rect 24582 15000 24638 15056
rect 24766 14864 24822 14920
rect 23662 12688 23718 12744
rect 23570 12300 23626 12336
rect 23570 12280 23572 12300
rect 23572 12280 23624 12300
rect 23624 12280 23626 12300
rect 22834 11464 22890 11520
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 13776 24822 13832
rect 24582 13388 24638 13424
rect 24582 13368 24584 13388
rect 24584 13368 24636 13388
rect 24636 13368 24638 13388
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24766 13096 24822 13152
rect 24766 12588 24768 12608
rect 24768 12588 24820 12608
rect 24820 12588 24822 12608
rect 23846 10376 23902 10432
rect 23570 9832 23626 9888
rect 22006 4664 22062 4720
rect 23846 9424 23902 9480
rect 23754 9288 23810 9344
rect 22742 5072 22798 5128
rect 22374 3712 22430 3768
rect 22558 4120 22614 4176
rect 22742 3612 22744 3632
rect 22744 3612 22796 3632
rect 22796 3612 22798 3632
rect 22742 3576 22798 3612
rect 22742 3032 22798 3088
rect 22650 2796 22652 2816
rect 22652 2796 22704 2816
rect 22704 2796 22706 2816
rect 22650 2760 22706 2796
rect 22098 2352 22154 2408
rect 20718 1944 20774 2000
rect 21914 1400 21970 1456
rect 22834 2080 22890 2136
rect 23662 3848 23718 3904
rect 24766 12552 24822 12588
rect 25042 13932 25098 13968
rect 25042 13912 25044 13932
rect 25044 13912 25096 13932
rect 25096 13912 25098 13932
rect 25410 13640 25466 13696
rect 25410 12416 25466 12472
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24766 11872 24822 11928
rect 25226 11348 25282 11384
rect 25226 11328 25228 11348
rect 25228 11328 25280 11348
rect 25280 11328 25282 11348
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 25594 10240 25650 10296
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24674 9036 24730 9072
rect 24674 9016 24676 9036
rect 24676 9016 24728 9036
rect 24728 9016 24730 9036
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24766 8880 24822 8936
rect 24674 8472 24730 8528
rect 23846 7248 23902 7304
rect 24766 7928 24822 7984
rect 24122 7792 24178 7848
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 25226 6860 25282 6896
rect 25226 6840 25228 6860
rect 25228 6840 25280 6860
rect 25280 6840 25282 6860
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 23846 4700 23848 4720
rect 23848 4700 23900 4720
rect 23900 4700 23902 4720
rect 23846 4664 23902 4700
rect 23754 3576 23810 3632
rect 24674 6024 24730 6080
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24030 3984 24086 4040
rect 23754 3304 23810 3360
rect 23570 3168 23626 3224
rect 23938 3440 23994 3496
rect 24122 3712 24178 3768
rect 24030 1536 24086 1592
rect 23570 856 23626 912
rect 24950 4392 25006 4448
rect 25410 4120 25466 4176
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24766 2896 24822 2952
rect 27526 2896 27582 2952
rect 25502 2760 25558 2816
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24582 1264 24638 1320
rect 24766 1264 24822 1320
rect 26790 1400 26846 1456
rect 24582 312 24638 368
<< metal3 >>
rect 23197 27706 23263 27709
rect 27520 27706 28000 27736
rect 23197 27704 28000 27706
rect 23197 27648 23202 27704
rect 23258 27648 28000 27704
rect 23197 27646 28000 27648
rect 23197 27643 23263 27646
rect 27520 27616 28000 27646
rect 24209 27162 24275 27165
rect 27520 27162 28000 27192
rect 24209 27160 28000 27162
rect 24209 27104 24214 27160
rect 24270 27104 28000 27160
rect 24209 27102 28000 27104
rect 24209 27099 24275 27102
rect 27520 27072 28000 27102
rect 23289 26618 23355 26621
rect 27520 26618 28000 26648
rect 23289 26616 28000 26618
rect 23289 26560 23294 26616
rect 23350 26560 28000 26616
rect 23289 26558 28000 26560
rect 23289 26555 23355 26558
rect 27520 26528 28000 26558
rect 23657 25938 23723 25941
rect 27520 25938 28000 25968
rect 23657 25936 28000 25938
rect 23657 25880 23662 25936
rect 23718 25880 28000 25936
rect 23657 25878 28000 25880
rect 23657 25875 23723 25878
rect 27520 25848 28000 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24761 25394 24827 25397
rect 27520 25394 28000 25424
rect 24761 25392 28000 25394
rect 24761 25336 24766 25392
rect 24822 25336 28000 25392
rect 24761 25334 28000 25336
rect 24761 25331 24827 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 2957 24850 3023 24853
rect 12341 24850 12407 24853
rect 2957 24848 12407 24850
rect 2957 24792 2962 24848
rect 3018 24792 12346 24848
rect 12402 24792 12407 24848
rect 2957 24790 12407 24792
rect 2957 24787 3023 24790
rect 12341 24787 12407 24790
rect 14549 24850 14615 24853
rect 15929 24850 15995 24853
rect 14549 24848 15995 24850
rect 14549 24792 14554 24848
rect 14610 24792 15934 24848
rect 15990 24792 15995 24848
rect 14549 24790 15995 24792
rect 14549 24787 14615 24790
rect 15929 24787 15995 24790
rect 20161 24850 20227 24853
rect 21357 24850 21423 24853
rect 20161 24848 21423 24850
rect 20161 24792 20166 24848
rect 20222 24792 21362 24848
rect 21418 24792 21423 24848
rect 20161 24790 21423 24792
rect 20161 24787 20227 24790
rect 21357 24787 21423 24790
rect 23749 24850 23815 24853
rect 27520 24850 28000 24880
rect 23749 24848 28000 24850
rect 23749 24792 23754 24848
rect 23810 24792 28000 24848
rect 23749 24790 28000 24792
rect 23749 24787 23815 24790
rect 27520 24760 28000 24790
rect 1577 24714 1643 24717
rect 12985 24714 13051 24717
rect 14457 24714 14523 24717
rect 1577 24712 12818 24714
rect 1577 24656 1582 24712
rect 1638 24656 12818 24712
rect 1577 24654 12818 24656
rect 1577 24651 1643 24654
rect 12758 24578 12818 24654
rect 12985 24712 14523 24714
rect 12985 24656 12990 24712
rect 13046 24656 14462 24712
rect 14518 24656 14523 24712
rect 12985 24654 14523 24656
rect 12985 24651 13051 24654
rect 14457 24651 14523 24654
rect 21265 24714 21331 24717
rect 23473 24714 23539 24717
rect 21265 24712 23539 24714
rect 21265 24656 21270 24712
rect 21326 24656 23478 24712
rect 23534 24656 23539 24712
rect 21265 24654 23539 24656
rect 21265 24651 21331 24654
rect 23473 24651 23539 24654
rect 15377 24578 15443 24581
rect 12758 24576 15443 24578
rect 12758 24520 15382 24576
rect 15438 24520 15443 24576
rect 12758 24518 15443 24520
rect 15377 24515 15443 24518
rect 23657 24578 23723 24581
rect 25497 24578 25563 24581
rect 23657 24576 25563 24578
rect 23657 24520 23662 24576
rect 23718 24520 25502 24576
rect 25558 24520 25563 24576
rect 23657 24518 25563 24520
rect 23657 24515 23723 24518
rect 25497 24515 25563 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 11881 24442 11947 24445
rect 13537 24442 13603 24445
rect 11881 24440 13603 24442
rect 11881 24384 11886 24440
rect 11942 24384 13542 24440
rect 13598 24384 13603 24440
rect 11881 24382 13603 24384
rect 11881 24379 11947 24382
rect 13537 24379 13603 24382
rect 24761 24442 24827 24445
rect 26877 24442 26943 24445
rect 24761 24440 26943 24442
rect 24761 24384 24766 24440
rect 24822 24384 26882 24440
rect 26938 24384 26943 24440
rect 24761 24382 26943 24384
rect 24761 24379 24827 24382
rect 26877 24379 26943 24382
rect 23933 24306 23999 24309
rect 23933 24304 24962 24306
rect 23933 24248 23938 24304
rect 23994 24248 24962 24304
rect 23933 24246 24962 24248
rect 23933 24243 23999 24246
rect 4981 24170 5047 24173
rect 11513 24170 11579 24173
rect 4981 24168 11579 24170
rect 4981 24112 4986 24168
rect 5042 24112 11518 24168
rect 11574 24112 11579 24168
rect 4981 24110 11579 24112
rect 4981 24107 5047 24110
rect 11513 24107 11579 24110
rect 22645 24170 22711 24173
rect 24669 24170 24735 24173
rect 22645 24168 24735 24170
rect 22645 24112 22650 24168
rect 22706 24112 24674 24168
rect 24730 24112 24735 24168
rect 22645 24110 24735 24112
rect 24902 24170 24962 24246
rect 27520 24170 28000 24200
rect 24902 24110 28000 24170
rect 22645 24107 22711 24110
rect 24669 24107 24735 24110
rect 27520 24080 28000 24110
rect 15653 24034 15719 24037
rect 20621 24034 20687 24037
rect 15653 24032 20687 24034
rect 15653 23976 15658 24032
rect 15714 23976 20626 24032
rect 20682 23976 20687 24032
rect 15653 23974 20687 23976
rect 15653 23971 15719 23974
rect 20621 23971 20687 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 6361 23898 6427 23901
rect 11421 23898 11487 23901
rect 14549 23898 14615 23901
rect 6361 23896 11487 23898
rect 6361 23840 6366 23896
rect 6422 23840 11426 23896
rect 11482 23840 11487 23896
rect 6361 23838 11487 23840
rect 6361 23835 6427 23838
rect 11421 23835 11487 23838
rect 12942 23896 14615 23898
rect 12942 23840 14554 23896
rect 14610 23840 14615 23896
rect 12942 23838 14615 23840
rect 4337 23762 4403 23765
rect 12942 23762 13002 23838
rect 14549 23835 14615 23838
rect 17033 23898 17099 23901
rect 19425 23898 19491 23901
rect 17033 23896 19491 23898
rect 17033 23840 17038 23896
rect 17094 23840 19430 23896
rect 19486 23840 19491 23896
rect 17033 23838 19491 23840
rect 17033 23835 17099 23838
rect 19425 23835 19491 23838
rect 24761 23898 24827 23901
rect 27521 23898 27587 23901
rect 24761 23896 27587 23898
rect 24761 23840 24766 23896
rect 24822 23840 27526 23896
rect 27582 23840 27587 23896
rect 24761 23838 27587 23840
rect 24761 23835 24827 23838
rect 27521 23835 27587 23838
rect 4337 23760 13002 23762
rect 4337 23704 4342 23760
rect 4398 23704 13002 23760
rect 4337 23702 13002 23704
rect 13169 23762 13235 23765
rect 16113 23762 16179 23765
rect 13169 23760 16179 23762
rect 13169 23704 13174 23760
rect 13230 23704 16118 23760
rect 16174 23704 16179 23760
rect 13169 23702 16179 23704
rect 4337 23699 4403 23702
rect 13169 23699 13235 23702
rect 16113 23699 16179 23702
rect 17769 23762 17835 23765
rect 20529 23762 20595 23765
rect 17769 23760 20595 23762
rect 17769 23704 17774 23760
rect 17830 23704 20534 23760
rect 20590 23704 20595 23760
rect 17769 23702 20595 23704
rect 17769 23699 17835 23702
rect 20529 23699 20595 23702
rect 12525 23626 12591 23629
rect 16297 23626 16363 23629
rect 12525 23624 16363 23626
rect 12525 23568 12530 23624
rect 12586 23568 16302 23624
rect 16358 23568 16363 23624
rect 12525 23566 16363 23568
rect 12525 23563 12591 23566
rect 16297 23563 16363 23566
rect 18137 23626 18203 23629
rect 20897 23626 20963 23629
rect 18137 23624 20963 23626
rect 18137 23568 18142 23624
rect 18198 23568 20902 23624
rect 20958 23568 20963 23624
rect 18137 23566 20963 23568
rect 18137 23563 18203 23566
rect 20897 23563 20963 23566
rect 23657 23626 23723 23629
rect 27520 23626 28000 23656
rect 23657 23624 28000 23626
rect 23657 23568 23662 23624
rect 23718 23568 28000 23624
rect 23657 23566 28000 23568
rect 23657 23563 23723 23566
rect 27520 23536 28000 23566
rect 17033 23490 17099 23493
rect 18689 23490 18755 23493
rect 17033 23488 18755 23490
rect 17033 23432 17038 23488
rect 17094 23432 18694 23488
rect 18750 23432 18755 23488
rect 17033 23430 18755 23432
rect 17033 23427 17099 23430
rect 18689 23427 18755 23430
rect 24669 23490 24735 23493
rect 26141 23490 26207 23493
rect 24669 23488 26207 23490
rect 24669 23432 24674 23488
rect 24730 23432 26146 23488
rect 26202 23432 26207 23488
rect 24669 23430 26207 23432
rect 24669 23427 24735 23430
rect 26141 23427 26207 23430
rect 10277 23424 10597 23425
rect 0 23354 480 23384
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 22737 23354 22803 23357
rect 23841 23354 23907 23357
rect 0 23294 1226 23354
rect 0 23264 480 23294
rect 1166 22402 1226 23294
rect 22737 23352 23907 23354
rect 22737 23296 22742 23352
rect 22798 23296 23846 23352
rect 23902 23296 23907 23352
rect 22737 23294 23907 23296
rect 22737 23291 22803 23294
rect 23841 23291 23907 23294
rect 10685 23218 10751 23221
rect 12525 23218 12591 23221
rect 22921 23218 22987 23221
rect 10685 23216 22987 23218
rect 10685 23160 10690 23216
rect 10746 23160 12530 23216
rect 12586 23160 22926 23216
rect 22982 23160 22987 23216
rect 10685 23158 22987 23160
rect 10685 23155 10751 23158
rect 12525 23155 12591 23158
rect 22921 23155 22987 23158
rect 14457 23082 14523 23085
rect 20713 23082 20779 23085
rect 14457 23080 20779 23082
rect 14457 23024 14462 23080
rect 14518 23024 20718 23080
rect 20774 23024 20779 23080
rect 14457 23022 20779 23024
rect 14457 23019 14523 23022
rect 20713 23019 20779 23022
rect 20989 23082 21055 23085
rect 24209 23082 24275 23085
rect 20989 23080 24275 23082
rect 20989 23024 20994 23080
rect 21050 23024 24214 23080
rect 24270 23024 24275 23080
rect 20989 23022 24275 23024
rect 20989 23019 21055 23022
rect 24209 23019 24275 23022
rect 25405 23082 25471 23085
rect 27520 23082 28000 23112
rect 25405 23080 28000 23082
rect 25405 23024 25410 23080
rect 25466 23024 28000 23080
rect 25405 23022 28000 23024
rect 25405 23019 25471 23022
rect 27520 22992 28000 23022
rect 15469 22946 15535 22949
rect 21081 22946 21147 22949
rect 15469 22944 21147 22946
rect 15469 22888 15474 22944
rect 15530 22888 21086 22944
rect 21142 22888 21147 22944
rect 15469 22886 21147 22888
rect 15469 22883 15535 22886
rect 21081 22883 21147 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1485 22674 1551 22677
rect 16481 22674 16547 22677
rect 1485 22672 16547 22674
rect 1485 22616 1490 22672
rect 1546 22616 16486 22672
rect 16542 22616 16547 22672
rect 1485 22614 16547 22616
rect 1485 22611 1551 22614
rect 16481 22611 16547 22614
rect 3693 22538 3759 22541
rect 17401 22538 17467 22541
rect 19149 22538 19215 22541
rect 23933 22538 23999 22541
rect 27520 22538 28000 22568
rect 3693 22536 17467 22538
rect 3693 22480 3698 22536
rect 3754 22480 17406 22536
rect 17462 22480 17467 22536
rect 3693 22478 17467 22480
rect 3693 22475 3759 22478
rect 17401 22475 17467 22478
rect 17542 22536 23999 22538
rect 17542 22480 19154 22536
rect 19210 22480 23938 22536
rect 23994 22480 23999 22536
rect 17542 22478 23999 22480
rect 15377 22402 15443 22405
rect 17542 22402 17602 22478
rect 19149 22475 19215 22478
rect 23933 22475 23999 22478
rect 24902 22478 28000 22538
rect 1166 22342 2698 22402
rect 2638 22266 2698 22342
rect 15377 22400 17602 22402
rect 15377 22344 15382 22400
rect 15438 22344 17602 22400
rect 15377 22342 17602 22344
rect 20069 22402 20135 22405
rect 23289 22402 23355 22405
rect 20069 22400 23355 22402
rect 20069 22344 20074 22400
rect 20130 22344 23294 22400
rect 23350 22344 23355 22400
rect 20069 22342 23355 22344
rect 15377 22339 15443 22342
rect 20069 22339 20135 22342
rect 23289 22339 23355 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 9949 22266 10015 22269
rect 2638 22264 10015 22266
rect 2638 22208 9954 22264
rect 10010 22208 10015 22264
rect 2638 22206 10015 22208
rect 9949 22203 10015 22206
rect 14089 22130 14155 22133
rect 24902 22130 24962 22478
rect 27520 22448 28000 22478
rect 14089 22128 24962 22130
rect 14089 22072 14094 22128
rect 14150 22072 24962 22128
rect 14089 22070 24962 22072
rect 14089 22067 14155 22070
rect 15285 21994 15351 21997
rect 18505 21994 18571 21997
rect 15285 21992 18571 21994
rect 15285 21936 15290 21992
rect 15346 21936 18510 21992
rect 18566 21936 18571 21992
rect 15285 21934 18571 21936
rect 15285 21931 15351 21934
rect 18505 21931 18571 21934
rect 16021 21858 16087 21861
rect 23473 21858 23539 21861
rect 16021 21856 23539 21858
rect 16021 21800 16026 21856
rect 16082 21800 23478 21856
rect 23534 21800 23539 21856
rect 16021 21798 23539 21800
rect 16021 21795 16087 21798
rect 23473 21795 23539 21798
rect 24761 21858 24827 21861
rect 27520 21858 28000 21888
rect 24761 21856 28000 21858
rect 24761 21800 24766 21856
rect 24822 21800 28000 21856
rect 24761 21798 28000 21800
rect 24761 21795 24827 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 27520 21768 28000 21798
rect 24277 21727 24597 21728
rect 5993 21722 6059 21725
rect 11053 21722 11119 21725
rect 5993 21720 11119 21722
rect 5993 21664 5998 21720
rect 6054 21664 11058 21720
rect 11114 21664 11119 21720
rect 5993 21662 11119 21664
rect 5993 21659 6059 21662
rect 11053 21659 11119 21662
rect 22553 21314 22619 21317
rect 27520 21314 28000 21344
rect 22553 21312 28000 21314
rect 22553 21256 22558 21312
rect 22614 21256 28000 21312
rect 22553 21254 28000 21256
rect 22553 21251 22619 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 27520 21224 28000 21254
rect 19610 21183 19930 21184
rect 9765 21042 9831 21045
rect 11697 21042 11763 21045
rect 9765 21040 11763 21042
rect 9765 20984 9770 21040
rect 9826 20984 11702 21040
rect 11758 20984 11763 21040
rect 9765 20982 11763 20984
rect 9765 20979 9831 20982
rect 11697 20979 11763 20982
rect 13629 21042 13695 21045
rect 24209 21042 24275 21045
rect 13629 21040 24275 21042
rect 13629 20984 13634 21040
rect 13690 20984 24214 21040
rect 24270 20984 24275 21040
rect 13629 20982 24275 20984
rect 13629 20979 13695 20982
rect 24209 20979 24275 20982
rect 1577 20906 1643 20909
rect 14089 20906 14155 20909
rect 1577 20904 14155 20906
rect 1577 20848 1582 20904
rect 1638 20848 14094 20904
rect 14150 20848 14155 20904
rect 1577 20846 14155 20848
rect 1577 20843 1643 20846
rect 14089 20843 14155 20846
rect 9121 20770 9187 20773
rect 14089 20770 14155 20773
rect 9121 20768 14155 20770
rect 9121 20712 9126 20768
rect 9182 20712 14094 20768
rect 14150 20712 14155 20768
rect 9121 20710 14155 20712
rect 9121 20707 9187 20710
rect 14089 20707 14155 20710
rect 18781 20770 18847 20773
rect 21909 20770 21975 20773
rect 18781 20768 21975 20770
rect 18781 20712 18786 20768
rect 18842 20712 21914 20768
rect 21970 20712 21975 20768
rect 18781 20710 21975 20712
rect 18781 20707 18847 20710
rect 21909 20707 21975 20710
rect 24761 20770 24827 20773
rect 27520 20770 28000 20800
rect 24761 20768 28000 20770
rect 24761 20712 24766 20768
rect 24822 20712 28000 20768
rect 24761 20710 28000 20712
rect 24761 20707 24827 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 10317 20498 10383 20501
rect 15653 20498 15719 20501
rect 16573 20498 16639 20501
rect 10317 20496 16639 20498
rect 10317 20440 10322 20496
rect 10378 20440 15658 20496
rect 15714 20440 16578 20496
rect 16634 20440 16639 20496
rect 10317 20438 16639 20440
rect 10317 20435 10383 20438
rect 15653 20435 15719 20438
rect 16573 20435 16639 20438
rect 1577 20362 1643 20365
rect 24669 20362 24735 20365
rect 1577 20360 24735 20362
rect 1577 20304 1582 20360
rect 1638 20304 24674 20360
rect 24730 20304 24735 20360
rect 1577 20302 24735 20304
rect 1577 20299 1643 20302
rect 24669 20299 24735 20302
rect 12709 20226 12775 20229
rect 14181 20226 14247 20229
rect 12709 20224 14247 20226
rect 12709 20168 12714 20224
rect 12770 20168 14186 20224
rect 14242 20168 14247 20224
rect 12709 20166 14247 20168
rect 12709 20163 12775 20166
rect 14181 20163 14247 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 13169 20090 13235 20093
rect 15745 20090 15811 20093
rect 16021 20090 16087 20093
rect 27520 20090 28000 20120
rect 13169 20088 16087 20090
rect 13169 20032 13174 20088
rect 13230 20032 15750 20088
rect 15806 20032 16026 20088
rect 16082 20032 16087 20088
rect 13169 20030 16087 20032
rect 13169 20027 13235 20030
rect 15745 20027 15811 20030
rect 16021 20027 16087 20030
rect 24902 20030 28000 20090
rect 12065 19954 12131 19957
rect 24761 19954 24827 19957
rect 12065 19952 24827 19954
rect 12065 19896 12070 19952
rect 12126 19896 24766 19952
rect 24822 19896 24827 19952
rect 12065 19894 24827 19896
rect 12065 19891 12131 19894
rect 24761 19891 24827 19894
rect 9949 19818 10015 19821
rect 15929 19818 15995 19821
rect 24902 19818 24962 20030
rect 27520 20000 28000 20030
rect 9949 19816 15394 19818
rect 9949 19760 9954 19816
rect 10010 19760 15394 19816
rect 9949 19758 15394 19760
rect 9949 19755 10015 19758
rect 15334 19682 15394 19758
rect 15929 19816 24962 19818
rect 15929 19760 15934 19816
rect 15990 19760 24962 19816
rect 15929 19758 24962 19760
rect 15929 19755 15995 19758
rect 21817 19682 21883 19685
rect 15334 19680 21883 19682
rect 15334 19624 21822 19680
rect 21878 19624 21883 19680
rect 15334 19622 21883 19624
rect 21817 19619 21883 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 27520 19546 28000 19576
rect 24718 19486 28000 19546
rect 18689 19410 18755 19413
rect 20437 19410 20503 19413
rect 18689 19408 20503 19410
rect 18689 19352 18694 19408
rect 18750 19352 20442 19408
rect 20498 19352 20503 19408
rect 18689 19350 20503 19352
rect 18689 19347 18755 19350
rect 20437 19347 20503 19350
rect 20621 19410 20687 19413
rect 23657 19410 23723 19413
rect 20621 19408 23723 19410
rect 20621 19352 20626 19408
rect 20682 19352 23662 19408
rect 23718 19352 23723 19408
rect 20621 19350 23723 19352
rect 20621 19347 20687 19350
rect 23657 19347 23723 19350
rect 24025 19410 24091 19413
rect 24718 19410 24778 19486
rect 27520 19456 28000 19486
rect 24025 19408 24778 19410
rect 24025 19352 24030 19408
rect 24086 19352 24778 19408
rect 24025 19350 24778 19352
rect 24025 19347 24091 19350
rect 7097 19274 7163 19277
rect 10777 19274 10843 19277
rect 7097 19272 10843 19274
rect 7097 19216 7102 19272
rect 7158 19216 10782 19272
rect 10838 19216 10843 19272
rect 7097 19214 10843 19216
rect 7097 19211 7163 19214
rect 10777 19211 10843 19214
rect 12433 19274 12499 19277
rect 12801 19274 12867 19277
rect 12433 19272 12867 19274
rect 12433 19216 12438 19272
rect 12494 19216 12806 19272
rect 12862 19216 12867 19272
rect 12433 19214 12867 19216
rect 12433 19211 12499 19214
rect 12801 19211 12867 19214
rect 13169 19138 13235 19141
rect 18597 19138 18663 19141
rect 13169 19136 18663 19138
rect 13169 19080 13174 19136
rect 13230 19080 18602 19136
rect 18658 19080 18663 19136
rect 13169 19078 18663 19080
rect 13169 19075 13235 19078
rect 18597 19075 18663 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 24669 19002 24735 19005
rect 27520 19002 28000 19032
rect 24669 19000 28000 19002
rect 24669 18944 24674 19000
rect 24730 18944 28000 19000
rect 24669 18942 28000 18944
rect 24669 18939 24735 18942
rect 27520 18912 28000 18942
rect 19793 18866 19859 18869
rect 20345 18866 20411 18869
rect 23933 18866 23999 18869
rect 19793 18864 23999 18866
rect 19793 18808 19798 18864
rect 19854 18808 20350 18864
rect 20406 18808 23938 18864
rect 23994 18808 23999 18864
rect 19793 18806 23999 18808
rect 19793 18803 19859 18806
rect 20345 18803 20411 18806
rect 23933 18803 23999 18806
rect 14089 18730 14155 18733
rect 19425 18730 19491 18733
rect 14089 18728 19491 18730
rect 14089 18672 14094 18728
rect 14150 18672 19430 18728
rect 19486 18672 19491 18728
rect 14089 18670 19491 18672
rect 14089 18667 14155 18670
rect 19425 18667 19491 18670
rect 16297 18594 16363 18597
rect 20110 18594 20116 18596
rect 16297 18592 20116 18594
rect 16297 18536 16302 18592
rect 16358 18536 20116 18592
rect 16297 18534 20116 18536
rect 16297 18531 16363 18534
rect 20110 18532 20116 18534
rect 20180 18594 20186 18596
rect 23197 18594 23263 18597
rect 20180 18592 23263 18594
rect 20180 18536 23202 18592
rect 23258 18536 23263 18592
rect 20180 18534 23263 18536
rect 20180 18532 20186 18534
rect 23197 18531 23263 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 18597 18458 18663 18461
rect 21265 18458 21331 18461
rect 18597 18456 21331 18458
rect 18597 18400 18602 18456
rect 18658 18400 21270 18456
rect 21326 18400 21331 18456
rect 18597 18398 21331 18400
rect 18597 18395 18663 18398
rect 21265 18395 21331 18398
rect 25681 18458 25747 18461
rect 27520 18458 28000 18488
rect 25681 18456 28000 18458
rect 25681 18400 25686 18456
rect 25742 18400 28000 18456
rect 25681 18398 28000 18400
rect 25681 18395 25747 18398
rect 27520 18368 28000 18398
rect 13353 18322 13419 18325
rect 15377 18322 15443 18325
rect 13353 18320 15443 18322
rect 13353 18264 13358 18320
rect 13414 18264 15382 18320
rect 15438 18264 15443 18320
rect 13353 18262 15443 18264
rect 13353 18259 13419 18262
rect 15377 18259 15443 18262
rect 19977 18322 20043 18325
rect 25221 18322 25287 18325
rect 19977 18320 25287 18322
rect 19977 18264 19982 18320
rect 20038 18264 25226 18320
rect 25282 18264 25287 18320
rect 19977 18262 25287 18264
rect 19977 18259 20043 18262
rect 25221 18259 25287 18262
rect 11697 18186 11763 18189
rect 22093 18186 22159 18189
rect 11697 18184 22159 18186
rect 11697 18128 11702 18184
rect 11758 18128 22098 18184
rect 22154 18128 22159 18184
rect 11697 18126 22159 18128
rect 11697 18123 11763 18126
rect 22093 18123 22159 18126
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 11237 17914 11303 17917
rect 13997 17914 14063 17917
rect 11237 17912 14063 17914
rect 11237 17856 11242 17912
rect 11298 17856 14002 17912
rect 14058 17856 14063 17912
rect 11237 17854 14063 17856
rect 11237 17851 11303 17854
rect 13997 17851 14063 17854
rect 20069 17914 20135 17917
rect 25497 17914 25563 17917
rect 20069 17912 25563 17914
rect 20069 17856 20074 17912
rect 20130 17856 25502 17912
rect 25558 17856 25563 17912
rect 20069 17854 25563 17856
rect 20069 17851 20135 17854
rect 25497 17851 25563 17854
rect 7741 17778 7807 17781
rect 14273 17778 14339 17781
rect 7741 17776 14339 17778
rect 7741 17720 7746 17776
rect 7802 17720 14278 17776
rect 14334 17720 14339 17776
rect 7741 17718 14339 17720
rect 7741 17715 7807 17718
rect 14273 17715 14339 17718
rect 16849 17778 16915 17781
rect 20161 17778 20227 17781
rect 16849 17776 20227 17778
rect 16849 17720 16854 17776
rect 16910 17720 20166 17776
rect 20222 17720 20227 17776
rect 16849 17718 20227 17720
rect 16849 17715 16915 17718
rect 20161 17715 20227 17718
rect 25405 17778 25471 17781
rect 27520 17778 28000 17808
rect 25405 17776 28000 17778
rect 25405 17720 25410 17776
rect 25466 17720 28000 17776
rect 25405 17718 28000 17720
rect 25405 17715 25471 17718
rect 27520 17688 28000 17718
rect 17953 17642 18019 17645
rect 15518 17640 18019 17642
rect 15518 17584 17958 17640
rect 18014 17584 18019 17640
rect 15518 17582 18019 17584
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 10869 17234 10935 17237
rect 15518 17234 15578 17582
rect 17953 17579 18019 17582
rect 19793 17642 19859 17645
rect 20345 17642 20411 17645
rect 23197 17642 23263 17645
rect 19793 17640 23263 17642
rect 19793 17584 19798 17640
rect 19854 17584 20350 17640
rect 20406 17584 23202 17640
rect 23258 17584 23263 17640
rect 19793 17582 23263 17584
rect 19793 17579 19859 17582
rect 20345 17579 20411 17582
rect 23197 17579 23263 17582
rect 15653 17506 15719 17509
rect 21633 17506 21699 17509
rect 15653 17504 21699 17506
rect 15653 17448 15658 17504
rect 15714 17448 21638 17504
rect 21694 17448 21699 17504
rect 15653 17446 21699 17448
rect 15653 17443 15719 17446
rect 21633 17443 21699 17446
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 16021 17370 16087 17373
rect 19977 17370 20043 17373
rect 16021 17368 20043 17370
rect 16021 17312 16026 17368
rect 16082 17312 19982 17368
rect 20038 17312 20043 17368
rect 16021 17310 20043 17312
rect 16021 17307 16087 17310
rect 19977 17307 20043 17310
rect 10869 17232 15578 17234
rect 10869 17176 10874 17232
rect 10930 17176 15578 17232
rect 10869 17174 15578 17176
rect 19057 17234 19123 17237
rect 20253 17234 20319 17237
rect 22277 17234 22343 17237
rect 19057 17232 22343 17234
rect 19057 17176 19062 17232
rect 19118 17176 20258 17232
rect 20314 17176 22282 17232
rect 22338 17176 22343 17232
rect 19057 17174 22343 17176
rect 10869 17171 10935 17174
rect 19057 17171 19123 17174
rect 20253 17171 20319 17174
rect 22277 17171 22343 17174
rect 24945 17234 25011 17237
rect 27520 17234 28000 17264
rect 24945 17232 28000 17234
rect 24945 17176 24950 17232
rect 25006 17176 28000 17232
rect 24945 17174 28000 17176
rect 24945 17171 25011 17174
rect 27520 17144 28000 17174
rect 17401 17098 17467 17101
rect 23197 17098 23263 17101
rect 17401 17096 23263 17098
rect 17401 17040 17406 17096
rect 17462 17040 23202 17096
rect 23258 17040 23263 17096
rect 17401 17038 23263 17040
rect 17401 17035 17467 17038
rect 23197 17035 23263 17038
rect 14273 16962 14339 16965
rect 14406 16962 14412 16964
rect 14273 16960 14412 16962
rect 14273 16904 14278 16960
rect 14334 16904 14412 16960
rect 14273 16902 14412 16904
rect 14273 16899 14339 16902
rect 14406 16900 14412 16902
rect 14476 16900 14482 16964
rect 15469 16962 15535 16965
rect 19333 16962 19399 16965
rect 15469 16960 19399 16962
rect 15469 16904 15474 16960
rect 15530 16904 19338 16960
rect 19394 16904 19399 16960
rect 15469 16902 19399 16904
rect 15469 16899 15535 16902
rect 19333 16899 19399 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 18229 16690 18295 16693
rect 25037 16690 25103 16693
rect 18229 16688 25103 16690
rect 18229 16632 18234 16688
rect 18290 16632 25042 16688
rect 25098 16632 25103 16688
rect 18229 16630 25103 16632
rect 18229 16627 18295 16630
rect 25037 16627 25103 16630
rect 25221 16690 25287 16693
rect 27520 16690 28000 16720
rect 25221 16688 28000 16690
rect 25221 16632 25226 16688
rect 25282 16632 28000 16688
rect 25221 16630 28000 16632
rect 25221 16627 25287 16630
rect 27520 16600 28000 16630
rect 13353 16554 13419 16557
rect 15561 16554 15627 16557
rect 13353 16552 15627 16554
rect 13353 16496 13358 16552
rect 13414 16496 15566 16552
rect 15622 16496 15627 16552
rect 13353 16494 15627 16496
rect 13353 16491 13419 16494
rect 15561 16491 15627 16494
rect 17217 16418 17283 16421
rect 20989 16418 21055 16421
rect 17217 16416 21055 16418
rect 17217 16360 17222 16416
rect 17278 16360 20994 16416
rect 21050 16360 21055 16416
rect 17217 16358 21055 16360
rect 17217 16355 17283 16358
rect 20989 16355 21055 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 9581 16146 9647 16149
rect 14733 16146 14799 16149
rect 9581 16144 14799 16146
rect 9581 16088 9586 16144
rect 9642 16088 14738 16144
rect 14794 16088 14799 16144
rect 9581 16086 14799 16088
rect 9581 16083 9647 16086
rect 14733 16083 14799 16086
rect 16757 16146 16823 16149
rect 20529 16146 20595 16149
rect 16757 16144 20595 16146
rect 16757 16088 16762 16144
rect 16818 16088 20534 16144
rect 20590 16088 20595 16144
rect 16757 16086 20595 16088
rect 16757 16083 16823 16086
rect 20529 16083 20595 16086
rect 13537 16010 13603 16013
rect 24577 16010 24643 16013
rect 13537 16008 24643 16010
rect 13537 15952 13542 16008
rect 13598 15952 24582 16008
rect 24638 15952 24643 16008
rect 13537 15950 24643 15952
rect 13537 15947 13603 15950
rect 24577 15947 24643 15950
rect 24761 16010 24827 16013
rect 27520 16010 28000 16040
rect 24761 16008 28000 16010
rect 24761 15952 24766 16008
rect 24822 15952 28000 16008
rect 24761 15950 28000 15952
rect 24761 15947 24827 15950
rect 27520 15920 28000 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 15193 15738 15259 15741
rect 15193 15736 18476 15738
rect 15193 15680 15198 15736
rect 15254 15680 18476 15736
rect 15193 15678 18476 15680
rect 15193 15675 15259 15678
rect 16205 15602 16271 15605
rect 18229 15602 18295 15605
rect 16205 15600 18295 15602
rect 16205 15544 16210 15600
rect 16266 15544 18234 15600
rect 18290 15544 18295 15600
rect 16205 15542 18295 15544
rect 18416 15602 18476 15678
rect 20713 15602 20779 15605
rect 18416 15600 20779 15602
rect 18416 15544 20718 15600
rect 20774 15544 20779 15600
rect 18416 15542 20779 15544
rect 16205 15539 16271 15542
rect 18229 15539 18295 15542
rect 20713 15539 20779 15542
rect 15101 15466 15167 15469
rect 24577 15466 24643 15469
rect 15101 15464 24643 15466
rect 15101 15408 15106 15464
rect 15162 15408 24582 15464
rect 24638 15408 24643 15464
rect 15101 15406 24643 15408
rect 15101 15403 15167 15406
rect 24577 15403 24643 15406
rect 24761 15466 24827 15469
rect 27520 15466 28000 15496
rect 24761 15464 28000 15466
rect 24761 15408 24766 15464
rect 24822 15408 28000 15464
rect 24761 15406 28000 15408
rect 24761 15403 24827 15406
rect 27520 15376 28000 15406
rect 20302 15270 21466 15330
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 9489 15194 9555 15197
rect 14181 15194 14247 15197
rect 9489 15192 14247 15194
rect 9489 15136 9494 15192
rect 9550 15136 14186 15192
rect 14242 15136 14247 15192
rect 9489 15134 14247 15136
rect 9489 15131 9555 15134
rect 14181 15131 14247 15134
rect 15745 15194 15811 15197
rect 20302 15194 20362 15270
rect 15745 15192 20362 15194
rect 15745 15136 15750 15192
rect 15806 15136 20362 15192
rect 15745 15134 20362 15136
rect 20437 15194 20503 15197
rect 21265 15194 21331 15197
rect 20437 15192 21331 15194
rect 20437 15136 20442 15192
rect 20498 15136 21270 15192
rect 21326 15136 21331 15192
rect 20437 15134 21331 15136
rect 21406 15194 21466 15270
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 23565 15194 23631 15197
rect 23841 15194 23907 15197
rect 21406 15192 23907 15194
rect 21406 15136 23570 15192
rect 23626 15136 23846 15192
rect 23902 15136 23907 15192
rect 21406 15134 23907 15136
rect 15745 15131 15811 15134
rect 20437 15131 20503 15134
rect 21265 15131 21331 15134
rect 23565 15131 23631 15134
rect 23841 15131 23907 15134
rect 13721 15058 13787 15061
rect 24577 15058 24643 15061
rect 13721 15056 24643 15058
rect 13721 15000 13726 15056
rect 13782 15000 24582 15056
rect 24638 15000 24643 15056
rect 13721 14998 24643 15000
rect 13721 14995 13787 14998
rect 24577 14995 24643 14998
rect 19057 14922 19123 14925
rect 21357 14922 21423 14925
rect 19057 14920 21423 14922
rect 19057 14864 19062 14920
rect 19118 14864 21362 14920
rect 21418 14864 21423 14920
rect 19057 14862 21423 14864
rect 19057 14859 19123 14862
rect 21357 14859 21423 14862
rect 24761 14922 24827 14925
rect 27520 14922 28000 14952
rect 24761 14920 28000 14922
rect 24761 14864 24766 14920
rect 24822 14864 28000 14920
rect 24761 14862 28000 14864
rect 24761 14859 24827 14862
rect 27520 14832 28000 14862
rect 13445 14786 13511 14789
rect 15745 14786 15811 14789
rect 13445 14784 15811 14786
rect 13445 14728 13450 14784
rect 13506 14728 15750 14784
rect 15806 14728 15811 14784
rect 13445 14726 15811 14728
rect 13445 14723 13511 14726
rect 15745 14723 15811 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 10777 14650 10843 14653
rect 15469 14650 15535 14653
rect 10777 14648 15535 14650
rect 10777 14592 10782 14648
rect 10838 14592 15474 14648
rect 15530 14592 15535 14648
rect 10777 14590 15535 14592
rect 10777 14587 10843 14590
rect 15469 14587 15535 14590
rect 11605 14514 11671 14517
rect 14089 14514 14155 14517
rect 11605 14512 14155 14514
rect 11605 14456 11610 14512
rect 11666 14456 14094 14512
rect 14150 14456 14155 14512
rect 11605 14454 14155 14456
rect 11605 14451 11671 14454
rect 14089 14451 14155 14454
rect 11605 14378 11671 14381
rect 13261 14378 13327 14381
rect 11605 14376 13327 14378
rect 11605 14320 11610 14376
rect 11666 14320 13266 14376
rect 13322 14320 13327 14376
rect 11605 14318 13327 14320
rect 11605 14315 11671 14318
rect 13261 14315 13327 14318
rect 14273 14378 14339 14381
rect 27520 14378 28000 14408
rect 14273 14376 28000 14378
rect 14273 14320 14278 14376
rect 14334 14320 28000 14376
rect 14273 14318 28000 14320
rect 14273 14315 14339 14318
rect 27520 14288 28000 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 19149 14106 19215 14109
rect 22185 14106 22251 14109
rect 19149 14104 22251 14106
rect 19149 14048 19154 14104
rect 19210 14048 22190 14104
rect 22246 14048 22251 14104
rect 19149 14046 22251 14048
rect 19149 14043 19215 14046
rect 22185 14043 22251 14046
rect 0 13970 480 14000
rect 1669 13970 1735 13973
rect 0 13968 1735 13970
rect 0 13912 1674 13968
rect 1730 13912 1735 13968
rect 0 13910 1735 13912
rect 0 13880 480 13910
rect 1669 13907 1735 13910
rect 13261 13970 13327 13973
rect 25037 13970 25103 13973
rect 13261 13968 25103 13970
rect 13261 13912 13266 13968
rect 13322 13912 25042 13968
rect 25098 13912 25103 13968
rect 13261 13910 25103 13912
rect 13261 13907 13327 13910
rect 25037 13907 25103 13910
rect 13997 13834 14063 13837
rect 15561 13834 15627 13837
rect 13997 13832 15627 13834
rect 13997 13776 14002 13832
rect 14058 13776 15566 13832
rect 15622 13776 15627 13832
rect 13997 13774 15627 13776
rect 13997 13771 14063 13774
rect 15561 13771 15627 13774
rect 21081 13834 21147 13837
rect 24761 13834 24827 13837
rect 21081 13832 24827 13834
rect 21081 13776 21086 13832
rect 21142 13776 24766 13832
rect 24822 13776 24827 13832
rect 21081 13774 24827 13776
rect 21081 13771 21147 13774
rect 24761 13771 24827 13774
rect 20713 13698 20779 13701
rect 23105 13698 23171 13701
rect 20713 13696 23171 13698
rect 20713 13640 20718 13696
rect 20774 13640 23110 13696
rect 23166 13640 23171 13696
rect 20713 13638 23171 13640
rect 20713 13635 20779 13638
rect 23105 13635 23171 13638
rect 25405 13698 25471 13701
rect 27520 13698 28000 13728
rect 25405 13696 28000 13698
rect 25405 13640 25410 13696
rect 25466 13640 28000 13696
rect 25405 13638 28000 13640
rect 25405 13635 25471 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 27520 13608 28000 13638
rect 19610 13567 19930 13568
rect 22921 13562 22987 13565
rect 20072 13560 22987 13562
rect 20072 13504 22926 13560
rect 22982 13504 22987 13560
rect 20072 13502 22987 13504
rect 14181 13426 14247 13429
rect 20072 13426 20132 13502
rect 22921 13499 22987 13502
rect 14181 13424 20132 13426
rect 14181 13368 14186 13424
rect 14242 13368 20132 13424
rect 14181 13366 20132 13368
rect 21541 13426 21607 13429
rect 24577 13426 24643 13429
rect 21541 13424 24643 13426
rect 21541 13368 21546 13424
rect 21602 13368 24582 13424
rect 24638 13368 24643 13424
rect 21541 13366 24643 13368
rect 14181 13363 14247 13366
rect 21541 13363 21607 13366
rect 24577 13363 24643 13366
rect 2313 13290 2379 13293
rect 13077 13290 13143 13293
rect 2313 13288 13143 13290
rect 2313 13232 2318 13288
rect 2374 13232 13082 13288
rect 13138 13232 13143 13288
rect 2313 13230 13143 13232
rect 2313 13227 2379 13230
rect 13077 13227 13143 13230
rect 14273 13290 14339 13293
rect 17033 13290 17099 13293
rect 14273 13288 17099 13290
rect 14273 13232 14278 13288
rect 14334 13232 17038 13288
rect 17094 13232 17099 13288
rect 14273 13230 17099 13232
rect 14273 13227 14339 13230
rect 17033 13227 17099 13230
rect 24761 13154 24827 13157
rect 27520 13154 28000 13184
rect 24761 13152 28000 13154
rect 24761 13096 24766 13152
rect 24822 13096 28000 13152
rect 24761 13094 28000 13096
rect 24761 13091 24827 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 13077 12882 13143 12885
rect 18873 12882 18939 12885
rect 13077 12880 18939 12882
rect 13077 12824 13082 12880
rect 13138 12824 18878 12880
rect 18934 12824 18939 12880
rect 13077 12822 18939 12824
rect 13077 12819 13143 12822
rect 18873 12819 18939 12822
rect 13353 12746 13419 12749
rect 20805 12746 20871 12749
rect 23657 12746 23723 12749
rect 13353 12744 23723 12746
rect 13353 12688 13358 12744
rect 13414 12688 20810 12744
rect 20866 12688 23662 12744
rect 23718 12688 23723 12744
rect 13353 12686 23723 12688
rect 13353 12683 13419 12686
rect 20805 12683 20871 12686
rect 23657 12683 23723 12686
rect 12341 12610 12407 12613
rect 13905 12610 13971 12613
rect 12341 12608 13971 12610
rect 12341 12552 12346 12608
rect 12402 12552 13910 12608
rect 13966 12552 13971 12608
rect 12341 12550 13971 12552
rect 12341 12547 12407 12550
rect 13905 12547 13971 12550
rect 24761 12610 24827 12613
rect 27520 12610 28000 12640
rect 24761 12608 28000 12610
rect 24761 12552 24766 12608
rect 24822 12552 28000 12608
rect 24761 12550 28000 12552
rect 24761 12547 24827 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 23197 12474 23263 12477
rect 25405 12474 25471 12477
rect 23197 12472 25471 12474
rect 23197 12416 23202 12472
rect 23258 12416 25410 12472
rect 25466 12416 25471 12472
rect 23197 12414 25471 12416
rect 23197 12411 23263 12414
rect 25405 12411 25471 12414
rect 16205 12338 16271 12341
rect 18137 12338 18203 12341
rect 16205 12336 18203 12338
rect 16205 12280 16210 12336
rect 16266 12280 18142 12336
rect 18198 12280 18203 12336
rect 16205 12278 18203 12280
rect 16205 12275 16271 12278
rect 18137 12275 18203 12278
rect 20110 12276 20116 12340
rect 20180 12338 20186 12340
rect 20253 12338 20319 12341
rect 20180 12336 20319 12338
rect 20180 12280 20258 12336
rect 20314 12280 20319 12336
rect 20180 12278 20319 12280
rect 20180 12276 20186 12278
rect 20253 12275 20319 12278
rect 22001 12338 22067 12341
rect 23565 12338 23631 12341
rect 22001 12336 23631 12338
rect 22001 12280 22006 12336
rect 22062 12280 23570 12336
rect 23626 12280 23631 12336
rect 22001 12278 23631 12280
rect 22001 12275 22067 12278
rect 23565 12275 23631 12278
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 24761 11930 24827 11933
rect 27520 11930 28000 11960
rect 24761 11928 28000 11930
rect 24761 11872 24766 11928
rect 24822 11872 28000 11928
rect 24761 11870 28000 11872
rect 24761 11867 24827 11870
rect 27520 11840 28000 11870
rect 12065 11794 12131 11797
rect 17585 11794 17651 11797
rect 12065 11792 17651 11794
rect 12065 11736 12070 11792
rect 12126 11736 17590 11792
rect 17646 11736 17651 11792
rect 12065 11734 17651 11736
rect 12065 11731 12131 11734
rect 17585 11731 17651 11734
rect 4981 11658 5047 11661
rect 12341 11658 12407 11661
rect 4981 11656 12407 11658
rect 4981 11600 4986 11656
rect 5042 11600 12346 11656
rect 12402 11600 12407 11656
rect 4981 11598 12407 11600
rect 4981 11595 5047 11598
rect 12341 11595 12407 11598
rect 20069 11522 20135 11525
rect 22829 11522 22895 11525
rect 20069 11520 22895 11522
rect 20069 11464 20074 11520
rect 20130 11464 22834 11520
rect 22890 11464 22895 11520
rect 20069 11462 22895 11464
rect 20069 11459 20135 11462
rect 22829 11459 22895 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 15469 11386 15535 11389
rect 18229 11386 18295 11389
rect 15469 11384 18295 11386
rect 15469 11328 15474 11384
rect 15530 11328 18234 11384
rect 18290 11328 18295 11384
rect 15469 11326 18295 11328
rect 15469 11323 15535 11326
rect 18229 11323 18295 11326
rect 21909 11386 21975 11389
rect 25221 11386 25287 11389
rect 27520 11386 28000 11416
rect 21909 11384 28000 11386
rect 21909 11328 21914 11384
rect 21970 11328 25226 11384
rect 25282 11328 28000 11384
rect 21909 11326 28000 11328
rect 21909 11323 21975 11326
rect 25221 11323 25287 11326
rect 27520 11296 28000 11326
rect 12525 11114 12591 11117
rect 18045 11114 18111 11117
rect 12525 11112 18111 11114
rect 12525 11056 12530 11112
rect 12586 11056 18050 11112
rect 18106 11056 18111 11112
rect 12525 11054 18111 11056
rect 12525 11051 12591 11054
rect 18045 11051 18111 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 17769 10842 17835 10845
rect 20437 10842 20503 10845
rect 27520 10842 28000 10872
rect 17769 10840 20503 10842
rect 17769 10784 17774 10840
rect 17830 10784 20442 10840
rect 20498 10784 20503 10840
rect 17769 10782 20503 10784
rect 17769 10779 17835 10782
rect 20437 10779 20503 10782
rect 24902 10782 28000 10842
rect 10869 10706 10935 10709
rect 12433 10706 12499 10709
rect 18413 10706 18479 10709
rect 10869 10704 18479 10706
rect 10869 10648 10874 10704
rect 10930 10648 12438 10704
rect 12494 10648 18418 10704
rect 18474 10648 18479 10704
rect 10869 10646 18479 10648
rect 10869 10643 10935 10646
rect 12433 10643 12499 10646
rect 18413 10643 18479 10646
rect 19241 10706 19307 10709
rect 24902 10706 24962 10782
rect 27520 10752 28000 10782
rect 19241 10704 24962 10706
rect 19241 10648 19246 10704
rect 19302 10648 24962 10704
rect 19241 10646 24962 10648
rect 19241 10643 19307 10646
rect 13629 10570 13695 10573
rect 15469 10570 15535 10573
rect 13629 10568 15535 10570
rect 13629 10512 13634 10568
rect 13690 10512 15474 10568
rect 15530 10512 15535 10568
rect 13629 10510 15535 10512
rect 13629 10507 13695 10510
rect 15469 10507 15535 10510
rect 15837 10570 15903 10573
rect 18781 10570 18847 10573
rect 20805 10570 20871 10573
rect 15837 10568 20871 10570
rect 15837 10512 15842 10568
rect 15898 10512 18786 10568
rect 18842 10512 20810 10568
rect 20866 10512 20871 10568
rect 15837 10510 20871 10512
rect 15837 10507 15903 10510
rect 18781 10507 18847 10510
rect 20805 10507 20871 10510
rect 14549 10434 14615 10437
rect 17493 10434 17559 10437
rect 14549 10432 17559 10434
rect 14549 10376 14554 10432
rect 14610 10376 17498 10432
rect 17554 10376 17559 10432
rect 14549 10374 17559 10376
rect 14549 10371 14615 10374
rect 17493 10371 17559 10374
rect 21909 10434 21975 10437
rect 23841 10434 23907 10437
rect 21909 10432 23907 10434
rect 21909 10376 21914 10432
rect 21970 10376 23846 10432
rect 23902 10376 23907 10432
rect 21909 10374 23907 10376
rect 21909 10371 21975 10374
rect 23841 10371 23907 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 20069 10298 20135 10301
rect 25589 10298 25655 10301
rect 20069 10296 25655 10298
rect 20069 10240 20074 10296
rect 20130 10240 25594 10296
rect 25650 10240 25655 10296
rect 20069 10238 25655 10240
rect 20069 10235 20135 10238
rect 25589 10235 25655 10238
rect 4337 10162 4403 10165
rect 13537 10162 13603 10165
rect 14457 10164 14523 10165
rect 14406 10162 14412 10164
rect 4337 10160 13603 10162
rect 4337 10104 4342 10160
rect 4398 10104 13542 10160
rect 13598 10104 13603 10160
rect 4337 10102 13603 10104
rect 14366 10102 14412 10162
rect 14476 10160 14523 10164
rect 14518 10104 14523 10160
rect 4337 10099 4403 10102
rect 13537 10099 13603 10102
rect 14406 10100 14412 10102
rect 14476 10100 14523 10104
rect 14457 10099 14523 10100
rect 16757 10162 16823 10165
rect 27520 10162 28000 10192
rect 16757 10160 28000 10162
rect 16757 10104 16762 10160
rect 16818 10104 28000 10160
rect 16757 10102 28000 10104
rect 16757 10099 16823 10102
rect 27520 10072 28000 10102
rect 13629 10026 13695 10029
rect 17953 10026 18019 10029
rect 13629 10024 18019 10026
rect 13629 9968 13634 10024
rect 13690 9968 17958 10024
rect 18014 9968 18019 10024
rect 13629 9966 18019 9968
rect 13629 9963 13695 9966
rect 17953 9963 18019 9966
rect 15561 9890 15627 9893
rect 23565 9890 23631 9893
rect 15561 9888 23631 9890
rect 15561 9832 15566 9888
rect 15622 9832 23570 9888
rect 23626 9832 23631 9888
rect 15561 9830 23631 9832
rect 15561 9827 15627 9830
rect 23565 9827 23631 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 1485 9754 1551 9757
rect 2865 9754 2931 9757
rect 1485 9752 2931 9754
rect 1485 9696 1490 9752
rect 1546 9696 2870 9752
rect 2926 9696 2931 9752
rect 1485 9694 2931 9696
rect 1485 9691 1551 9694
rect 2865 9691 2931 9694
rect 18689 9754 18755 9757
rect 21541 9754 21607 9757
rect 18689 9752 21607 9754
rect 18689 9696 18694 9752
rect 18750 9696 21546 9752
rect 21602 9696 21607 9752
rect 18689 9694 21607 9696
rect 18689 9691 18755 9694
rect 21541 9691 21607 9694
rect 2773 9618 2839 9621
rect 10133 9618 10199 9621
rect 2773 9616 10199 9618
rect 2773 9560 2778 9616
rect 2834 9560 10138 9616
rect 10194 9560 10199 9616
rect 2773 9558 10199 9560
rect 2773 9555 2839 9558
rect 10133 9555 10199 9558
rect 10961 9618 11027 9621
rect 13905 9618 13971 9621
rect 10961 9616 13971 9618
rect 10961 9560 10966 9616
rect 11022 9560 13910 9616
rect 13966 9560 13971 9616
rect 10961 9558 13971 9560
rect 10961 9555 11027 9558
rect 13905 9555 13971 9558
rect 18505 9618 18571 9621
rect 27520 9618 28000 9648
rect 18505 9616 28000 9618
rect 18505 9560 18510 9616
rect 18566 9560 28000 9616
rect 18505 9558 28000 9560
rect 18505 9555 18571 9558
rect 27520 9528 28000 9558
rect 21081 9482 21147 9485
rect 23841 9482 23907 9485
rect 21081 9480 23907 9482
rect 21081 9424 21086 9480
rect 21142 9424 23846 9480
rect 23902 9424 23907 9480
rect 21081 9422 23907 9424
rect 21081 9419 21147 9422
rect 23841 9419 23907 9422
rect 2865 9346 2931 9349
rect 9673 9346 9739 9349
rect 2865 9344 9739 9346
rect 2865 9288 2870 9344
rect 2926 9288 9678 9344
rect 9734 9288 9739 9344
rect 2865 9286 9739 9288
rect 2865 9283 2931 9286
rect 9673 9283 9739 9286
rect 13905 9346 13971 9349
rect 17769 9346 17835 9349
rect 13905 9344 17835 9346
rect 13905 9288 13910 9344
rect 13966 9288 17774 9344
rect 17830 9288 17835 9344
rect 13905 9286 17835 9288
rect 13905 9283 13971 9286
rect 17769 9283 17835 9286
rect 21173 9346 21239 9349
rect 23749 9346 23815 9349
rect 21173 9344 23815 9346
rect 21173 9288 21178 9344
rect 21234 9288 23754 9344
rect 23810 9288 23815 9344
rect 21173 9286 23815 9288
rect 21173 9283 21239 9286
rect 23749 9283 23815 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 12709 9074 12775 9077
rect 19333 9074 19399 9077
rect 20989 9074 21055 9077
rect 12709 9072 21055 9074
rect 12709 9016 12714 9072
rect 12770 9016 19338 9072
rect 19394 9016 20994 9072
rect 21050 9016 21055 9072
rect 12709 9014 21055 9016
rect 12709 9011 12775 9014
rect 19333 9011 19399 9014
rect 20989 9011 21055 9014
rect 21173 9074 21239 9077
rect 24669 9074 24735 9077
rect 27520 9074 28000 9104
rect 21173 9072 24735 9074
rect 21173 9016 21178 9072
rect 21234 9016 24674 9072
rect 24730 9016 24735 9072
rect 21173 9014 24735 9016
rect 21173 9011 21239 9014
rect 24669 9011 24735 9014
rect 24902 9014 28000 9074
rect 9121 8938 9187 8941
rect 12249 8938 12315 8941
rect 9121 8936 12315 8938
rect 9121 8880 9126 8936
rect 9182 8880 12254 8936
rect 12310 8880 12315 8936
rect 9121 8878 12315 8880
rect 9121 8875 9187 8878
rect 12249 8875 12315 8878
rect 13629 8938 13695 8941
rect 17033 8938 17099 8941
rect 13629 8936 17099 8938
rect 13629 8880 13634 8936
rect 13690 8880 17038 8936
rect 17094 8880 17099 8936
rect 13629 8878 17099 8880
rect 13629 8875 13695 8878
rect 17033 8875 17099 8878
rect 24761 8938 24827 8941
rect 24902 8938 24962 9014
rect 27520 8984 28000 9014
rect 24761 8936 24962 8938
rect 24761 8880 24766 8936
rect 24822 8880 24962 8936
rect 24761 8878 24962 8880
rect 24761 8875 24827 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 18229 8666 18295 8669
rect 20069 8666 20135 8669
rect 18229 8664 20135 8666
rect 18229 8608 18234 8664
rect 18290 8608 20074 8664
rect 20130 8608 20135 8664
rect 18229 8606 20135 8608
rect 18229 8603 18295 8606
rect 20069 8603 20135 8606
rect 11053 8530 11119 8533
rect 21725 8530 21791 8533
rect 11053 8528 21791 8530
rect 11053 8472 11058 8528
rect 11114 8472 21730 8528
rect 21786 8472 21791 8528
rect 11053 8470 21791 8472
rect 11053 8467 11119 8470
rect 21725 8467 21791 8470
rect 24669 8530 24735 8533
rect 27520 8530 28000 8560
rect 24669 8528 28000 8530
rect 24669 8472 24674 8528
rect 24730 8472 28000 8528
rect 24669 8470 28000 8472
rect 24669 8467 24735 8470
rect 27520 8440 28000 8470
rect 18413 8394 18479 8397
rect 12344 8392 18479 8394
rect 12344 8336 18418 8392
rect 18474 8336 18479 8392
rect 12344 8334 18479 8336
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 12344 8122 12404 8334
rect 18413 8331 18479 8334
rect 20069 8394 20135 8397
rect 22553 8394 22619 8397
rect 20069 8392 22619 8394
rect 20069 8336 20074 8392
rect 20130 8336 22558 8392
rect 22614 8336 22619 8392
rect 20069 8334 22619 8336
rect 20069 8331 20135 8334
rect 22553 8331 22619 8334
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 10734 8062 12404 8122
rect 3693 7986 3759 7989
rect 10734 7986 10794 8062
rect 3693 7984 10794 7986
rect 3693 7928 3698 7984
rect 3754 7928 10794 7984
rect 3693 7926 10794 7928
rect 12525 7986 12591 7989
rect 15561 7986 15627 7989
rect 12525 7984 15627 7986
rect 12525 7928 12530 7984
rect 12586 7928 15566 7984
rect 15622 7928 15627 7984
rect 12525 7926 15627 7928
rect 3693 7923 3759 7926
rect 12525 7923 12591 7926
rect 15561 7923 15627 7926
rect 18505 7986 18571 7989
rect 24761 7986 24827 7989
rect 18505 7984 24827 7986
rect 18505 7928 18510 7984
rect 18566 7928 24766 7984
rect 24822 7928 24827 7984
rect 18505 7926 24827 7928
rect 18505 7923 18571 7926
rect 20164 7853 20224 7926
rect 24761 7923 24827 7926
rect 19517 7850 19583 7853
rect 14782 7848 19583 7850
rect 14782 7792 19522 7848
rect 19578 7792 19583 7848
rect 14782 7790 19583 7792
rect 12249 7714 12315 7717
rect 14782 7714 14842 7790
rect 19517 7787 19583 7790
rect 20161 7848 20227 7853
rect 20161 7792 20166 7848
rect 20222 7792 20227 7848
rect 20161 7787 20227 7792
rect 24117 7850 24183 7853
rect 27520 7850 28000 7880
rect 24117 7848 28000 7850
rect 24117 7792 24122 7848
rect 24178 7792 28000 7848
rect 24117 7790 28000 7792
rect 24117 7787 24183 7790
rect 27520 7760 28000 7790
rect 12249 7712 14842 7714
rect 12249 7656 12254 7712
rect 12310 7656 14842 7712
rect 12249 7654 14842 7656
rect 12249 7651 12315 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 6913 7578 6979 7581
rect 12433 7578 12499 7581
rect 6913 7576 12499 7578
rect 6913 7520 6918 7576
rect 6974 7520 12438 7576
rect 12494 7520 12499 7576
rect 6913 7518 12499 7520
rect 6913 7515 6979 7518
rect 12433 7515 12499 7518
rect 17309 7306 17375 7309
rect 23841 7306 23907 7309
rect 27520 7306 28000 7336
rect 17309 7304 20178 7306
rect 17309 7248 17314 7304
rect 17370 7248 20178 7304
rect 17309 7246 20178 7248
rect 17309 7243 17375 7246
rect 20118 7170 20178 7246
rect 23841 7304 28000 7306
rect 23841 7248 23846 7304
rect 23902 7248 28000 7304
rect 23841 7246 28000 7248
rect 23841 7243 23907 7246
rect 27520 7216 28000 7246
rect 21265 7170 21331 7173
rect 22093 7170 22159 7173
rect 20118 7168 22159 7170
rect 20118 7112 21270 7168
rect 21326 7112 22098 7168
rect 22154 7112 22159 7168
rect 20118 7110 22159 7112
rect 21265 7107 21331 7110
rect 22093 7107 22159 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 22001 6898 22067 6901
rect 25221 6898 25287 6901
rect 22001 6896 25287 6898
rect 22001 6840 22006 6896
rect 22062 6840 25226 6896
rect 25282 6840 25287 6896
rect 22001 6838 25287 6840
rect 22001 6835 22067 6838
rect 25221 6835 25287 6838
rect 13537 6762 13603 6765
rect 15285 6762 15351 6765
rect 13537 6760 15351 6762
rect 13537 6704 13542 6760
rect 13598 6704 15290 6760
rect 15346 6704 15351 6760
rect 13537 6702 15351 6704
rect 13537 6699 13603 6702
rect 15285 6699 15351 6702
rect 18873 6762 18939 6765
rect 27520 6762 28000 6792
rect 18873 6760 28000 6762
rect 18873 6704 18878 6760
rect 18934 6704 28000 6760
rect 18873 6702 28000 6704
rect 18873 6699 18939 6702
rect 27520 6672 28000 6702
rect 12249 6626 12315 6629
rect 14181 6626 14247 6629
rect 12249 6624 14247 6626
rect 12249 6568 12254 6624
rect 12310 6568 14186 6624
rect 14242 6568 14247 6624
rect 12249 6566 14247 6568
rect 12249 6563 12315 6566
rect 14181 6563 14247 6566
rect 16481 6626 16547 6629
rect 16941 6626 17007 6629
rect 17769 6626 17835 6629
rect 16481 6624 17835 6626
rect 16481 6568 16486 6624
rect 16542 6568 16946 6624
rect 17002 6568 17774 6624
rect 17830 6568 17835 6624
rect 16481 6566 17835 6568
rect 16481 6563 16547 6566
rect 16941 6563 17007 6566
rect 17769 6563 17835 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 22185 6490 22251 6493
rect 16070 6488 22251 6490
rect 16070 6432 22190 6488
rect 22246 6432 22251 6488
rect 16070 6430 22251 6432
rect 2313 6354 2379 6357
rect 12893 6354 12959 6357
rect 2313 6352 12959 6354
rect 2313 6296 2318 6352
rect 2374 6296 12898 6352
rect 12954 6296 12959 6352
rect 2313 6294 12959 6296
rect 2313 6291 2379 6294
rect 12893 6291 12959 6294
rect 14457 6354 14523 6357
rect 16070 6354 16130 6430
rect 22185 6427 22251 6430
rect 14457 6352 16130 6354
rect 14457 6296 14462 6352
rect 14518 6296 16130 6352
rect 14457 6294 16130 6296
rect 16205 6354 16271 6357
rect 21081 6354 21147 6357
rect 16205 6352 21147 6354
rect 16205 6296 16210 6352
rect 16266 6296 21086 6352
rect 21142 6296 21147 6352
rect 16205 6294 21147 6296
rect 14457 6291 14523 6294
rect 16205 6291 16271 6294
rect 21081 6291 21147 6294
rect 19149 6218 19215 6221
rect 21357 6218 21423 6221
rect 19149 6216 21423 6218
rect 19149 6160 19154 6216
rect 19210 6160 21362 6216
rect 21418 6160 21423 6216
rect 19149 6158 21423 6160
rect 19149 6155 19215 6158
rect 21357 6155 21423 6158
rect 21541 6082 21607 6085
rect 24669 6082 24735 6085
rect 27520 6082 28000 6112
rect 21541 6080 24735 6082
rect 21541 6024 21546 6080
rect 21602 6024 24674 6080
rect 24730 6024 24735 6080
rect 21541 6022 24735 6024
rect 21541 6019 21607 6022
rect 24669 6019 24735 6022
rect 24902 6022 28000 6082
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 13445 5810 13511 5813
rect 17585 5810 17651 5813
rect 13445 5808 17651 5810
rect 13445 5752 13450 5808
rect 13506 5752 17590 5808
rect 17646 5752 17651 5808
rect 13445 5750 17651 5752
rect 13445 5747 13511 5750
rect 17585 5747 17651 5750
rect 19057 5810 19123 5813
rect 20897 5810 20963 5813
rect 19057 5808 20963 5810
rect 19057 5752 19062 5808
rect 19118 5752 20902 5808
rect 20958 5752 20963 5808
rect 19057 5750 20963 5752
rect 19057 5747 19123 5750
rect 20897 5747 20963 5750
rect 21081 5810 21147 5813
rect 24902 5810 24962 6022
rect 27520 5992 28000 6022
rect 21081 5808 24962 5810
rect 21081 5752 21086 5808
rect 21142 5752 24962 5808
rect 21081 5750 24962 5752
rect 21081 5747 21147 5750
rect 11881 5674 11947 5677
rect 21265 5674 21331 5677
rect 11881 5672 21331 5674
rect 11881 5616 11886 5672
rect 11942 5616 21270 5672
rect 21326 5616 21331 5672
rect 11881 5614 21331 5616
rect 11881 5611 11947 5614
rect 21265 5611 21331 5614
rect 27520 5538 28000 5568
rect 24764 5478 28000 5538
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 14089 5266 14155 5269
rect 16849 5266 16915 5269
rect 14089 5264 16915 5266
rect 14089 5208 14094 5264
rect 14150 5208 16854 5264
rect 16910 5208 16915 5264
rect 14089 5206 16915 5208
rect 14089 5203 14155 5206
rect 16849 5203 16915 5206
rect 18873 5266 18939 5269
rect 20345 5266 20411 5269
rect 21633 5266 21699 5269
rect 18873 5264 21699 5266
rect 18873 5208 18878 5264
rect 18934 5208 20350 5264
rect 20406 5208 21638 5264
rect 21694 5208 21699 5264
rect 18873 5206 21699 5208
rect 18873 5203 18939 5206
rect 20345 5203 20411 5206
rect 21633 5203 21699 5206
rect 2957 5130 3023 5133
rect 22737 5130 22803 5133
rect 24764 5130 24824 5478
rect 27520 5448 28000 5478
rect 2957 5128 22803 5130
rect 2957 5072 2962 5128
rect 3018 5072 22742 5128
rect 22798 5072 22803 5128
rect 2957 5070 22803 5072
rect 2957 5067 3023 5070
rect 22737 5067 22803 5070
rect 23798 5070 24824 5130
rect 10777 4994 10843 4997
rect 10777 4992 17050 4994
rect 10777 4936 10782 4992
rect 10838 4936 17050 4992
rect 10777 4934 17050 4936
rect 10777 4931 10843 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 14641 4858 14707 4861
rect 16757 4858 16823 4861
rect 14641 4856 16823 4858
rect 14641 4800 14646 4856
rect 14702 4800 16762 4856
rect 16818 4800 16823 4856
rect 14641 4798 16823 4800
rect 14641 4795 14707 4798
rect 16757 4795 16823 4798
rect 0 4722 480 4752
rect 2865 4722 2931 4725
rect 0 4720 2931 4722
rect 0 4664 2870 4720
rect 2926 4664 2931 4720
rect 0 4662 2931 4664
rect 0 4632 480 4662
rect 2865 4659 2931 4662
rect 8293 4722 8359 4725
rect 16021 4722 16087 4725
rect 8293 4720 16087 4722
rect 8293 4664 8298 4720
rect 8354 4664 16026 4720
rect 16082 4664 16087 4720
rect 8293 4662 16087 4664
rect 16990 4722 17050 4934
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 20069 4858 20135 4861
rect 23798 4858 23858 5070
rect 27520 4994 28000 5024
rect 20069 4856 23858 4858
rect 20069 4800 20074 4856
rect 20130 4800 23858 4856
rect 20069 4798 23858 4800
rect 23982 4934 28000 4994
rect 20069 4795 20135 4798
rect 20897 4722 20963 4725
rect 16990 4720 20963 4722
rect 16990 4664 20902 4720
rect 20958 4664 20963 4720
rect 16990 4662 20963 4664
rect 8293 4659 8359 4662
rect 16021 4659 16087 4662
rect 20897 4659 20963 4662
rect 22001 4722 22067 4725
rect 23841 4722 23907 4725
rect 22001 4720 23907 4722
rect 22001 4664 22006 4720
rect 22062 4664 23846 4720
rect 23902 4664 23907 4720
rect 22001 4662 23907 4664
rect 22001 4659 22067 4662
rect 23841 4659 23907 4662
rect 9765 4586 9831 4589
rect 14641 4586 14707 4589
rect 9765 4584 14707 4586
rect 9765 4528 9770 4584
rect 9826 4528 14646 4584
rect 14702 4528 14707 4584
rect 9765 4526 14707 4528
rect 9765 4523 9831 4526
rect 14641 4523 14707 4526
rect 18597 4586 18663 4589
rect 20897 4586 20963 4589
rect 18597 4584 20963 4586
rect 18597 4528 18602 4584
rect 18658 4528 20902 4584
rect 20958 4528 20963 4584
rect 18597 4526 20963 4528
rect 18597 4523 18663 4526
rect 20897 4523 20963 4526
rect 18689 4450 18755 4453
rect 21173 4450 21239 4453
rect 23982 4450 24042 4934
rect 27520 4904 28000 4934
rect 18689 4448 24042 4450
rect 18689 4392 18694 4448
rect 18750 4392 21178 4448
rect 21234 4392 24042 4448
rect 18689 4390 24042 4392
rect 24945 4450 25011 4453
rect 27520 4450 28000 4480
rect 24945 4448 28000 4450
rect 24945 4392 24950 4448
rect 25006 4392 28000 4448
rect 24945 4390 28000 4392
rect 18689 4387 18755 4390
rect 21173 4387 21239 4390
rect 24945 4387 25011 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 17033 4314 17099 4317
rect 19333 4314 19399 4317
rect 17033 4312 19399 4314
rect 17033 4256 17038 4312
rect 17094 4256 19338 4312
rect 19394 4256 19399 4312
rect 17033 4254 19399 4256
rect 17033 4251 17099 4254
rect 19333 4251 19399 4254
rect 10685 4178 10751 4181
rect 15377 4178 15443 4181
rect 10685 4176 15443 4178
rect 10685 4120 10690 4176
rect 10746 4120 15382 4176
rect 15438 4120 15443 4176
rect 10685 4118 15443 4120
rect 10685 4115 10751 4118
rect 15377 4115 15443 4118
rect 16021 4178 16087 4181
rect 18689 4178 18755 4181
rect 16021 4176 18755 4178
rect 16021 4120 16026 4176
rect 16082 4120 18694 4176
rect 18750 4120 18755 4176
rect 16021 4118 18755 4120
rect 16021 4115 16087 4118
rect 18689 4115 18755 4118
rect 22553 4178 22619 4181
rect 25405 4178 25471 4181
rect 22553 4176 25471 4178
rect 22553 4120 22558 4176
rect 22614 4120 25410 4176
rect 25466 4120 25471 4176
rect 22553 4118 25471 4120
rect 22553 4115 22619 4118
rect 25405 4115 25471 4118
rect 7097 4042 7163 4045
rect 11053 4042 11119 4045
rect 7097 4040 11119 4042
rect 7097 3984 7102 4040
rect 7158 3984 11058 4040
rect 11114 3984 11119 4040
rect 7097 3982 11119 3984
rect 7097 3979 7163 3982
rect 11053 3979 11119 3982
rect 14733 4042 14799 4045
rect 16573 4042 16639 4045
rect 14733 4040 16639 4042
rect 14733 3984 14738 4040
rect 14794 3984 16578 4040
rect 16634 3984 16639 4040
rect 14733 3982 16639 3984
rect 14733 3979 14799 3982
rect 16573 3979 16639 3982
rect 19149 4042 19215 4045
rect 24025 4042 24091 4045
rect 19149 4040 24091 4042
rect 19149 3984 19154 4040
rect 19210 3984 24030 4040
rect 24086 3984 24091 4040
rect 19149 3982 24091 3984
rect 19149 3979 19215 3982
rect 24025 3979 24091 3982
rect 23657 3906 23723 3909
rect 23657 3904 24410 3906
rect 23657 3848 23662 3904
rect 23718 3848 24410 3904
rect 23657 3846 24410 3848
rect 23657 3843 23723 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 12709 3770 12775 3773
rect 16573 3770 16639 3773
rect 12709 3768 16639 3770
rect 12709 3712 12714 3768
rect 12770 3712 16578 3768
rect 16634 3712 16639 3768
rect 12709 3710 16639 3712
rect 12709 3707 12775 3710
rect 16573 3707 16639 3710
rect 22369 3770 22435 3773
rect 24117 3770 24183 3773
rect 22369 3768 24183 3770
rect 22369 3712 22374 3768
rect 22430 3712 24122 3768
rect 24178 3712 24183 3768
rect 22369 3710 24183 3712
rect 24350 3770 24410 3846
rect 27520 3770 28000 3800
rect 24350 3710 28000 3770
rect 22369 3707 22435 3710
rect 24117 3707 24183 3710
rect 27520 3680 28000 3710
rect 12433 3634 12499 3637
rect 16113 3634 16179 3637
rect 22737 3634 22803 3637
rect 12433 3632 16179 3634
rect 12433 3576 12438 3632
rect 12494 3576 16118 3632
rect 16174 3576 16179 3632
rect 12433 3574 16179 3576
rect 12433 3571 12499 3574
rect 16113 3571 16179 3574
rect 19198 3632 22803 3634
rect 19198 3576 22742 3632
rect 22798 3576 22803 3632
rect 19198 3574 22803 3576
rect 19198 3501 19258 3574
rect 22737 3571 22803 3574
rect 23749 3634 23815 3637
rect 23749 3632 24824 3634
rect 23749 3576 23754 3632
rect 23810 3576 24824 3632
rect 23749 3574 24824 3576
rect 23749 3571 23815 3574
rect 933 3498 999 3501
rect 1945 3498 2011 3501
rect 933 3496 2011 3498
rect 933 3440 938 3496
rect 994 3440 1950 3496
rect 2006 3440 2011 3496
rect 933 3438 2011 3440
rect 933 3435 999 3438
rect 1945 3435 2011 3438
rect 13629 3498 13695 3501
rect 19149 3498 19258 3501
rect 23933 3498 23999 3501
rect 13629 3496 19258 3498
rect 13629 3440 13634 3496
rect 13690 3440 19154 3496
rect 19210 3440 19258 3496
rect 13629 3438 19258 3440
rect 19382 3496 23999 3498
rect 19382 3440 23938 3496
rect 23994 3440 23999 3496
rect 19382 3438 23999 3440
rect 13629 3435 13695 3438
rect 19149 3435 19215 3438
rect 15377 3362 15443 3365
rect 19382 3362 19442 3438
rect 23933 3435 23999 3438
rect 15377 3360 19442 3362
rect 15377 3304 15382 3360
rect 15438 3304 19442 3360
rect 15377 3302 19442 3304
rect 19517 3362 19583 3365
rect 23749 3362 23815 3365
rect 19517 3360 23815 3362
rect 19517 3304 19522 3360
rect 19578 3304 23754 3360
rect 23810 3304 23815 3360
rect 19517 3302 23815 3304
rect 15377 3299 15443 3302
rect 19517 3299 19583 3302
rect 23749 3299 23815 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 10133 3226 10199 3229
rect 14733 3226 14799 3229
rect 10133 3224 14799 3226
rect 10133 3168 10138 3224
rect 10194 3168 14738 3224
rect 14794 3168 14799 3224
rect 10133 3166 14799 3168
rect 10133 3163 10199 3166
rect 14733 3163 14799 3166
rect 15469 3226 15535 3229
rect 20437 3226 20503 3229
rect 15469 3224 20503 3226
rect 15469 3168 15474 3224
rect 15530 3168 20442 3224
rect 20498 3168 20503 3224
rect 15469 3166 20503 3168
rect 15469 3163 15535 3166
rect 20437 3163 20503 3166
rect 21449 3226 21515 3229
rect 23565 3226 23631 3229
rect 21449 3224 23631 3226
rect 21449 3168 21454 3224
rect 21510 3168 23570 3224
rect 23626 3168 23631 3224
rect 21449 3166 23631 3168
rect 24764 3226 24824 3574
rect 27520 3226 28000 3256
rect 24764 3166 28000 3226
rect 21449 3163 21515 3166
rect 23565 3163 23631 3166
rect 27520 3136 28000 3166
rect 11421 3090 11487 3093
rect 15929 3090 15995 3093
rect 11421 3088 15995 3090
rect 11421 3032 11426 3088
rect 11482 3032 15934 3088
rect 15990 3032 15995 3088
rect 11421 3030 15995 3032
rect 11421 3027 11487 3030
rect 15929 3027 15995 3030
rect 20253 3090 20319 3093
rect 22737 3090 22803 3093
rect 20253 3088 22803 3090
rect 20253 3032 20258 3088
rect 20314 3032 22742 3088
rect 22798 3032 22803 3088
rect 20253 3030 22803 3032
rect 20253 3027 20319 3030
rect 22737 3027 22803 3030
rect 13629 2954 13695 2957
rect 17953 2954 18019 2957
rect 19517 2954 19583 2957
rect 13629 2952 18019 2954
rect 13629 2896 13634 2952
rect 13690 2896 17958 2952
rect 18014 2896 18019 2952
rect 13629 2894 18019 2896
rect 13629 2891 13695 2894
rect 17953 2891 18019 2894
rect 19382 2952 19583 2954
rect 19382 2896 19522 2952
rect 19578 2896 19583 2952
rect 19382 2894 19583 2896
rect 11605 2818 11671 2821
rect 14549 2818 14615 2821
rect 11605 2816 14615 2818
rect 11605 2760 11610 2816
rect 11666 2760 14554 2816
rect 14610 2760 14615 2816
rect 11605 2758 14615 2760
rect 11605 2755 11671 2758
rect 14549 2755 14615 2758
rect 15745 2818 15811 2821
rect 19382 2818 19442 2894
rect 19517 2891 19583 2894
rect 24761 2954 24827 2957
rect 27521 2954 27587 2957
rect 24761 2952 27587 2954
rect 24761 2896 24766 2952
rect 24822 2896 27526 2952
rect 27582 2896 27587 2952
rect 24761 2894 27587 2896
rect 24761 2891 24827 2894
rect 27521 2891 27587 2894
rect 15745 2816 19442 2818
rect 15745 2760 15750 2816
rect 15806 2760 19442 2816
rect 15745 2758 19442 2760
rect 22645 2818 22711 2821
rect 25497 2818 25563 2821
rect 22645 2816 25563 2818
rect 22645 2760 22650 2816
rect 22706 2760 25502 2816
rect 25558 2760 25563 2816
rect 22645 2758 25563 2760
rect 15745 2755 15811 2758
rect 22645 2755 22711 2758
rect 25497 2755 25563 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 13077 2682 13143 2685
rect 16113 2682 16179 2685
rect 18873 2682 18939 2685
rect 27520 2682 28000 2712
rect 13077 2680 18939 2682
rect 13077 2624 13082 2680
rect 13138 2624 16118 2680
rect 16174 2624 18878 2680
rect 18934 2624 18939 2680
rect 13077 2622 18939 2624
rect 13077 2619 13143 2622
rect 16113 2619 16179 2622
rect 18873 2619 18939 2622
rect 26742 2622 28000 2682
rect 5717 2546 5783 2549
rect 11697 2546 11763 2549
rect 5717 2544 11763 2546
rect 5717 2488 5722 2544
rect 5778 2488 11702 2544
rect 11758 2488 11763 2544
rect 5717 2486 11763 2488
rect 5717 2483 5783 2486
rect 11697 2483 11763 2486
rect 14825 2546 14891 2549
rect 18045 2546 18111 2549
rect 14825 2544 18111 2546
rect 14825 2488 14830 2544
rect 14886 2488 18050 2544
rect 18106 2488 18111 2544
rect 14825 2486 18111 2488
rect 14825 2483 14891 2486
rect 18045 2483 18111 2486
rect 18781 2546 18847 2549
rect 26742 2546 26802 2622
rect 27520 2592 28000 2622
rect 18781 2544 26802 2546
rect 18781 2488 18786 2544
rect 18842 2488 26802 2544
rect 18781 2486 26802 2488
rect 18781 2483 18847 2486
rect 14457 2410 14523 2413
rect 22093 2410 22159 2413
rect 14457 2408 22159 2410
rect 14457 2352 14462 2408
rect 14518 2352 22098 2408
rect 22154 2352 22159 2408
rect 14457 2350 22159 2352
rect 14457 2347 14523 2350
rect 22093 2347 22159 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 16941 2138 17007 2141
rect 22829 2138 22895 2141
rect 16941 2136 22895 2138
rect 16941 2080 16946 2136
rect 17002 2080 22834 2136
rect 22890 2080 22895 2136
rect 16941 2078 22895 2080
rect 16941 2075 17007 2078
rect 22829 2075 22895 2078
rect 13353 2002 13419 2005
rect 20713 2002 20779 2005
rect 27520 2002 28000 2032
rect 13353 2000 20779 2002
rect 13353 1944 13358 2000
rect 13414 1944 20718 2000
rect 20774 1944 20779 2000
rect 13353 1942 20779 1944
rect 13353 1939 13419 1942
rect 20713 1939 20779 1942
rect 26926 1942 28000 2002
rect 289 1730 355 1733
rect 12617 1730 12683 1733
rect 26926 1730 26986 1942
rect 27520 1912 28000 1942
rect 289 1728 12683 1730
rect 289 1672 294 1728
rect 350 1672 12622 1728
rect 12678 1672 12683 1728
rect 289 1670 12683 1672
rect 289 1667 355 1670
rect 12617 1667 12683 1670
rect 21406 1670 26986 1730
rect 11605 1594 11671 1597
rect 17309 1594 17375 1597
rect 11605 1592 17375 1594
rect 11605 1536 11610 1592
rect 11666 1536 17314 1592
rect 17370 1536 17375 1592
rect 11605 1534 17375 1536
rect 11605 1531 11671 1534
rect 17309 1531 17375 1534
rect 10961 1458 11027 1461
rect 15285 1458 15351 1461
rect 10961 1456 15351 1458
rect 10961 1400 10966 1456
rect 11022 1400 15290 1456
rect 15346 1400 15351 1456
rect 10961 1398 15351 1400
rect 10961 1395 11027 1398
rect 15285 1395 15351 1398
rect 15837 1458 15903 1461
rect 21406 1458 21466 1670
rect 24025 1594 24091 1597
rect 24025 1592 26986 1594
rect 24025 1536 24030 1592
rect 24086 1536 26986 1592
rect 24025 1534 26986 1536
rect 24025 1531 24091 1534
rect 15837 1456 21466 1458
rect 15837 1400 15842 1456
rect 15898 1400 21466 1456
rect 15837 1398 21466 1400
rect 21909 1458 21975 1461
rect 26785 1458 26851 1461
rect 21909 1456 26851 1458
rect 21909 1400 21914 1456
rect 21970 1400 26790 1456
rect 26846 1400 26851 1456
rect 21909 1398 26851 1400
rect 26926 1458 26986 1534
rect 27520 1458 28000 1488
rect 26926 1398 28000 1458
rect 15837 1395 15903 1398
rect 21909 1395 21975 1398
rect 26785 1395 26851 1398
rect 27520 1368 28000 1398
rect 24577 1322 24643 1325
rect 24761 1322 24827 1325
rect 24577 1320 24827 1322
rect 24577 1264 24582 1320
rect 24638 1264 24766 1320
rect 24822 1264 24827 1320
rect 24577 1262 24827 1264
rect 24577 1259 24643 1262
rect 24761 1259 24827 1262
rect 23565 914 23631 917
rect 27520 914 28000 944
rect 23565 912 28000 914
rect 23565 856 23570 912
rect 23626 856 28000 912
rect 23565 854 28000 856
rect 23565 851 23631 854
rect 27520 824 28000 854
rect 24577 370 24643 373
rect 27520 370 28000 400
rect 24577 368 28000 370
rect 24577 312 24582 368
rect 24638 312 28000 368
rect 24577 310 28000 312
rect 24577 307 24643 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 20116 18532 20180 18596
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 14412 16900 14476 16964
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 20116 12276 20180 12340
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 14412 10160 14476 10164
rect 14412 10104 14462 10160
rect 14462 10104 14476 10160
rect 14412 10100 14476 10104
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14411 16964 14477 16965
rect 14411 16900 14412 16964
rect 14476 16900 14477 16964
rect 14411 16899 14477 16900
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 14414 10165 14474 16899
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14411 10164 14477 10165
rect 14411 10100 14412 10164
rect 14476 10100 14477 10164
rect 14411 10099 14477 10100
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 20115 18596 20181 18597
rect 20115 18532 20116 18596
rect 20180 18532 20181 18596
rect 20115 18531 20181 18532
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 20118 12341 20178 18531
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 20115 12340 20181 12341
rect 20115 12276 20116 12340
rect 20180 12276 20181 12340
rect 20115 12275 20181 12276
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_buf_2  _059_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__059__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3312 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_22 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_26 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3496 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_30 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _060_
timestamp 1586364061
transform 1 0 5520 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_52
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _061_
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_80
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_1.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_91
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_92
timestamp 1586364061
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_104
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_108
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_conb_1  _049_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_126
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_130
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_135
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_139
timestamp 1586364061
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 15640 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_165
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l3_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_169
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_171
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_192
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_205
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_209
timestamp 1586364061
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_215
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20700 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_222
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_222
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21344 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_226
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_230
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_228
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_243
timestamp 1586364061
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23276 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23828 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_267
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_263
timestamp 1586364061
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_259
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_271
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_1  mux_bottom_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_116
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_128
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_132
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_162
timestamp 1586364061
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_185
timestamp 1586364061
transform 1 0 18124 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_191
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22356 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22724 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_229
timestamp 1586364061
transform 1 0 22172 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_233
timestamp 1586364061
transform 1 0 22540 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_237
timestamp 1586364061
transform 1 0 22908 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24288 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_250
timestamp 1586364061
transform 1 0 24104 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_254
timestamp 1586364061
transform 1 0 24472 0 -1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_224
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_228
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_237
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_241
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_264
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_139
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_164
timestamp 1586364061
transform 1 0 16192 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_181
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_198
timestamp 1586364061
transform 1 0 19320 0 -1 4896
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_203
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_207
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_234
timestamp 1586364061
transform 1 0 22632 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_238
timestamp 1586364061
transform 1 0 23000 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23368 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_261
timestamp 1586364061
transform 1 0 25116 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_4_273
timestamp 1586364061
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 774 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_106
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12512 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_133
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_137
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_164
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_201
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_218
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_222
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23828 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_270
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_148
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_139
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_142
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_152
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_187
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_192
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_196
timestamp 1586364061
transform 1 0 19136 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18952 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _083_
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19504 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_223
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_219
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_236
timestamp 1586364061
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23000 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_240
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_254
timestamp 1586364061
transform 1 0 24472 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24656 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24196 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_260
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_265
timestamp 1586364061
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_276
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_273
timestamp 1586364061
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_264
timestamp 1586364061
transform 1 0 25392 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15364 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_168
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_181
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_4  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21160 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22724 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22172 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22540 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_231
timestamp 1586364061
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  mux_bottom_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_265
timestamp 1586364061
transform 1 0 25484 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_191
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_195
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_222
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_265
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_126
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_130
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 406 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_161
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_177
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_183
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_194
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_198
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_201
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22632 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22356 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_226
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_233
timestamp 1586364061
transform 1 0 22540 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_257
timestamp 1586364061
transform 1 0 24748 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_261
timestamp 1586364061
transform 1 0 25116 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_10_273
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 774 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_146
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_169
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_201
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_223
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 24104 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_133
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_173
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_177
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 590 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_226
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_230
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_243
timestamp 1586364061
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_260
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_264
timestamp 1586364061
transform 1 0 25392 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_144
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_180
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_197
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_201
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_209
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_222
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_226
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_230
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22080 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_235
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22908 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 25392 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_262
timestamp 1586364061
transform 1 0 25208 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_266
timestamp 1586364061
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1786 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 590 592
use scs8hd_buf_1  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_137
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18952 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_213
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_230
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_234
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_238
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_264
timestamp 1586364061
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_268
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_272
timestamp 1586364061
transform 1 0 26128 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_115
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_128
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_196
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_200
timestamp 1586364061
transform 1 0 19504 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 1786 592
use scs8hd_buf_1  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_222
timestamp 1586364061
transform 1 0 21528 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_226
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 24748 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_249
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_253
timestamp 1586364061
transform 1 0 24380 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_266
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_128
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_155
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_203
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_207
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_230
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_17_270
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_128
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_177
timestamp 1586364061
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 18124 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_181
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_188
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_192
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21068 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_236
timestamp 1586364061
transform 1 0 22816 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_1  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_165
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_161
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_169
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_187
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_buf_1  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_193
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_191
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_204
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_228
timestamp 1586364061
transform 1 0 22080 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_225
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_221
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_231
timestamp 1586364061
transform 1 0 22356 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22172 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 22632 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_1  mux_right_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22172 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_243
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _062_
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_129
timestamp 1586364061
transform 1 0 12972 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 774 592
use scs8hd_buf_1  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_149
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_155
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_168
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_176
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_180
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_224
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 590 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_266
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_270
timestamp 1586364061
transform 1 0 25944 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_1  mux_right_track_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_133
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 774 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_4  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 15732 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_161
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_181
timestamp 1586364061
transform 1 0 17756 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_191
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_204
timestamp 1586364061
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 22724 0 -1 14688
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_22_219
timestamp 1586364061
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_231
timestamp 1586364061
transform 1 0 22356 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_254
timestamp 1586364061
transform 1 0 24472 0 -1 14688
box -38 -48 774 592
use scs8hd_buf_2  _063_
timestamp 1586364061
transform 1 0 25208 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_266
timestamp 1586364061
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_buf_1  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 590 592
use scs8hd_conb_1  _031_
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_156
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_160
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_173
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_177
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_26.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_181
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_23_219
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_223
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_228
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_259
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_263
timestamp 1586364061
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_1  mux_right_track_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_26.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_170
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_193
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_197
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 406 592
use scs8hd_conb_1  _032_
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_26.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20148 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_209
timestamp 1586364061
transform 1 0 20332 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_213
timestamp 1586364061
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_218
timestamp 1586364061
transform 1 0 21160 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21344 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_222
timestamp 1586364061
transform 1 0 21528 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_245
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_253
timestamp 1586364061
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 774 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_106
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_130
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_160
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18584 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_199
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_216
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21712 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_233
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_237
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 406 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24196 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_241
timestamp 1586364061
transform 1 0 23276 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_249
timestamp 1586364061
transform 1 0 24012 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_263
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_267
timestamp 1586364061
transform 1 0 25668 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_275
timestamp 1586364061
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 11316 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_120
timestamp 1586364061
transform 1 0 12144 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_133
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_146
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_142
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_168
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_169
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_178
timestamp 1586364061
transform 1 0 17480 0 1 16864
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_194
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_188
timestamp 1586364061
transform 1 0 18400 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_214
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21160 0 1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 22540 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 22908 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_234
timestamp 1586364061
transform 1 0 22632 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_238
timestamp 1586364061
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_227
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_231
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_235
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_239
timestamp 1586364061
transform 1 0 23092 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_242
timestamp 1586364061
transform 1 0 23368 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23460 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_26_256
timestamp 1586364061
transform 1 0 24656 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_252
timestamp 1586364061
transform 1 0 24288 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24472 0 -1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_22.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_264
timestamp 1586364061
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_264
timestamp 1586364061
transform 1 0 25392 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _067_
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_27_268
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_272
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_132
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16928 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_167
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_171
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_191
timestamp 1586364061
transform 1 0 18676 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_28_197
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 590 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_buf_1  mux_right_track_22.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_228
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_236
timestamp 1586364061
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_2  _066_
timestamp 1586364061
transform 1 0 24748 0 -1 17952
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23184 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_249
timestamp 1586364061
transform 1 0 24012 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_253
timestamp 1586364061
transform 1 0 24380 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_261
timestamp 1586364061
transform 1 0 25116 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_273
timestamp 1586364061
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_94
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use scs8hd_buf_1  mux_right_track_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13340 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16284 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_163
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_167
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_178
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 1786 592
use scs8hd_buf_1  mux_right_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_187
timestamp 1586364061
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_191
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_214
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 22908 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_231
timestamp 1586364061
transform 1 0 22356 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_235
timestamp 1586364061
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_239
timestamp 1586364061
transform 1 0 23092 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_254
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _065_
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_270
timestamp 1586364061
transform 1 0 25944 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_276
timestamp 1586364061
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10580 0 -1 19040
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_30_101
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12512 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_122
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_126
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_134
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15364 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_164
timestamp 1586364061
transform 1 0 16192 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_170
timestamp 1586364061
transform 1 0 16744 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_192
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_196
timestamp 1586364061
transform 1 0 19136 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 866 592
use scs8hd_buf_1  mux_right_track_20.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_200
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_conb_1  _030_
timestamp 1586364061
transform 1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22172 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22540 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_231
timestamp 1586364061
transform 1 0 22356 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_235
timestamp 1586364061
transform 1 0 22724 0 -1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_22.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_266
timestamp 1586364061
transform 1 0 25576 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_91
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_108
timestamp 1586364061
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_112
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_138
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _028_
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_165
timestamp 1586364061
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_169
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19688 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_211
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21252 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22264 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_228
timestamp 1586364061
transform 1 0 22080 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_236
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23920 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _064_
timestamp 1586364061
transform 1 0 25484 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25300 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 26036 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_261
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_273
timestamp 1586364061
transform 1 0 26220 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10028 0 -1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_32_116
timestamp 1586364061
transform 1 0 11776 0 -1 20128
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15364 0 -1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_174
timestamp 1586364061
transform 1 0 17112 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17664 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_182
timestamp 1586364061
transform 1 0 17848 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_199
timestamp 1586364061
transform 1 0 19412 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_204
timestamp 1586364061
transform 1 0 19872 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_208
timestamp 1586364061
transform 1 0 20240 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22816 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_234
timestamp 1586364061
transform 1 0 22632 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_238
timestamp 1586364061
transform 1 0 23000 0 -1 20128
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_20.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23920 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23736 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_267
timestamp 1586364061
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_buf_2  _057_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use scs8hd_buf_2  _058_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_19
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 314 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_103
timestamp 1586364061
transform 1 0 10580 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_136
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_132
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_143
timestamp 1586364061
transform 1 0 14260 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_144
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_140
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 13984 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_34_167
timestamp 1586364061
transform 1 0 16468 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_166
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16560 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16560 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_174
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_170
timestamp 1586364061
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_174
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_170
timestamp 1586364061
transform 1 0 16744 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16928 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17204 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18768 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_184
timestamp 1586364061
transform 1 0 18032 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_188
timestamp 1586364061
transform 1 0 18400 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_191
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_205
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_201
timestamp 1586364061
transform 1 0 19596 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_207
timestamp 1586364061
transform 1 0 20148 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_203
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19780 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20516 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_227
timestamp 1586364061
transform 1 0 21988 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_224
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21620 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21804 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_236
timestamp 1586364061
transform 1 0 22816 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_231
timestamp 1586364061
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22172 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _029_
timestamp 1586364061
transform 1 0 22540 0 1 20128
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_18.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21804 0 -1 21216
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_34_244
timestamp 1586364061
transform 1 0 23552 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23736 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_248
timestamp 1586364061
transform 1 0 23920 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24104 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23920 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24104 0 1 20128
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24288 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_267
timestamp 1586364061
transform 1 0 25668 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_263
timestamp 1586364061
transform 1 0 25300 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_259
timestamp 1586364061
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 25484 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 25116 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_273
timestamp 1586364061
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_271
timestamp 1586364061
transform 1 0 26036 0 1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_261
timestamp 1586364061
transform 1 0 25116 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10672 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_141
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_145
timestamp 1586364061
transform 1 0 14444 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_158
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17296 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_170
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_174
timestamp 1586364061
transform 1 0 17112 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_178
timestamp 1586364061
transform 1 0 17480 0 1 21216
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18952 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 18768 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18400 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_190
timestamp 1586364061
transform 1 0 18584 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_213
timestamp 1586364061
transform 1 0 20700 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_223
timestamp 1586364061
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_20.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24104 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23920 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23092 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_241
timestamp 1586364061
transform 1 0 23276 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12052 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15364 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14904 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13892 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16928 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_164
timestamp 1586364061
transform 1 0 16192 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_168
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18492 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_181
timestamp 1586364061
transform 1 0 17756 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_198
timestamp 1586364061
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 20976 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20148 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19504 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_206
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_209
timestamp 1586364061
transform 1 0 20332 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_1  mux_right_track_18.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22080 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21528 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22908 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22540 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_220
timestamp 1586364061
transform 1 0 21344 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_224
timestamp 1586364061
transform 1 0 21712 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_231
timestamp 1586364061
transform 1 0 22356 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_235
timestamp 1586364061
transform 1 0 22724 0 -1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_18.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1786 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_258
timestamp 1586364061
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_270
timestamp 1586364061
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_104
timestamp 1586364061
transform 1 0 10672 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_107
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_111
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_119
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1586364061
transform 1 0 14904 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_142
timestamp 1586364061
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_146
timestamp 1586364061
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16284 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_163
timestamp 1586364061
transform 1 0 16100 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_167
timestamp 1586364061
transform 1 0 16468 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_193
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_197
timestamp 1586364061
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20148 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19964 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_201
timestamp 1586364061
transform 1 0 19596 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22908 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22540 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 22080 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_226
timestamp 1586364061
transform 1 0 21896 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_230
timestamp 1586364061
transform 1 0 22264 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_235
timestamp 1586364061
transform 1 0 22724 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_239
timestamp 1586364061
transform 1 0 23092 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_254
timestamp 1586364061
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _056_
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_37_266
timestamp 1586364061
transform 1 0 25576 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_37_274
timestamp 1586364061
transform 1 0 26312 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13248 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13064 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_124
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_128
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14260 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_152
timestamp 1586364061
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_149
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 14904 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_158
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 15456 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15824 0 -1 23392
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18308 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_179
timestamp 1586364061
transform 1 0 17572 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_183
timestamp 1586364061
transform 1 0 17940 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_186
timestamp 1586364061
transform 1 0 18216 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_206
timestamp 1586364061
transform 1 0 20056 0 -1 23392
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1586364061
transform 1 0 22908 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_12  FILLER_38_224
timestamp 1586364061
transform 1 0 21712 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_236
timestamp 1586364061
transform 1 0 22816 0 -1 23392
box -38 -48 130 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 24472 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23920 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24288 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_246
timestamp 1586364061
transform 1 0 23736 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_250
timestamp 1586364061
transform 1 0 24104 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_258
timestamp 1586364061
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_270
timestamp 1586364061
transform 1 0 25944 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11868 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_106
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_119
timestamp 1586364061
transform 1 0 12052 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13432 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13248 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_126
timestamp 1586364061
transform 1 0 12696 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_130
timestamp 1586364061
transform 1 0 13064 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_143
timestamp 1586364061
transform 1 0 14260 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_146
timestamp 1586364061
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_152
timestamp 1586364061
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_149
timestamp 1586364061
transform 1 0 14812 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 14904 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1586364061
transform 1 0 14904 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_167
timestamp 1586364061
transform 1 0 16468 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_163
timestamp 1586364061
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15824 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_177
timestamp 1586364061
transform 1 0 17388 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_169
timestamp 1586364061
transform 1 0 16652 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17204 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17572 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 17756 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_196
timestamp 1586364061
transform 1 0 19136 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_190
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18952 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18952 0 1 23392
box -38 -48 1786 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 19596 0 -1 24480
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_213
timestamp 1586364061
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_217
timestamp 1586364061
transform 1 0 21068 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_200
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_205
timestamp 1586364061
transform 1 0 19964 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_224
timestamp 1586364061
transform 1 0 21712 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_224
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 21252 0 1 23392
box -38 -48 222 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 21436 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_235
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_228
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 22448 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_236
timestamp 1586364061
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 23460 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_247
timestamp 1586364061
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 23828 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_259
timestamp 1586364061
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 12788 0 1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 13340 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_131
timestamp 1586364061
transform 1 0 13156 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 314 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 14352 0 1 24480
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15456 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 15272 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_140
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_148
timestamp 1586364061
transform 1 0 14720 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_152
timestamp 1586364061
transform 1 0 15088 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 16652 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_165
timestamp 1586364061
transform 1 0 16284 0 1 24480
box -38 -48 406 592
use scs8hd_decap_6  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 590 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_179
timestamp 1586364061
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_193
timestamp 1586364061
transform 1 0 18860 0 1 24480
box -38 -48 590 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 21068 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 19964 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 20516 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 19412 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_201
timestamp 1586364061
transform 1 0 19596 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_209
timestamp 1586364061
transform 1 0 20332 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_213
timestamp 1586364061
transform 1 0 20700 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 22172 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 21620 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 22724 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 21988 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_221
timestamp 1586364061
transform 1 0 21436 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_225
timestamp 1586364061
transform 1 0 21804 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_233
timestamp 1586364061
transform 1 0 22540 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_237
timestamp 1586364061
transform 1 0 22908 0 1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_243
timestamp 1586364061
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 590 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 14260 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_147
timestamp 1586364061
transform 1 0 14628 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 16652 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16008 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_160
timestamp 1586364061
transform 1 0 15824 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_164
timestamp 1586364061
transform 1 0 16192 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_173
timestamp 1586364061
transform 1 0 17020 0 -1 25568
box -38 -48 774 592
use scs8hd_conb_1  _033_
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_181
timestamp 1586364061
transform 1 0 17756 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_190
timestamp 1586364061
transform 1 0 18584 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_198
timestamp 1586364061
transform 1 0 19320 0 -1 25568
box -38 -48 130 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_203
timestamp 1586364061
transform 1 0 19780 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_42_215
timestamp 1586364061
transform 1 0 20884 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 21988 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_226
timestamp 1586364061
transform 1 0 21896 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_231
timestamp 1586364061
transform 1 0 22356 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_243
timestamp 1586364061
transform 1 0 23460 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_247
timestamp 1586364061
transform 1 0 23828 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 13880 480 14000 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 23264 480 23384 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 27520 280 28000 400 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 27520 6672 28000 6792 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 27520 11296 28000 11416 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 27520 824 28000 944 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 27520 5448 28000 5568 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 27520 17688 28000 17808 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 27520 18368 28000 18488 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 27520 19456 28000 19576 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 27520 21224 28000 21344 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 27520 17144 28000 17264 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1582 0 1638 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 24122 0 24178 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 26146 0 26202 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 26882 0 26938 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 27526 0 27582 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 938 27520 994 28000 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 7746 27520 7802 28000 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 9126 27520 9182 28000 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 11150 27520 11206 28000 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1582 27520 1638 28000 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2962 27520 3018 28000 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4986 27520 5042 28000 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 5722 27520 5778 28000 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 22742 27520 22798 28000 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 23478 27520 23534 28000 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 25502 27520 25558 28000 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 26146 27520 26202 28000 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 26882 27520 26938 28000 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 27526 27520 27582 28000 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 15290 27520 15346 28000 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 17314 27520 17370 28000 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 19338 27520 19394 28000 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 20718 27520 20774 28000 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 prog_clk
port 123 nsew default input
rlabel metal3 s 27520 23536 28000 23656 6 right_top_grid_pin_42_
port 124 nsew default input
rlabel metal3 s 27520 24080 28000 24200 6 right_top_grid_pin_43_
port 125 nsew default input
rlabel metal3 s 27520 24760 28000 24880 6 right_top_grid_pin_44_
port 126 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_top_grid_pin_45_
port 127 nsew default input
rlabel metal3 s 27520 25848 28000 25968 6 right_top_grid_pin_46_
port 128 nsew default input
rlabel metal3 s 27520 26528 28000 26648 6 right_top_grid_pin_47_
port 129 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_top_grid_pin_48_
port 130 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_49_
port 131 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 133 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
