magic
tech EFS8A
magscale 1 2
timestamp 1603803961
<< locali >>
rect 7205 33371 7239 33609
rect 9873 23511 9907 23613
rect 9229 12087 9263 12393
rect 9137 11611 9171 11849
rect 8953 6103 8987 6409
<< viali >>
rect 9664 36669 9698 36703
rect 9735 36533 9769 36567
rect 10149 36533 10183 36567
rect 8677 36329 8711 36363
rect 8309 36261 8343 36295
rect 7516 36193 7550 36227
rect 8493 36193 8527 36227
rect 9756 36193 9790 36227
rect 7619 36057 7653 36091
rect 9827 35989 9861 36023
rect 10241 35989 10275 36023
rect 7757 35785 7791 35819
rect 9321 35785 9355 35819
rect 7021 35717 7055 35751
rect 8769 35649 8803 35683
rect 10333 35649 10367 35683
rect 10793 35649 10827 35683
rect 6837 35581 6871 35615
rect 7389 35581 7423 35615
rect 8309 35513 8343 35547
rect 8401 35513 8435 35547
rect 10149 35513 10183 35547
rect 10425 35513 10459 35547
rect 9781 35445 9815 35479
rect 6055 35241 6089 35275
rect 9045 35241 9079 35275
rect 10241 35241 10275 35275
rect 13185 35241 13219 35275
rect 8217 35173 8251 35207
rect 10609 35173 10643 35207
rect 5984 35105 6018 35139
rect 6929 35105 6963 35139
rect 12056 35105 12090 35139
rect 13001 35105 13035 35139
rect 8125 35037 8159 35071
rect 8401 35037 8435 35071
rect 10517 35037 10551 35071
rect 11161 35037 11195 35071
rect 7113 34969 7147 35003
rect 7573 34901 7607 34935
rect 12127 34901 12161 34935
rect 8953 34697 8987 34731
rect 9321 34697 9355 34731
rect 12633 34697 12667 34731
rect 5825 34629 5859 34663
rect 7665 34561 7699 34595
rect 8033 34561 8067 34595
rect 10333 34561 10367 34595
rect 10793 34561 10827 34595
rect 5641 34493 5675 34527
rect 6193 34493 6227 34527
rect 6653 34493 6687 34527
rect 8677 34493 8711 34527
rect 9137 34493 9171 34527
rect 9689 34493 9723 34527
rect 12081 34493 12115 34527
rect 12449 34493 12483 34527
rect 13001 34493 13035 34527
rect 13369 34493 13403 34527
rect 7481 34425 7515 34459
rect 7757 34425 7791 34459
rect 10425 34425 10459 34459
rect 7113 34357 7147 34391
rect 10149 34357 10183 34391
rect 11253 34357 11287 34391
rect 5319 34153 5353 34187
rect 13185 34153 13219 34187
rect 6377 34085 6411 34119
rect 7941 34085 7975 34119
rect 10051 34085 10085 34119
rect 11621 34085 11655 34119
rect 5248 34017 5282 34051
rect 10609 34017 10643 34051
rect 13001 34017 13035 34051
rect 6285 33949 6319 33983
rect 7849 33949 7883 33983
rect 8493 33949 8527 33983
rect 9689 33949 9723 33983
rect 11529 33949 11563 33983
rect 11805 33949 11839 33983
rect 6837 33881 6871 33915
rect 7573 33813 7607 33847
rect 10977 33813 11011 33847
rect 4859 33609 4893 33643
rect 6561 33609 6595 33643
rect 7205 33609 7239 33643
rect 7297 33609 7331 33643
rect 10241 33609 10275 33643
rect 11253 33609 11287 33643
rect 13461 33609 13495 33643
rect 5871 33541 5905 33575
rect 4756 33405 4790 33439
rect 5273 33405 5307 33439
rect 5800 33405 5834 33439
rect 7573 33473 7607 33507
rect 8033 33473 8067 33507
rect 8861 33473 8895 33507
rect 12541 33473 12575 33507
rect 12817 33473 12851 33507
rect 9321 33405 9355 33439
rect 11069 33405 11103 33439
rect 11621 33405 11655 33439
rect 5549 33337 5583 33371
rect 7205 33337 7239 33371
rect 7665 33337 7699 33371
rect 9683 33337 9717 33371
rect 12173 33337 12207 33371
rect 12633 33337 12667 33371
rect 6285 33269 6319 33303
rect 9229 33269 9263 33303
rect 10517 33269 10551 33303
rect 10977 33269 11011 33303
rect 5871 33065 5905 33099
rect 6193 33065 6227 33099
rect 7665 33065 7699 33099
rect 7941 33065 7975 33099
rect 8309 33065 8343 33099
rect 8631 33065 8665 33099
rect 10609 33065 10643 33099
rect 12541 33065 12575 33099
rect 7107 32997 7141 33031
rect 10010 32997 10044 33031
rect 11621 32997 11655 33031
rect 5800 32929 5834 32963
rect 8560 32929 8594 32963
rect 13068 32929 13102 32963
rect 6745 32861 6779 32895
rect 9689 32861 9723 32895
rect 11529 32861 11563 32895
rect 11805 32861 11839 32895
rect 8953 32725 8987 32759
rect 9321 32725 9355 32759
rect 11345 32725 11379 32759
rect 13139 32725 13173 32759
rect 7757 32521 7791 32555
rect 9505 32521 9539 32555
rect 11713 32521 11747 32555
rect 12587 32521 12621 32555
rect 8493 32453 8527 32487
rect 8585 32385 8619 32419
rect 6837 32317 6871 32351
rect 10609 32317 10643 32351
rect 10793 32317 10827 32351
rect 12484 32317 12518 32351
rect 7199 32249 7233 32283
rect 8125 32249 8159 32283
rect 8947 32249 8981 32283
rect 9781 32249 9815 32283
rect 10241 32249 10275 32283
rect 5825 32181 5859 32215
rect 6285 32181 6319 32215
rect 6561 32181 6595 32215
rect 10425 32181 10459 32215
rect 11345 32181 11379 32215
rect 12173 32181 12207 32215
rect 13093 32181 13127 32215
rect 9781 31977 9815 32011
rect 11391 31977 11425 32011
rect 11713 31977 11747 32011
rect 6837 31909 6871 31943
rect 7481 31909 7515 31943
rect 8401 31909 8435 31943
rect 10701 31909 10735 31943
rect 6101 31841 6135 31875
rect 6653 31841 6687 31875
rect 7941 31841 7975 31875
rect 8125 31841 8159 31875
rect 9965 31841 9999 31875
rect 10241 31841 10275 31875
rect 11288 31841 11322 31875
rect 7205 31637 7239 31671
rect 8677 31637 8711 31671
rect 5825 31433 5859 31467
rect 9781 31433 9815 31467
rect 7389 31297 7423 31331
rect 9321 31297 9355 31331
rect 10701 31297 10735 31331
rect 6929 31229 6963 31263
rect 7297 31229 7331 31263
rect 8677 31229 8711 31263
rect 9229 31229 9263 31263
rect 10149 31229 10183 31263
rect 8585 31161 8619 31195
rect 10517 31161 10551 31195
rect 10793 31161 10827 31195
rect 11345 31161 11379 31195
rect 6193 31093 6227 31127
rect 6653 31093 6687 31127
rect 7849 31093 7883 31127
rect 11621 31093 11655 31127
rect 7757 30889 7791 30923
rect 9505 30889 9539 30923
rect 10793 30889 10827 30923
rect 8217 30821 8251 30855
rect 9781 30821 9815 30855
rect 9873 30821 9907 30855
rect 11437 30821 11471 30855
rect 7021 30685 7055 30719
rect 8125 30685 8159 30719
rect 8401 30685 8435 30719
rect 10057 30685 10091 30719
rect 11345 30685 11379 30719
rect 11989 30685 12023 30719
rect 6929 30549 6963 30583
rect 11345 30345 11379 30379
rect 8999 30277 9033 30311
rect 10793 30277 10827 30311
rect 11621 30209 11655 30243
rect 7481 30141 7515 30175
rect 7757 30141 7791 30175
rect 8769 30141 8803 30175
rect 8896 30141 8930 30175
rect 9873 30141 9907 30175
rect 10235 30073 10269 30107
rect 7113 30005 7147 30039
rect 7573 30005 7607 30039
rect 8309 30005 8343 30039
rect 9321 30005 9355 30039
rect 9689 30005 9723 30039
rect 7481 29801 7515 29835
rect 7941 29801 7975 29835
rect 10977 29801 11011 29835
rect 10419 29733 10453 29767
rect 11989 29733 12023 29767
rect 6561 29665 6595 29699
rect 6929 29665 6963 29699
rect 8217 29665 8251 29699
rect 8585 29665 8619 29699
rect 7205 29597 7239 29631
rect 8769 29597 8803 29631
rect 9137 29597 9171 29631
rect 10057 29597 10091 29631
rect 11897 29597 11931 29631
rect 12173 29597 12207 29631
rect 5273 29461 5307 29495
rect 9965 29461 9999 29495
rect 8309 29257 8343 29291
rect 8677 29257 8711 29291
rect 9045 29257 9079 29291
rect 10425 29257 10459 29291
rect 11897 29257 11931 29291
rect 5089 29121 5123 29155
rect 5273 29121 5307 29155
rect 5917 29121 5951 29155
rect 7389 29121 7423 29155
rect 9137 29121 9171 29155
rect 10885 29121 10919 29155
rect 6561 29053 6595 29087
rect 10057 29053 10091 29087
rect 12173 29053 12207 29087
rect 5365 28985 5399 29019
rect 7297 28985 7331 29019
rect 7751 28985 7785 29019
rect 9499 28985 9533 29019
rect 10701 28917 10735 28951
rect 7481 28713 7515 28747
rect 8585 28713 8619 28747
rect 9965 28713 9999 28747
rect 11437 28713 11471 28747
rect 8027 28645 8061 28679
rect 4880 28577 4914 28611
rect 6377 28577 6411 28611
rect 6653 28577 6687 28611
rect 7665 28577 7699 28611
rect 8861 28577 8895 28611
rect 9689 28577 9723 28611
rect 10149 28577 10183 28611
rect 11253 28577 11287 28611
rect 6837 28509 6871 28543
rect 4951 28373 4985 28407
rect 5273 28373 5307 28407
rect 5641 28373 5675 28407
rect 7205 28373 7239 28407
rect 6193 28169 6227 28203
rect 8401 28169 8435 28203
rect 9137 28169 9171 28203
rect 10333 28169 10367 28203
rect 11069 28169 11103 28203
rect 7757 28101 7791 28135
rect 8125 28101 8159 28135
rect 5089 28033 5123 28067
rect 6837 28033 6871 28067
rect 8769 28033 8803 28067
rect 10057 28033 10091 28067
rect 4020 27965 4054 27999
rect 4445 27965 4479 27999
rect 9413 27965 9447 27999
rect 9781 27965 9815 27999
rect 10885 27965 10919 27999
rect 11713 27965 11747 27999
rect 5181 27897 5215 27931
rect 5733 27897 5767 27931
rect 6653 27897 6687 27931
rect 7199 27897 7233 27931
rect 4123 27829 4157 27863
rect 4905 27829 4939 27863
rect 11345 27829 11379 27863
rect 4813 27625 4847 27659
rect 5181 27625 5215 27659
rect 6377 27625 6411 27659
rect 6745 27625 6779 27659
rect 4399 27557 4433 27591
rect 5457 27557 5491 27591
rect 7021 27557 7055 27591
rect 9873 27557 9907 27591
rect 11437 27557 11471 27591
rect 4312 27489 4346 27523
rect 8436 27489 8470 27523
rect 12852 27489 12886 27523
rect 5365 27421 5399 27455
rect 5733 27421 5767 27455
rect 6929 27421 6963 27455
rect 9781 27421 9815 27455
rect 10425 27421 10459 27455
rect 11345 27421 11379 27455
rect 11989 27421 12023 27455
rect 7481 27353 7515 27387
rect 8539 27285 8573 27319
rect 9413 27285 9447 27319
rect 12955 27285 12989 27319
rect 3203 27081 3237 27115
rect 6285 27081 6319 27115
rect 7849 27081 7883 27115
rect 8539 27081 8573 27115
rect 11989 27081 12023 27115
rect 13277 27081 13311 27115
rect 13599 27081 13633 27115
rect 4537 27013 4571 27047
rect 5733 27013 5767 27047
rect 8861 27013 8895 27047
rect 10241 27013 10275 27047
rect 5181 26945 5215 26979
rect 6929 26945 6963 26979
rect 7205 26945 7239 26979
rect 10977 26945 11011 26979
rect 12587 26945 12621 26979
rect 3100 26877 3134 26911
rect 3525 26877 3559 26911
rect 4144 26877 4178 26911
rect 6561 26877 6595 26911
rect 8436 26877 8470 26911
rect 9229 26877 9263 26911
rect 11196 26877 11230 26911
rect 11621 26877 11655 26911
rect 12500 26877 12534 26911
rect 12909 26877 12943 26911
rect 13528 26877 13562 26911
rect 13921 26877 13955 26911
rect 5273 26809 5307 26843
rect 7021 26809 7055 26843
rect 9689 26809 9723 26843
rect 9781 26809 9815 26843
rect 10609 26809 10643 26843
rect 4215 26741 4249 26775
rect 4997 26741 5031 26775
rect 11299 26741 11333 26775
rect 5273 26537 5307 26571
rect 5641 26537 5675 26571
rect 7113 26537 7147 26571
rect 9505 26537 9539 26571
rect 11161 26537 11195 26571
rect 12909 26537 12943 26571
rect 4674 26469 4708 26503
rect 5917 26469 5951 26503
rect 6285 26469 6319 26503
rect 9137 26469 9171 26503
rect 9873 26469 9907 26503
rect 11345 26469 11379 26503
rect 11437 26469 11471 26503
rect 12449 26469 12483 26503
rect 7849 26401 7883 26435
rect 8309 26401 8343 26435
rect 10425 26401 10459 26435
rect 13093 26401 13127 26435
rect 13277 26401 13311 26435
rect 4353 26333 4387 26367
rect 6193 26333 6227 26367
rect 8401 26333 8435 26367
rect 9781 26333 9815 26367
rect 11621 26333 11655 26367
rect 6745 26265 6779 26299
rect 7573 26197 7607 26231
rect 10701 26197 10735 26231
rect 5181 25993 5215 26027
rect 6469 25993 6503 26027
rect 7481 25993 7515 26027
rect 9229 25993 9263 26027
rect 9597 25993 9631 26027
rect 10977 25993 11011 26027
rect 11621 25993 11655 26027
rect 6975 25925 7009 25959
rect 8125 25925 8159 25959
rect 9965 25925 9999 25959
rect 8309 25857 8343 25891
rect 12541 25857 12575 25891
rect 12817 25857 12851 25891
rect 4261 25789 4295 25823
rect 6904 25789 6938 25823
rect 10057 25789 10091 25823
rect 11345 25789 11379 25823
rect 4169 25721 4203 25755
rect 4623 25721 4657 25755
rect 8671 25721 8705 25755
rect 10378 25721 10412 25755
rect 12633 25721 12667 25755
rect 3801 25653 3835 25687
rect 5549 25653 5583 25687
rect 6101 25653 6135 25687
rect 7757 25653 7791 25687
rect 12173 25653 12207 25687
rect 13461 25653 13495 25687
rect 5825 25449 5859 25483
rect 8401 25449 8435 25483
rect 8953 25449 8987 25483
rect 9965 25449 9999 25483
rect 10977 25449 11011 25483
rect 13001 25449 13035 25483
rect 13691 25449 13725 25483
rect 3157 25381 3191 25415
rect 4353 25381 4387 25415
rect 5267 25381 5301 25415
rect 7107 25381 7141 25415
rect 10419 25381 10453 25415
rect 12126 25381 12160 25415
rect 2697 25313 2731 25347
rect 2973 25313 3007 25347
rect 10057 25313 10091 25347
rect 12725 25313 12759 25347
rect 13588 25313 13622 25347
rect 4905 25245 4939 25279
rect 6745 25245 6779 25279
rect 8493 25245 8527 25279
rect 11805 25245 11839 25279
rect 4721 25177 4755 25211
rect 6561 25109 6595 25143
rect 7665 25109 7699 25143
rect 7941 25109 7975 25143
rect 2513 24905 2547 24939
rect 2881 24905 2915 24939
rect 8217 24905 8251 24939
rect 10057 24905 10091 24939
rect 10333 24905 10367 24939
rect 11805 24905 11839 24939
rect 13553 24905 13587 24939
rect 5917 24769 5951 24803
rect 6193 24769 6227 24803
rect 7205 24769 7239 24803
rect 8861 24769 8895 24803
rect 9505 24769 9539 24803
rect 12173 24769 12207 24803
rect 3617 24701 3651 24735
rect 4169 24701 4203 24735
rect 5457 24701 5491 24735
rect 5641 24701 5675 24735
rect 10517 24701 10551 24735
rect 12541 24701 12575 24735
rect 12909 24701 12943 24735
rect 7297 24633 7331 24667
rect 7849 24633 7883 24667
rect 8677 24633 8711 24667
rect 8953 24633 8987 24667
rect 10838 24633 10872 24667
rect 3433 24565 3467 24599
rect 3893 24565 3927 24599
rect 4997 24565 5031 24599
rect 6653 24565 6687 24599
rect 11437 24565 11471 24599
rect 12541 24565 12575 24599
rect 8769 24361 8803 24395
rect 10517 24361 10551 24395
rect 12541 24361 12575 24395
rect 4813 24293 4847 24327
rect 6561 24293 6595 24327
rect 7205 24293 7239 24327
rect 10241 24293 10275 24327
rect 10977 24293 11011 24327
rect 11253 24293 11287 24327
rect 12771 24293 12805 24327
rect 2973 24225 3007 24259
rect 4077 24225 4111 24259
rect 4537 24225 4571 24259
rect 6009 24225 6043 24259
rect 8585 24225 8619 24259
rect 9689 24225 9723 24259
rect 12668 24225 12702 24259
rect 7113 24157 7147 24191
rect 11161 24157 11195 24191
rect 11529 24157 11563 24191
rect 6193 24089 6227 24123
rect 7665 24089 7699 24123
rect 9045 24089 9079 24123
rect 9873 24089 9907 24123
rect 3157 24021 3191 24055
rect 3709 24021 3743 24055
rect 5273 24021 5307 24055
rect 5549 24021 5583 24055
rect 6837 24021 6871 24055
rect 12081 24021 12115 24055
rect 2513 23817 2547 23851
rect 6653 23817 6687 23851
rect 11253 23817 11287 23851
rect 2789 23749 2823 23783
rect 11529 23749 11563 23783
rect 8953 23681 8987 23715
rect 10885 23681 10919 23715
rect 2605 23613 2639 23647
rect 3617 23613 3651 23647
rect 4169 23613 4203 23647
rect 5089 23613 5123 23647
rect 5457 23613 5491 23647
rect 5641 23613 5675 23647
rect 6285 23613 6319 23647
rect 6837 23613 6871 23647
rect 9873 23613 9907 23647
rect 10149 23613 10183 23647
rect 10609 23613 10643 23647
rect 12633 23613 12667 23647
rect 3065 23545 3099 23579
rect 5917 23545 5951 23579
rect 7158 23545 7192 23579
rect 8677 23545 8711 23579
rect 8769 23545 8803 23579
rect 9689 23545 9723 23579
rect 3433 23477 3467 23511
rect 3893 23477 3927 23511
rect 4721 23477 4755 23511
rect 7757 23477 7791 23511
rect 8033 23477 8067 23511
rect 8401 23477 8435 23511
rect 9873 23477 9907 23511
rect 10057 23477 10091 23511
rect 6193 23273 6227 23307
rect 7297 23273 7331 23307
rect 7941 23273 7975 23307
rect 8953 23273 8987 23307
rect 9873 23273 9907 23307
rect 12633 23273 12667 23307
rect 4997 23205 5031 23239
rect 6698 23205 6732 23239
rect 11161 23205 11195 23239
rect 11253 23205 11287 23239
rect 2973 23137 3007 23171
rect 6377 23137 6411 23171
rect 8125 23137 8159 23171
rect 9689 23137 9723 23171
rect 10149 23137 10183 23171
rect 4905 23069 4939 23103
rect 11529 23069 11563 23103
rect 5457 23001 5491 23035
rect 3157 22933 3191 22967
rect 3709 22933 3743 22967
rect 4261 22933 4295 22967
rect 4629 22933 4663 22967
rect 7573 22933 7607 22967
rect 8309 22933 8343 22967
rect 8585 22933 8619 22967
rect 2973 22729 3007 22763
rect 3525 22729 3559 22763
rect 5825 22729 5859 22763
rect 6469 22729 6503 22763
rect 8125 22729 8159 22763
rect 11437 22729 11471 22763
rect 12633 22729 12667 22763
rect 3801 22661 3835 22695
rect 13645 22661 13679 22695
rect 4629 22593 4663 22627
rect 7205 22593 7239 22627
rect 9873 22593 9907 22627
rect 10057 22593 10091 22627
rect 10425 22593 10459 22627
rect 3617 22525 3651 22559
rect 4077 22525 4111 22559
rect 5549 22525 5583 22559
rect 8493 22525 8527 22559
rect 8861 22525 8895 22559
rect 9505 22525 9539 22559
rect 9965 22525 9999 22559
rect 10241 22525 10275 22559
rect 12449 22525 12483 22559
rect 12909 22525 12943 22559
rect 13461 22525 13495 22559
rect 13921 22525 13955 22559
rect 4537 22457 4571 22491
rect 4991 22457 5025 22491
rect 6929 22457 6963 22491
rect 7021 22457 7055 22491
rect 9137 22457 9171 22491
rect 10977 22389 11011 22423
rect 11713 22389 11747 22423
rect 5457 22185 5491 22219
rect 6561 22185 6595 22219
rect 7665 22185 7699 22219
rect 9413 22185 9447 22219
rect 4899 22117 4933 22151
rect 10378 22117 10412 22151
rect 12541 22117 12575 22151
rect 6285 22049 6319 22083
rect 6837 22049 6871 22083
rect 8677 22049 8711 22083
rect 10057 22049 10091 22083
rect 11805 22049 11839 22083
rect 12081 22049 12115 22083
rect 4537 21981 4571 22015
rect 7389 21981 7423 22015
rect 8769 21981 8803 22015
rect 10977 21913 11011 21947
rect 11897 21913 11931 21947
rect 4353 21845 4387 21879
rect 9873 21845 9907 21879
rect 5273 21641 5307 21675
rect 9505 21641 9539 21675
rect 11069 21641 11103 21675
rect 6929 21573 6963 21607
rect 8493 21573 8527 21607
rect 10057 21573 10091 21607
rect 11345 21573 11379 21607
rect 12633 21573 12667 21607
rect 4813 21505 4847 21539
rect 7573 21505 7607 21539
rect 9137 21505 9171 21539
rect 4353 21437 4387 21471
rect 4721 21437 4755 21471
rect 6653 21437 6687 21471
rect 6837 21437 6871 21471
rect 7113 21437 7147 21471
rect 8401 21437 8435 21471
rect 8677 21437 8711 21471
rect 9965 21437 9999 21471
rect 10241 21437 10275 21471
rect 10701 21437 10735 21471
rect 12449 21437 12483 21471
rect 12909 21437 12943 21471
rect 6285 21369 6319 21403
rect 7941 21369 7975 21403
rect 12173 21369 12207 21403
rect 3801 21301 3835 21335
rect 4169 21301 4203 21335
rect 5825 21301 5859 21335
rect 8309 21301 8343 21335
rect 9781 21301 9815 21335
rect 11805 21301 11839 21335
rect 4261 21097 4295 21131
rect 6377 21097 6411 21131
rect 8677 21097 8711 21131
rect 10149 21097 10183 21131
rect 11713 21097 11747 21131
rect 12265 21097 12299 21131
rect 6745 21029 6779 21063
rect 10793 21029 10827 21063
rect 4445 20961 4479 20995
rect 4629 20961 4663 20995
rect 8160 20961 8194 20995
rect 10333 20961 10367 20995
rect 11253 20961 11287 20995
rect 11529 20961 11563 20995
rect 6653 20893 6687 20927
rect 8263 20893 8297 20927
rect 7205 20825 7239 20859
rect 11345 20825 11379 20859
rect 7573 20757 7607 20791
rect 9505 20757 9539 20791
rect 6285 20553 6319 20587
rect 9781 20553 9815 20587
rect 11989 20553 12023 20587
rect 5365 20485 5399 20519
rect 10057 20485 10091 20519
rect 7389 20417 7423 20451
rect 3776 20349 3810 20383
rect 8309 20349 8343 20383
rect 8769 20349 8803 20383
rect 9965 20349 9999 20383
rect 10241 20349 10275 20383
rect 3617 20281 3651 20315
rect 4813 20281 4847 20315
rect 4905 20281 4939 20315
rect 6929 20281 6963 20315
rect 7021 20281 7055 20315
rect 10701 20281 10735 20315
rect 11345 20281 11379 20315
rect 3847 20213 3881 20247
rect 4261 20213 4295 20247
rect 4629 20213 4663 20247
rect 6653 20213 6687 20247
rect 7849 20213 7883 20247
rect 8677 20213 8711 20247
rect 11713 20213 11747 20247
rect 4399 20009 4433 20043
rect 5089 20009 5123 20043
rect 6469 20009 6503 20043
rect 9505 20009 9539 20043
rect 2973 19941 3007 19975
rect 4721 19941 4755 19975
rect 5870 19941 5904 19975
rect 7481 19941 7515 19975
rect 4328 19873 4362 19907
rect 9873 19873 9907 19907
rect 10149 19873 10183 19907
rect 11437 19873 11471 19907
rect 5549 19805 5583 19839
rect 7389 19805 7423 19839
rect 10333 19805 10367 19839
rect 7941 19737 7975 19771
rect 9965 19737 9999 19771
rect 11621 19737 11655 19771
rect 6929 19669 6963 19703
rect 8401 19669 8435 19703
rect 5181 19465 5215 19499
rect 5641 19465 5675 19499
rect 7849 19465 7883 19499
rect 9689 19465 9723 19499
rect 10885 19465 10919 19499
rect 11529 19465 11563 19499
rect 6929 19329 6963 19363
rect 7573 19329 7607 19363
rect 8953 19329 8987 19363
rect 2697 19261 2731 19295
rect 3249 19261 3283 19295
rect 3801 19261 3835 19295
rect 4261 19261 4295 19295
rect 5917 19261 5951 19295
rect 8585 19261 8619 19295
rect 9229 19261 9263 19295
rect 10425 19261 10459 19295
rect 3433 19193 3467 19227
rect 4623 19193 4657 19227
rect 7021 19193 7055 19227
rect 8309 19193 8343 19227
rect 8401 19193 8435 19227
rect 10517 19193 10551 19227
rect 11161 19193 11195 19227
rect 2513 19125 2547 19159
rect 4169 19125 4203 19159
rect 6653 19125 6687 19159
rect 2789 18921 2823 18955
rect 3111 18921 3145 18955
rect 6469 18921 6503 18955
rect 8309 18921 8343 18955
rect 9413 18921 9447 18955
rect 10701 18921 10735 18955
rect 5870 18853 5904 18887
rect 7481 18853 7515 18887
rect 2028 18785 2062 18819
rect 3040 18785 3074 18819
rect 4572 18785 4606 18819
rect 9045 18785 9079 18819
rect 9689 18785 9723 18819
rect 9965 18785 9999 18819
rect 11345 18785 11379 18819
rect 3525 18717 3559 18751
rect 5549 18717 5583 18751
rect 7389 18717 7423 18751
rect 10425 18717 10459 18751
rect 4675 18649 4709 18683
rect 7941 18649 7975 18683
rect 9781 18649 9815 18683
rect 2099 18581 2133 18615
rect 4261 18581 4295 18615
rect 4997 18581 5031 18615
rect 5457 18581 5491 18615
rect 6837 18581 6871 18615
rect 11529 18581 11563 18615
rect 2605 18377 2639 18411
rect 3065 18377 3099 18411
rect 6009 18377 6043 18411
rect 6561 18377 6595 18411
rect 8033 18377 8067 18411
rect 8493 18377 8527 18411
rect 9597 18377 9631 18411
rect 9965 18377 9999 18411
rect 10425 18377 10459 18411
rect 11345 18377 11379 18411
rect 7757 18309 7791 18343
rect 8861 18309 8895 18343
rect 4169 18241 4203 18275
rect 9229 18241 9263 18275
rect 9689 18241 9723 18275
rect 2421 18173 2455 18207
rect 3433 18173 3467 18207
rect 3893 18173 3927 18207
rect 4997 18173 5031 18207
rect 5549 18173 5583 18207
rect 6837 18173 6871 18207
rect 9468 18173 9502 18207
rect 10885 18173 10919 18207
rect 11713 18173 11747 18207
rect 12449 18173 12483 18207
rect 12909 18173 12943 18207
rect 2053 18105 2087 18139
rect 5733 18105 5767 18139
rect 7158 18105 7192 18139
rect 9321 18105 9355 18139
rect 4537 18037 4571 18071
rect 10701 18037 10735 18071
rect 11069 18037 11103 18071
rect 12633 18037 12667 18071
rect 3157 17833 3191 17867
rect 3433 17833 3467 17867
rect 4215 17833 4249 17867
rect 6101 17833 6135 17867
rect 6561 17833 6595 17867
rect 9413 17833 9447 17867
rect 13277 17833 13311 17867
rect 4905 17765 4939 17799
rect 5825 17765 5859 17799
rect 6837 17765 6871 17799
rect 7389 17765 7423 17799
rect 8125 17765 8159 17799
rect 8217 17765 8251 17799
rect 10793 17765 10827 17799
rect 2973 17697 3007 17731
rect 4144 17697 4178 17731
rect 5089 17697 5123 17731
rect 5549 17697 5583 17731
rect 8401 17697 8435 17731
rect 9689 17697 9723 17731
rect 9965 17697 9999 17731
rect 11529 17697 11563 17731
rect 12817 17697 12851 17731
rect 13093 17697 13127 17731
rect 6745 17629 6779 17663
rect 10149 17629 10183 17663
rect 11253 17629 11287 17663
rect 7757 17561 7791 17595
rect 9781 17561 9815 17595
rect 12909 17561 12943 17595
rect 2513 17493 2547 17527
rect 4629 17493 4663 17527
rect 8493 17493 8527 17527
rect 4169 17289 4203 17323
rect 5273 17289 5307 17323
rect 5641 17289 5675 17323
rect 8309 17289 8343 17323
rect 10057 17289 10091 17323
rect 10425 17289 10459 17323
rect 11621 17289 11655 17323
rect 13553 17289 13587 17323
rect 3065 17221 3099 17255
rect 6285 17221 6319 17255
rect 10701 17221 10735 17255
rect 13185 17221 13219 17255
rect 3801 17153 3835 17187
rect 7573 17153 7607 17187
rect 9597 17153 9631 17187
rect 4537 17085 4571 17119
rect 4721 17085 4755 17119
rect 7113 17085 7147 17119
rect 7205 17085 7239 17119
rect 7389 17085 7423 17119
rect 8953 17085 8987 17119
rect 9505 17085 9539 17119
rect 10609 17085 10643 17119
rect 10885 17085 10919 17119
rect 4997 17017 5031 17051
rect 6653 17017 6687 17051
rect 9597 16949 9631 16983
rect 11069 16949 11103 16983
rect 12909 16949 12943 16983
rect 5273 16745 5307 16779
rect 5825 16745 5859 16779
rect 7205 16745 7239 16779
rect 8033 16745 8067 16779
rect 8769 16745 8803 16779
rect 9137 16745 9171 16779
rect 10793 16745 10827 16779
rect 13691 16745 13725 16779
rect 9505 16677 9539 16711
rect 11989 16677 12023 16711
rect 4261 16609 4295 16643
rect 4721 16609 4755 16643
rect 6653 16609 6687 16643
rect 7573 16609 7607 16643
rect 7849 16609 7883 16643
rect 9689 16609 9723 16643
rect 9965 16609 9999 16643
rect 11069 16609 11103 16643
rect 11897 16609 11931 16643
rect 13588 16609 13622 16643
rect 4813 16541 4847 16575
rect 6745 16541 6779 16575
rect 7665 16541 7699 16575
rect 10425 16541 10459 16575
rect 9781 16473 9815 16507
rect 3755 16201 3789 16235
rect 4537 16201 4571 16235
rect 6101 16201 6135 16235
rect 7941 16201 7975 16235
rect 10149 16201 10183 16235
rect 13553 16201 13587 16235
rect 6561 16133 6595 16167
rect 4169 16065 4203 16099
rect 4629 16065 4663 16099
rect 9413 16065 9447 16099
rect 10885 16065 10919 16099
rect 12449 16065 12483 16099
rect 3525 15997 3559 16031
rect 3652 15997 3686 16031
rect 6837 15997 6871 16031
rect 7389 15997 7423 16031
rect 8861 15997 8895 16031
rect 9505 15997 9539 16031
rect 4991 15929 5025 15963
rect 8585 15929 8619 15963
rect 10977 15929 11011 15963
rect 11529 15929 11563 15963
rect 5549 15861 5583 15895
rect 7113 15861 7147 15895
rect 9597 15861 9631 15895
rect 10701 15861 10735 15895
rect 11897 15861 11931 15895
rect 4353 15657 4387 15691
rect 7757 15657 7791 15691
rect 9045 15657 9079 15691
rect 9505 15657 9539 15691
rect 11161 15657 11195 15691
rect 4991 15589 5025 15623
rect 6561 15589 6595 15623
rect 10194 15589 10228 15623
rect 11805 15589 11839 15623
rect 4629 15521 4663 15555
rect 7941 15521 7975 15555
rect 8217 15521 8251 15555
rect 9873 15521 9907 15555
rect 10793 15521 10827 15555
rect 2973 15453 3007 15487
rect 6469 15453 6503 15487
rect 6929 15453 6963 15487
rect 8401 15453 8435 15487
rect 11713 15453 11747 15487
rect 11989 15453 12023 15487
rect 5549 15385 5583 15419
rect 8033 15385 8067 15419
rect 6193 15317 6227 15351
rect 7481 15317 7515 15351
rect 3893 15113 3927 15147
rect 5273 15113 5307 15147
rect 5549 15113 5583 15147
rect 6561 15113 6595 15147
rect 7941 15113 7975 15147
rect 8309 15113 8343 15147
rect 9413 15113 9447 15147
rect 10241 15113 10275 15147
rect 11069 15113 11103 15147
rect 11805 15113 11839 15147
rect 5917 15045 5951 15079
rect 6285 15045 6319 15079
rect 7205 14977 7239 15011
rect 2697 14909 2731 14943
rect 2973 14909 3007 14943
rect 3985 14909 4019 14943
rect 5733 14909 5767 14943
rect 8401 14909 8435 14943
rect 8861 14909 8895 14943
rect 10701 14909 10735 14943
rect 11437 14909 11471 14943
rect 2329 14841 2363 14875
rect 3157 14841 3191 14875
rect 3433 14841 3467 14875
rect 4306 14841 4340 14875
rect 6929 14841 6963 14875
rect 7021 14841 7055 14875
rect 4905 14773 4939 14807
rect 8493 14773 8527 14807
rect 9873 14773 9907 14807
rect 12173 14773 12207 14807
rect 2513 14569 2547 14603
rect 6837 14569 6871 14603
rect 7205 14569 7239 14603
rect 8861 14569 8895 14603
rect 9505 14569 9539 14603
rect 4721 14501 4755 14535
rect 7618 14501 7652 14535
rect 10010 14501 10044 14535
rect 6285 14433 6319 14467
rect 7297 14433 7331 14467
rect 9689 14433 9723 14467
rect 11472 14433 11506 14467
rect 4629 14365 4663 14399
rect 4905 14365 4939 14399
rect 6469 14297 6503 14331
rect 5549 14229 5583 14263
rect 6101 14229 6135 14263
rect 8217 14229 8251 14263
rect 8585 14229 8619 14263
rect 10609 14229 10643 14263
rect 11575 14229 11609 14263
rect 4629 14025 4663 14059
rect 6377 14025 6411 14059
rect 7205 14025 7239 14059
rect 9045 14025 9079 14059
rect 10977 14025 11011 14059
rect 5825 13957 5859 13991
rect 11437 13957 11471 13991
rect 3525 13889 3559 13923
rect 5273 13889 5307 13923
rect 7297 13889 7331 13923
rect 8493 13889 8527 13923
rect 9689 13889 9723 13923
rect 9965 13889 9999 13923
rect 3617 13821 3651 13855
rect 4077 13821 4111 13855
rect 8217 13821 8251 13855
rect 9413 13821 9447 13855
rect 5365 13753 5399 13787
rect 7618 13753 7652 13787
rect 10057 13753 10091 13787
rect 10609 13753 10643 13787
rect 3893 13685 3927 13719
rect 5089 13685 5123 13719
rect 3111 13481 3145 13515
rect 4629 13481 4663 13515
rect 7389 13481 7423 13515
rect 7757 13481 7791 13515
rect 3617 13413 3651 13447
rect 5410 13413 5444 13447
rect 8217 13413 8251 13447
rect 10057 13413 10091 13447
rect 10609 13413 10643 13447
rect 3008 13345 3042 13379
rect 4144 13345 4178 13379
rect 11472 13345 11506 13379
rect 5089 13277 5123 13311
rect 6837 13277 6871 13311
rect 8125 13277 8159 13311
rect 8769 13277 8803 13311
rect 9965 13277 9999 13311
rect 11575 13277 11609 13311
rect 4215 13209 4249 13243
rect 4905 13141 4939 13175
rect 6009 13141 6043 13175
rect 9045 13141 9079 13175
rect 2973 12937 3007 12971
rect 3433 12937 3467 12971
rect 6193 12937 6227 12971
rect 8125 12937 8159 12971
rect 8401 12937 8435 12971
rect 5089 12869 5123 12903
rect 11437 12869 11471 12903
rect 4353 12801 4387 12835
rect 5273 12801 5307 12835
rect 5641 12801 5675 12835
rect 6837 12801 6871 12835
rect 8677 12801 8711 12835
rect 8953 12801 8987 12835
rect 9965 12801 9999 12835
rect 10149 12801 10183 12835
rect 3617 12733 3651 12767
rect 4169 12733 4203 12767
rect 6561 12733 6595 12767
rect 10701 12733 10735 12767
rect 5365 12665 5399 12699
rect 7158 12665 7192 12699
rect 8769 12665 8803 12699
rect 4721 12597 4755 12631
rect 7757 12597 7791 12631
rect 3111 12393 3145 12427
rect 3709 12393 3743 12427
rect 4721 12393 4755 12427
rect 6009 12393 6043 12427
rect 7757 12393 7791 12427
rect 9045 12393 9079 12427
rect 9229 12393 9263 12427
rect 9505 12393 9539 12427
rect 9781 12393 9815 12427
rect 10701 12393 10735 12427
rect 5089 12325 5123 12359
rect 6653 12325 6687 12359
rect 8217 12325 8251 12359
rect 3040 12257 3074 12291
rect 4997 12189 5031 12223
rect 5641 12189 5675 12223
rect 6561 12189 6595 12223
rect 8125 12189 8159 12223
rect 7113 12121 7147 12155
rect 8677 12121 8711 12155
rect 9965 12257 9999 12291
rect 10149 12257 10183 12291
rect 11320 12257 11354 12291
rect 11391 12121 11425 12155
rect 9229 12053 9263 12087
rect 3065 11849 3099 11883
rect 4629 11849 4663 11883
rect 4997 11849 5031 11883
rect 6561 11849 6595 11883
rect 7021 11849 7055 11883
rect 7481 11849 7515 11883
rect 8585 11849 8619 11883
rect 8861 11849 8895 11883
rect 9137 11849 9171 11883
rect 9321 11849 9355 11883
rect 11437 11849 11471 11883
rect 5181 11713 5215 11747
rect 6101 11713 6135 11747
rect 7665 11713 7699 11747
rect 3433 11645 3467 11679
rect 3801 11645 3835 11679
rect 4077 11645 4111 11679
rect 10057 11781 10091 11815
rect 9505 11713 9539 11747
rect 10793 11713 10827 11747
rect 11115 11713 11149 11747
rect 11012 11645 11046 11679
rect 4261 11577 4295 11611
rect 5273 11577 5307 11611
rect 5825 11577 5859 11611
rect 7986 11577 8020 11611
rect 9137 11577 9171 11611
rect 9597 11577 9631 11611
rect 10425 11509 10459 11543
rect 11897 11509 11931 11543
rect 3617 11305 3651 11339
rect 5181 11305 5215 11339
rect 8585 11305 8619 11339
rect 9505 11305 9539 11339
rect 4623 11237 4657 11271
rect 7618 11237 7652 11271
rect 9873 11237 9907 11271
rect 10425 11237 10459 11271
rect 11437 11237 11471 11271
rect 2421 11169 2455 11203
rect 2973 11169 3007 11203
rect 3157 11169 3191 11203
rect 6320 11169 6354 11203
rect 4261 11101 4295 11135
rect 7297 11101 7331 11135
rect 9781 11101 9815 11135
rect 11345 11101 11379 11135
rect 11621 11101 11655 11135
rect 5549 11033 5583 11067
rect 6423 11033 6457 11067
rect 8217 10965 8251 10999
rect 2881 10761 2915 10795
rect 3571 10761 3605 10795
rect 4353 10761 4387 10795
rect 5641 10761 5675 10795
rect 7389 10761 7423 10795
rect 8677 10761 8711 10795
rect 10241 10761 10275 10795
rect 10609 10761 10643 10795
rect 10931 10761 10965 10795
rect 11621 10761 11655 10795
rect 4445 10625 4479 10659
rect 9965 10625 9999 10659
rect 3500 10557 3534 10591
rect 7481 10557 7515 10591
rect 8401 10557 8435 10591
rect 10828 10557 10862 10591
rect 11253 10557 11287 10591
rect 4766 10489 4800 10523
rect 7802 10489 7836 10523
rect 9321 10489 9355 10523
rect 9413 10489 9447 10523
rect 2421 10421 2455 10455
rect 3893 10421 3927 10455
rect 5365 10421 5399 10455
rect 6285 10421 6319 10455
rect 9137 10421 9171 10455
rect 11989 10421 12023 10455
rect 3111 10217 3145 10251
rect 5089 10217 5123 10251
rect 7481 10217 7515 10251
rect 9321 10217 9355 10251
rect 9827 10217 9861 10251
rect 4721 10149 4755 10183
rect 5457 10149 5491 10183
rect 8217 10149 8251 10183
rect 8769 10149 8803 10183
rect 3040 10081 3074 10115
rect 4312 10081 4346 10115
rect 9756 10081 9790 10115
rect 4399 10013 4433 10047
rect 5365 10013 5399 10047
rect 5641 10013 5675 10047
rect 6837 10013 6871 10047
rect 8125 10013 8159 10047
rect 7849 9877 7883 9911
rect 4629 9673 4663 9707
rect 8125 9673 8159 9707
rect 4077 9605 4111 9639
rect 5825 9605 5859 9639
rect 9229 9605 9263 9639
rect 6561 9537 6595 9571
rect 7573 9537 7607 9571
rect 8539 9537 8573 9571
rect 4220 9469 4254 9503
rect 5089 9469 5123 9503
rect 6837 9469 6871 9503
rect 7389 9469 7423 9503
rect 8452 9469 8486 9503
rect 3709 9401 3743 9435
rect 4307 9401 4341 9435
rect 5273 9401 5307 9435
rect 5365 9401 5399 9435
rect 6285 9401 6319 9435
rect 8953 9401 8987 9435
rect 3065 9333 3099 9367
rect 9781 9333 9815 9367
rect 5641 9129 5675 9163
rect 6009 9129 6043 9163
rect 6469 9061 6503 9095
rect 7297 9061 7331 9095
rect 4537 8993 4571 9027
rect 4721 8993 4755 9027
rect 6561 8993 6595 9027
rect 7113 8993 7147 9027
rect 8125 8993 8159 9027
rect 4813 8925 4847 8959
rect 8309 8857 8343 8891
rect 8585 8857 8619 8891
rect 5365 8789 5399 8823
rect 7665 8789 7699 8823
rect 8953 8789 8987 8823
rect 4997 8585 5031 8619
rect 8217 8585 8251 8619
rect 4629 8517 4663 8551
rect 3525 8449 3559 8483
rect 6837 8449 6871 8483
rect 9137 8449 9171 8483
rect 3893 8381 3927 8415
rect 4169 8381 4203 8415
rect 5181 8381 5215 8415
rect 5641 8381 5675 8415
rect 6193 8381 6227 8415
rect 6653 8381 6687 8415
rect 8677 8381 8711 8415
rect 9045 8381 9079 8415
rect 4353 8313 4387 8347
rect 5917 8313 5951 8347
rect 7199 8313 7233 8347
rect 7757 8245 7791 8279
rect 3249 8041 3283 8075
rect 3709 8041 3743 8075
rect 4261 8041 4295 8075
rect 4813 8041 4847 8075
rect 7757 8041 7791 8075
rect 9781 8041 9815 8075
rect 6653 7973 6687 8007
rect 8217 7973 8251 8007
rect 4905 7905 4939 7939
rect 5365 7905 5399 7939
rect 9965 7905 9999 7939
rect 10149 7905 10183 7939
rect 5457 7837 5491 7871
rect 6561 7837 6595 7871
rect 7021 7837 7055 7871
rect 8125 7837 8159 7871
rect 8769 7837 8803 7871
rect 9505 7701 9539 7735
rect 7021 7497 7055 7531
rect 7481 7497 7515 7531
rect 8585 7497 8619 7531
rect 8861 7497 8895 7531
rect 10425 7497 10459 7531
rect 6561 7429 6595 7463
rect 4721 7361 4755 7395
rect 7665 7361 7699 7395
rect 9505 7361 9539 7395
rect 11115 7361 11149 7395
rect 3065 7293 3099 7327
rect 3433 7293 3467 7327
rect 3617 7293 3651 7327
rect 11028 7293 11062 7327
rect 11437 7293 11471 7327
rect 3893 7225 3927 7259
rect 4629 7225 4663 7259
rect 5083 7225 5117 7259
rect 7986 7225 8020 7259
rect 9597 7225 9631 7259
rect 10149 7225 10183 7259
rect 4261 7157 4295 7191
rect 5641 7157 5675 7191
rect 9229 7157 9263 7191
rect 4445 6953 4479 6987
rect 4905 6953 4939 6987
rect 9505 6953 9539 6987
rect 5594 6885 5628 6919
rect 7843 6885 7877 6919
rect 9873 6885 9907 6919
rect 2697 6817 2731 6851
rect 2973 6817 3007 6851
rect 4261 6817 4295 6851
rect 6469 6817 6503 6851
rect 7481 6817 7515 6851
rect 3157 6749 3191 6783
rect 5273 6749 5307 6783
rect 9781 6749 9815 6783
rect 10057 6749 10091 6783
rect 6193 6613 6227 6647
rect 8401 6613 8435 6647
rect 8769 6613 8803 6647
rect 2559 6409 2593 6443
rect 2973 6409 3007 6443
rect 3249 6409 3283 6443
rect 4537 6409 4571 6443
rect 6193 6409 6227 6443
rect 6653 6409 6687 6443
rect 7389 6409 7423 6443
rect 8953 6409 8987 6443
rect 9045 6409 9079 6443
rect 10609 6409 10643 6443
rect 4905 6341 4939 6375
rect 8401 6341 8435 6375
rect 2329 6273 2363 6307
rect 4997 6273 5031 6307
rect 7481 6273 7515 6307
rect 8677 6273 8711 6307
rect 2488 6205 2522 6239
rect 3433 6205 3467 6239
rect 3985 6205 4019 6239
rect 4169 6137 4203 6171
rect 5359 6137 5393 6171
rect 7802 6137 7836 6171
rect 10241 6341 10275 6375
rect 9689 6273 9723 6307
rect 9321 6137 9355 6171
rect 9413 6137 9447 6171
rect 5917 6069 5951 6103
rect 8953 6069 8987 6103
rect 2513 5865 2547 5899
rect 3525 5865 3559 5899
rect 5365 5865 5399 5899
rect 7297 5865 7331 5899
rect 8217 5865 8251 5899
rect 9827 5865 9861 5899
rect 5825 5797 5859 5831
rect 4261 5729 4295 5763
rect 4537 5729 4571 5763
rect 7205 5729 7239 5763
rect 7665 5729 7699 5763
rect 9724 5729 9758 5763
rect 4813 5661 4847 5695
rect 5733 5661 5767 5695
rect 6285 5593 6319 5627
rect 9229 5525 9263 5559
rect 4629 5321 4663 5355
rect 6193 5321 6227 5355
rect 7757 5321 7791 5355
rect 9689 5321 9723 5355
rect 6561 5253 6595 5287
rect 3525 5185 3559 5219
rect 8769 5185 8803 5219
rect 3893 5117 3927 5151
rect 4077 5117 4111 5151
rect 6837 5117 6871 5151
rect 7389 5117 7423 5151
rect 9908 5117 9942 5151
rect 10333 5117 10367 5151
rect 4353 5049 4387 5083
rect 5273 5049 5307 5083
rect 5365 5049 5399 5083
rect 5917 5049 5951 5083
rect 8401 5049 8435 5083
rect 8493 5049 8527 5083
rect 5089 4981 5123 5015
rect 7021 4981 7055 5015
rect 8217 4981 8251 5015
rect 10011 4981 10045 5015
rect 3709 4777 3743 4811
rect 4353 4777 4387 4811
rect 5917 4777 5951 4811
rect 7113 4777 7147 4811
rect 8217 4777 8251 4811
rect 5083 4709 5117 4743
rect 7618 4709 7652 4743
rect 3008 4641 3042 4675
rect 7297 4641 7331 4675
rect 9740 4641 9774 4675
rect 10736 4641 10770 4675
rect 4721 4573 4755 4607
rect 8585 4573 8619 4607
rect 9827 4573 9861 4607
rect 8953 4505 8987 4539
rect 10839 4505 10873 4539
rect 3111 4437 3145 4471
rect 5641 4437 5675 4471
rect 6285 4437 6319 4471
rect 3433 4233 3467 4267
rect 4813 4233 4847 4267
rect 8677 4233 8711 4267
rect 9965 4233 9999 4267
rect 10333 4233 10367 4267
rect 10977 4233 11011 4267
rect 3157 4165 3191 4199
rect 2743 4097 2777 4131
rect 5273 4097 5307 4131
rect 6193 4097 6227 4131
rect 6653 4097 6687 4131
rect 7113 4097 7147 4131
rect 8953 4097 8987 4131
rect 9229 4097 9263 4131
rect 1660 4029 1694 4063
rect 2656 4029 2690 4063
rect 10425 4029 10459 4063
rect 2513 3961 2547 3995
rect 3709 3961 3743 3995
rect 3801 3961 3835 3995
rect 4353 3961 4387 3995
rect 5365 3961 5399 3995
rect 5917 3961 5951 3995
rect 7434 3961 7468 3995
rect 9045 3961 9079 3995
rect 1731 3893 1765 3927
rect 2145 3893 2179 3927
rect 8033 3893 8067 3927
rect 10609 3893 10643 3927
rect 3709 3689 3743 3723
rect 5641 3689 5675 3723
rect 7205 3689 7239 3723
rect 7481 3689 7515 3723
rect 7941 3689 7975 3723
rect 10931 3689 10965 3723
rect 1869 3621 1903 3655
rect 4439 3621 4473 3655
rect 5365 3621 5399 3655
rect 6009 3621 6043 3655
rect 8217 3621 8251 3655
rect 8769 3621 8803 3655
rect 2012 3553 2046 3587
rect 4077 3553 4111 3587
rect 9689 3553 9723 3587
rect 10860 3553 10894 3587
rect 2099 3485 2133 3519
rect 2973 3485 3007 3519
rect 5917 3485 5951 3519
rect 6193 3485 6227 3519
rect 8125 3485 8159 3519
rect 2697 3349 2731 3383
rect 4997 3349 5031 3383
rect 9873 3349 9907 3383
rect 2421 3145 2455 3179
rect 5365 3145 5399 3179
rect 5917 3145 5951 3179
rect 8033 3145 8067 3179
rect 9229 3145 9263 3179
rect 10241 3145 10275 3179
rect 11621 3145 11655 3179
rect 8769 3077 8803 3111
rect 2697 3009 2731 3043
rect 3341 3009 3375 3043
rect 4169 3009 4203 3043
rect 6193 3009 6227 3043
rect 8217 3009 8251 3043
rect 9597 3009 9631 3043
rect 1660 2941 1694 2975
rect 2053 2941 2087 2975
rect 3709 2941 3743 2975
rect 4077 2941 4111 2975
rect 6837 2941 6871 2975
rect 7389 2941 7423 2975
rect 9689 2941 9723 2975
rect 10828 2941 10862 2975
rect 11253 2941 11287 2975
rect 2789 2873 2823 2907
rect 4490 2873 4524 2907
rect 8309 2873 8343 2907
rect 1731 2805 1765 2839
rect 5089 2805 5123 2839
rect 7021 2805 7055 2839
rect 9873 2805 9907 2839
rect 10931 2805 10965 2839
rect 1547 2601 1581 2635
rect 4261 2601 4295 2635
rect 4721 2601 4755 2635
rect 6653 2601 6687 2635
rect 8125 2601 8159 2635
rect 9137 2601 9171 2635
rect 12081 2601 12115 2635
rect 1961 2533 1995 2567
rect 2605 2533 2639 2567
rect 3525 2533 3559 2567
rect 4997 2533 5031 2567
rect 5089 2533 5123 2567
rect 5641 2533 5675 2567
rect 6377 2533 6411 2567
rect 7021 2533 7055 2567
rect 7113 2533 7147 2567
rect 1476 2465 1510 2499
rect 8493 2465 8527 2499
rect 10333 2465 10367 2499
rect 10885 2465 10919 2499
rect 11437 2465 11471 2499
rect 13185 2465 13219 2499
rect 13737 2465 13771 2499
rect 2329 2397 2363 2431
rect 2513 2397 2547 2431
rect 2973 2397 3007 2431
rect 5917 2397 5951 2431
rect 7297 2397 7331 2431
rect 10517 2329 10551 2363
rect 13369 2329 13403 2363
rect 8677 2261 8711 2295
rect 11621 2261 11655 2295
<< metal1 >>
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 4062 37272 4068 37324
rect 4120 37312 4126 37324
rect 5994 37312 6000 37324
rect 4120 37284 6000 37312
rect 4120 37272 4126 37284
rect 5994 37272 6000 37284
rect 6052 37272 6058 37324
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 9652 36703 9710 36709
rect 9652 36669 9664 36703
rect 9698 36700 9710 36703
rect 9698 36672 10180 36700
rect 9698 36669 9710 36672
rect 9652 36663 9710 36669
rect 9723 36567 9781 36573
rect 9723 36533 9735 36567
rect 9769 36564 9781 36567
rect 9950 36564 9956 36576
rect 9769 36536 9956 36564
rect 9769 36533 9781 36536
rect 9723 36527 9781 36533
rect 9950 36524 9956 36536
rect 10008 36524 10014 36576
rect 10152 36573 10180 36672
rect 10137 36567 10195 36573
rect 10137 36533 10149 36567
rect 10183 36564 10195 36567
rect 10686 36564 10692 36576
rect 10183 36536 10692 36564
rect 10183 36533 10195 36536
rect 10137 36527 10195 36533
rect 10686 36524 10692 36536
rect 10744 36524 10750 36576
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 8665 36363 8723 36369
rect 8665 36329 8677 36363
rect 8711 36360 8723 36363
rect 9306 36360 9312 36372
rect 8711 36332 9312 36360
rect 8711 36329 8723 36332
rect 8665 36323 8723 36329
rect 9306 36320 9312 36332
rect 9364 36320 9370 36372
rect 8297 36295 8355 36301
rect 8297 36261 8309 36295
rect 8343 36292 8355 36295
rect 8570 36292 8576 36304
rect 8343 36264 8576 36292
rect 8343 36261 8355 36264
rect 8297 36255 8355 36261
rect 8570 36252 8576 36264
rect 8628 36252 8634 36304
rect 7466 36184 7472 36236
rect 7524 36233 7530 36236
rect 7524 36227 7562 36233
rect 7550 36193 7562 36227
rect 7524 36187 7562 36193
rect 8481 36227 8539 36233
rect 8481 36193 8493 36227
rect 8527 36224 8539 36227
rect 9582 36224 9588 36236
rect 8527 36196 9588 36224
rect 8527 36193 8539 36196
rect 8481 36187 8539 36193
rect 7524 36184 7530 36187
rect 9582 36184 9588 36196
rect 9640 36184 9646 36236
rect 9766 36233 9772 36236
rect 9744 36227 9772 36233
rect 9744 36193 9756 36227
rect 9744 36187 9772 36193
rect 9766 36184 9772 36187
rect 9824 36184 9830 36236
rect 7607 36091 7665 36097
rect 7607 36057 7619 36091
rect 7653 36088 7665 36091
rect 8294 36088 8300 36100
rect 7653 36060 8300 36088
rect 7653 36057 7665 36060
rect 7607 36051 7665 36057
rect 8294 36048 8300 36060
rect 8352 36048 8358 36100
rect 9815 36023 9873 36029
rect 9815 35989 9827 36023
rect 9861 36020 9873 36023
rect 10229 36023 10287 36029
rect 10229 36020 10241 36023
rect 9861 35992 10241 36020
rect 9861 35989 9873 35992
rect 9815 35983 9873 35989
rect 10229 35989 10241 35992
rect 10275 36020 10287 36023
rect 10318 36020 10324 36032
rect 10275 35992 10324 36020
rect 10275 35989 10287 35992
rect 10229 35983 10287 35989
rect 10318 35980 10324 35992
rect 10376 35980 10382 36032
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 7466 35776 7472 35828
rect 7524 35816 7530 35828
rect 7745 35819 7803 35825
rect 7745 35816 7757 35819
rect 7524 35788 7757 35816
rect 7524 35776 7530 35788
rect 7745 35785 7757 35788
rect 7791 35785 7803 35819
rect 7745 35779 7803 35785
rect 9309 35819 9367 35825
rect 9309 35785 9321 35819
rect 9355 35816 9367 35819
rect 9582 35816 9588 35828
rect 9355 35788 9588 35816
rect 9355 35785 9367 35788
rect 9309 35779 9367 35785
rect 9582 35776 9588 35788
rect 9640 35776 9646 35828
rect 7006 35748 7012 35760
rect 6967 35720 7012 35748
rect 7006 35708 7012 35720
rect 7064 35708 7070 35760
rect 8754 35680 8760 35692
rect 8715 35652 8760 35680
rect 8754 35640 8760 35652
rect 8812 35640 8818 35692
rect 10318 35680 10324 35692
rect 10279 35652 10324 35680
rect 10318 35640 10324 35652
rect 10376 35640 10382 35692
rect 10778 35680 10784 35692
rect 10739 35652 10784 35680
rect 10778 35640 10784 35652
rect 10836 35640 10842 35692
rect 5626 35572 5632 35624
rect 5684 35612 5690 35624
rect 6825 35615 6883 35621
rect 6825 35612 6837 35615
rect 5684 35584 6837 35612
rect 5684 35572 5690 35584
rect 6825 35581 6837 35584
rect 6871 35612 6883 35615
rect 7377 35615 7435 35621
rect 7377 35612 7389 35615
rect 6871 35584 7389 35612
rect 6871 35581 6883 35584
rect 6825 35575 6883 35581
rect 7377 35581 7389 35584
rect 7423 35581 7435 35615
rect 7377 35575 7435 35581
rect 8294 35544 8300 35556
rect 8255 35516 8300 35544
rect 8294 35504 8300 35516
rect 8352 35504 8358 35556
rect 8389 35547 8447 35553
rect 8389 35513 8401 35547
rect 8435 35544 8447 35547
rect 8570 35544 8576 35556
rect 8435 35516 8576 35544
rect 8435 35513 8447 35516
rect 8389 35507 8447 35513
rect 8570 35504 8576 35516
rect 8628 35504 8634 35556
rect 10137 35547 10195 35553
rect 10137 35513 10149 35547
rect 10183 35544 10195 35547
rect 10410 35544 10416 35556
rect 10183 35516 10416 35544
rect 10183 35513 10195 35516
rect 10137 35507 10195 35513
rect 10410 35504 10416 35516
rect 10468 35504 10474 35556
rect 9766 35476 9772 35488
rect 9727 35448 9772 35476
rect 9766 35436 9772 35448
rect 9824 35436 9830 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 5994 35232 6000 35284
rect 6052 35281 6058 35284
rect 6052 35275 6101 35281
rect 6052 35241 6055 35275
rect 6089 35241 6101 35275
rect 6052 35235 6101 35241
rect 6052 35232 6058 35235
rect 8294 35232 8300 35284
rect 8352 35272 8358 35284
rect 9033 35275 9091 35281
rect 9033 35272 9045 35275
rect 8352 35244 9045 35272
rect 8352 35232 8358 35244
rect 9033 35241 9045 35244
rect 9079 35241 9091 35275
rect 9033 35235 9091 35241
rect 9950 35232 9956 35284
rect 10008 35272 10014 35284
rect 10229 35275 10287 35281
rect 10229 35272 10241 35275
rect 10008 35244 10241 35272
rect 10008 35232 10014 35244
rect 10229 35241 10241 35244
rect 10275 35241 10287 35275
rect 13170 35272 13176 35284
rect 13131 35244 13176 35272
rect 10229 35235 10287 35241
rect 13170 35232 13176 35244
rect 13228 35232 13234 35284
rect 8205 35207 8263 35213
rect 8205 35173 8217 35207
rect 8251 35204 8263 35207
rect 8570 35204 8576 35216
rect 8251 35176 8576 35204
rect 8251 35173 8263 35176
rect 8205 35167 8263 35173
rect 8570 35164 8576 35176
rect 8628 35164 8634 35216
rect 10594 35204 10600 35216
rect 10555 35176 10600 35204
rect 10594 35164 10600 35176
rect 10652 35164 10658 35216
rect 5972 35139 6030 35145
rect 5972 35105 5984 35139
rect 6018 35136 6030 35139
rect 6730 35136 6736 35148
rect 6018 35108 6736 35136
rect 6018 35105 6030 35108
rect 5972 35099 6030 35105
rect 6730 35096 6736 35108
rect 6788 35096 6794 35148
rect 6917 35139 6975 35145
rect 6917 35105 6929 35139
rect 6963 35136 6975 35139
rect 7282 35136 7288 35148
rect 6963 35108 7288 35136
rect 6963 35105 6975 35108
rect 6917 35099 6975 35105
rect 7282 35096 7288 35108
rect 7340 35096 7346 35148
rect 12066 35145 12072 35148
rect 12044 35139 12072 35145
rect 12044 35105 12056 35139
rect 12044 35099 12072 35105
rect 12066 35096 12072 35099
rect 12124 35096 12130 35148
rect 12989 35139 13047 35145
rect 12989 35105 13001 35139
rect 13035 35136 13047 35139
rect 13078 35136 13084 35148
rect 13035 35108 13084 35136
rect 13035 35105 13047 35108
rect 12989 35099 13047 35105
rect 13078 35096 13084 35108
rect 13136 35096 13142 35148
rect 8110 35068 8116 35080
rect 8071 35040 8116 35068
rect 8110 35028 8116 35040
rect 8168 35028 8174 35080
rect 8389 35071 8447 35077
rect 8389 35037 8401 35071
rect 8435 35037 8447 35071
rect 8389 35031 8447 35037
rect 10505 35071 10563 35077
rect 10505 35037 10517 35071
rect 10551 35068 10563 35071
rect 10962 35068 10968 35080
rect 10551 35040 10968 35068
rect 10551 35037 10563 35040
rect 10505 35031 10563 35037
rect 7101 35003 7159 35009
rect 7101 34969 7113 35003
rect 7147 35000 7159 35003
rect 8202 35000 8208 35012
rect 7147 34972 8208 35000
rect 7147 34969 7159 34972
rect 7101 34963 7159 34969
rect 8202 34960 8208 34972
rect 8260 34960 8266 35012
rect 7558 34932 7564 34944
rect 7519 34904 7564 34932
rect 7558 34892 7564 34904
rect 7616 34892 7622 34944
rect 8018 34892 8024 34944
rect 8076 34932 8082 34944
rect 8404 34932 8432 35031
rect 10962 35028 10968 35040
rect 11020 35028 11026 35080
rect 11149 35071 11207 35077
rect 11149 35037 11161 35071
rect 11195 35068 11207 35071
rect 11514 35068 11520 35080
rect 11195 35040 11520 35068
rect 11195 35037 11207 35040
rect 11149 35031 11207 35037
rect 11514 35028 11520 35040
rect 11572 35028 11578 35080
rect 8076 34904 8432 34932
rect 12115 34935 12173 34941
rect 8076 34892 8082 34904
rect 12115 34901 12127 34935
rect 12161 34932 12173 34935
rect 12526 34932 12532 34944
rect 12161 34904 12532 34932
rect 12161 34901 12173 34904
rect 12115 34895 12173 34901
rect 12526 34892 12532 34904
rect 12584 34892 12590 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 8110 34688 8116 34740
rect 8168 34728 8174 34740
rect 8941 34731 8999 34737
rect 8941 34728 8953 34731
rect 8168 34700 8953 34728
rect 8168 34688 8174 34700
rect 8941 34697 8953 34700
rect 8987 34697 8999 34731
rect 8941 34691 8999 34697
rect 9309 34731 9367 34737
rect 9309 34697 9321 34731
rect 9355 34728 9367 34731
rect 10134 34728 10140 34740
rect 9355 34700 10140 34728
rect 9355 34697 9367 34700
rect 9309 34691 9367 34697
rect 10134 34688 10140 34700
rect 10192 34688 10198 34740
rect 11054 34688 11060 34740
rect 11112 34728 11118 34740
rect 12621 34731 12679 34737
rect 12621 34728 12633 34731
rect 11112 34700 12633 34728
rect 11112 34688 11118 34700
rect 12621 34697 12633 34700
rect 12667 34697 12679 34731
rect 12621 34691 12679 34697
rect 5810 34660 5816 34672
rect 5771 34632 5816 34660
rect 5810 34620 5816 34632
rect 5868 34620 5874 34672
rect 7558 34620 7564 34672
rect 7616 34660 7622 34672
rect 7616 34632 7696 34660
rect 7616 34620 7622 34632
rect 7668 34601 7696 34632
rect 7653 34595 7711 34601
rect 7653 34561 7665 34595
rect 7699 34561 7711 34595
rect 8018 34592 8024 34604
rect 7979 34564 8024 34592
rect 7653 34555 7711 34561
rect 8018 34552 8024 34564
rect 8076 34552 8082 34604
rect 9950 34552 9956 34604
rect 10008 34592 10014 34604
rect 10321 34595 10379 34601
rect 10321 34592 10333 34595
rect 10008 34564 10333 34592
rect 10008 34552 10014 34564
rect 10321 34561 10333 34564
rect 10367 34561 10379 34595
rect 10778 34592 10784 34604
rect 10739 34564 10784 34592
rect 10321 34555 10379 34561
rect 10778 34552 10784 34564
rect 10836 34552 10842 34604
rect 5534 34484 5540 34536
rect 5592 34524 5598 34536
rect 5629 34527 5687 34533
rect 5629 34524 5641 34527
rect 5592 34496 5641 34524
rect 5592 34484 5598 34496
rect 5629 34493 5641 34496
rect 5675 34524 5687 34527
rect 6181 34527 6239 34533
rect 6181 34524 6193 34527
rect 5675 34496 6193 34524
rect 5675 34493 5687 34496
rect 5629 34487 5687 34493
rect 6181 34493 6193 34496
rect 6227 34493 6239 34527
rect 6181 34487 6239 34493
rect 6641 34527 6699 34533
rect 6641 34493 6653 34527
rect 6687 34524 6699 34527
rect 6730 34524 6736 34536
rect 6687 34496 6736 34524
rect 6687 34493 6699 34496
rect 6641 34487 6699 34493
rect 6730 34484 6736 34496
rect 6788 34484 6794 34536
rect 8662 34524 8668 34536
rect 8623 34496 8668 34524
rect 8662 34484 8668 34496
rect 8720 34484 8726 34536
rect 8846 34484 8852 34536
rect 8904 34524 8910 34536
rect 9125 34527 9183 34533
rect 9125 34524 9137 34527
rect 8904 34496 9137 34524
rect 8904 34484 8910 34496
rect 9125 34493 9137 34496
rect 9171 34524 9183 34527
rect 9677 34527 9735 34533
rect 9677 34524 9689 34527
rect 9171 34496 9689 34524
rect 9171 34493 9183 34496
rect 9125 34487 9183 34493
rect 9677 34493 9689 34496
rect 9723 34493 9735 34527
rect 12066 34524 12072 34536
rect 12027 34496 12072 34524
rect 9677 34487 9735 34493
rect 12066 34484 12072 34496
rect 12124 34484 12130 34536
rect 12434 34524 12440 34536
rect 12395 34496 12440 34524
rect 12434 34484 12440 34496
rect 12492 34524 12498 34536
rect 12989 34527 13047 34533
rect 12989 34524 13001 34527
rect 12492 34496 13001 34524
rect 12492 34484 12498 34496
rect 12989 34493 13001 34496
rect 13035 34493 13047 34527
rect 12989 34487 13047 34493
rect 13078 34484 13084 34536
rect 13136 34524 13142 34536
rect 13357 34527 13415 34533
rect 13357 34524 13369 34527
rect 13136 34496 13369 34524
rect 13136 34484 13142 34496
rect 13357 34493 13369 34496
rect 13403 34493 13415 34527
rect 13357 34487 13415 34493
rect 7469 34459 7527 34465
rect 7469 34425 7481 34459
rect 7515 34456 7527 34459
rect 7745 34459 7803 34465
rect 7745 34456 7757 34459
rect 7515 34428 7757 34456
rect 7515 34425 7527 34428
rect 7469 34419 7527 34425
rect 7745 34425 7757 34428
rect 7791 34456 7803 34459
rect 7926 34456 7932 34468
rect 7791 34428 7932 34456
rect 7791 34425 7803 34428
rect 7745 34419 7803 34425
rect 7926 34416 7932 34428
rect 7984 34416 7990 34468
rect 10413 34459 10471 34465
rect 10413 34425 10425 34459
rect 10459 34425 10471 34459
rect 10413 34419 10471 34425
rect 7101 34391 7159 34397
rect 7101 34357 7113 34391
rect 7147 34388 7159 34391
rect 7282 34388 7288 34400
rect 7147 34360 7288 34388
rect 7147 34357 7159 34360
rect 7101 34351 7159 34357
rect 7282 34348 7288 34360
rect 7340 34348 7346 34400
rect 10137 34391 10195 34397
rect 10137 34357 10149 34391
rect 10183 34388 10195 34391
rect 10226 34388 10232 34400
rect 10183 34360 10232 34388
rect 10183 34357 10195 34360
rect 10137 34351 10195 34357
rect 10226 34348 10232 34360
rect 10284 34388 10290 34400
rect 10428 34388 10456 34419
rect 10594 34388 10600 34400
rect 10284 34360 10600 34388
rect 10284 34348 10290 34360
rect 10594 34348 10600 34360
rect 10652 34388 10658 34400
rect 11241 34391 11299 34397
rect 11241 34388 11253 34391
rect 10652 34360 11253 34388
rect 10652 34348 10658 34360
rect 11241 34357 11253 34360
rect 11287 34357 11299 34391
rect 11241 34351 11299 34357
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 5350 34193 5356 34196
rect 5307 34187 5356 34193
rect 5307 34153 5319 34187
rect 5353 34153 5356 34187
rect 5307 34147 5356 34153
rect 5350 34144 5356 34147
rect 5408 34144 5414 34196
rect 13170 34184 13176 34196
rect 13131 34156 13176 34184
rect 13170 34144 13176 34156
rect 13228 34144 13234 34196
rect 6362 34116 6368 34128
rect 6323 34088 6368 34116
rect 6362 34076 6368 34088
rect 6420 34076 6426 34128
rect 7926 34116 7932 34128
rect 7887 34088 7932 34116
rect 7926 34076 7932 34088
rect 7984 34076 7990 34128
rect 10042 34125 10048 34128
rect 10039 34116 10048 34125
rect 10003 34088 10048 34116
rect 10039 34079 10048 34088
rect 10042 34076 10048 34079
rect 10100 34076 10106 34128
rect 11054 34116 11060 34128
rect 10612 34088 11060 34116
rect 5258 34057 5264 34060
rect 5236 34051 5264 34057
rect 5236 34017 5248 34051
rect 5236 34011 5264 34017
rect 5258 34008 5264 34011
rect 5316 34008 5322 34060
rect 10612 34057 10640 34088
rect 11054 34076 11060 34088
rect 11112 34116 11118 34128
rect 11609 34119 11667 34125
rect 11609 34116 11621 34119
rect 11112 34088 11621 34116
rect 11112 34076 11118 34088
rect 11609 34085 11621 34088
rect 11655 34085 11667 34119
rect 11609 34079 11667 34085
rect 10597 34051 10655 34057
rect 10597 34017 10609 34051
rect 10643 34017 10655 34051
rect 10597 34011 10655 34017
rect 12158 34008 12164 34060
rect 12216 34048 12222 34060
rect 12989 34051 13047 34057
rect 12989 34048 13001 34051
rect 12216 34020 13001 34048
rect 12216 34008 12222 34020
rect 12989 34017 13001 34020
rect 13035 34048 13047 34051
rect 13446 34048 13452 34060
rect 13035 34020 13452 34048
rect 13035 34017 13047 34020
rect 12989 34011 13047 34017
rect 13446 34008 13452 34020
rect 13504 34008 13510 34060
rect 6273 33983 6331 33989
rect 6273 33949 6285 33983
rect 6319 33949 6331 33983
rect 6273 33943 6331 33949
rect 7837 33983 7895 33989
rect 7837 33949 7849 33983
rect 7883 33980 7895 33983
rect 8294 33980 8300 33992
rect 7883 33952 8300 33980
rect 7883 33949 7895 33952
rect 7837 33943 7895 33949
rect 6178 33872 6184 33924
rect 6236 33912 6242 33924
rect 6288 33912 6316 33943
rect 8294 33940 8300 33952
rect 8352 33940 8358 33992
rect 8481 33983 8539 33989
rect 8481 33949 8493 33983
rect 8527 33980 8539 33983
rect 8754 33980 8760 33992
rect 8527 33952 8760 33980
rect 8527 33949 8539 33952
rect 8481 33943 8539 33949
rect 6236 33884 6316 33912
rect 6825 33915 6883 33921
rect 6236 33872 6242 33884
rect 6825 33881 6837 33915
rect 6871 33912 6883 33915
rect 8496 33912 8524 33943
rect 8754 33940 8760 33952
rect 8812 33980 8818 33992
rect 9490 33980 9496 33992
rect 8812 33952 9496 33980
rect 8812 33940 8818 33952
rect 9490 33940 9496 33952
rect 9548 33940 9554 33992
rect 9674 33980 9680 33992
rect 9635 33952 9680 33980
rect 9674 33940 9680 33952
rect 9732 33940 9738 33992
rect 11330 33940 11336 33992
rect 11388 33980 11394 33992
rect 11517 33983 11575 33989
rect 11517 33980 11529 33983
rect 11388 33952 11529 33980
rect 11388 33940 11394 33952
rect 11517 33949 11529 33952
rect 11563 33949 11575 33983
rect 11517 33943 11575 33949
rect 11793 33983 11851 33989
rect 11793 33949 11805 33983
rect 11839 33949 11851 33983
rect 11793 33943 11851 33949
rect 6871 33884 8524 33912
rect 6871 33881 6883 33884
rect 6825 33875 6883 33881
rect 10778 33872 10784 33924
rect 10836 33912 10842 33924
rect 11808 33912 11836 33943
rect 10836 33884 11836 33912
rect 10836 33872 10842 33884
rect 7558 33844 7564 33856
rect 7519 33816 7564 33844
rect 7558 33804 7564 33816
rect 7616 33804 7622 33856
rect 10962 33844 10968 33856
rect 10923 33816 10968 33844
rect 10962 33804 10968 33816
rect 11020 33804 11026 33856
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 4890 33649 4896 33652
rect 4847 33643 4896 33649
rect 4847 33609 4859 33643
rect 4893 33609 4896 33643
rect 4847 33603 4896 33609
rect 4890 33600 4896 33603
rect 4948 33600 4954 33652
rect 6362 33600 6368 33652
rect 6420 33640 6426 33652
rect 6549 33643 6607 33649
rect 6549 33640 6561 33643
rect 6420 33612 6561 33640
rect 6420 33600 6426 33612
rect 6549 33609 6561 33612
rect 6595 33640 6607 33643
rect 7193 33643 7251 33649
rect 7193 33640 7205 33643
rect 6595 33612 7205 33640
rect 6595 33609 6607 33612
rect 6549 33603 6607 33609
rect 7193 33609 7205 33612
rect 7239 33640 7251 33643
rect 7285 33643 7343 33649
rect 7285 33640 7297 33643
rect 7239 33612 7297 33640
rect 7239 33609 7251 33612
rect 7193 33603 7251 33609
rect 7285 33609 7297 33612
rect 7331 33609 7343 33643
rect 10226 33640 10232 33652
rect 10187 33612 10232 33640
rect 7285 33603 7343 33609
rect 10226 33600 10232 33612
rect 10284 33600 10290 33652
rect 11241 33643 11299 33649
rect 11241 33609 11253 33643
rect 11287 33640 11299 33643
rect 11974 33640 11980 33652
rect 11287 33612 11980 33640
rect 11287 33609 11299 33612
rect 11241 33603 11299 33609
rect 11974 33600 11980 33612
rect 12032 33600 12038 33652
rect 13446 33640 13452 33652
rect 13407 33612 13452 33640
rect 13446 33600 13452 33612
rect 13504 33600 13510 33652
rect 5859 33575 5917 33581
rect 5859 33541 5871 33575
rect 5905 33572 5917 33575
rect 5905 33544 6408 33572
rect 5905 33541 5917 33544
rect 5859 33535 5917 33541
rect 6380 33504 6408 33544
rect 7558 33504 7564 33516
rect 6380 33476 7564 33504
rect 7558 33464 7564 33476
rect 7616 33464 7622 33516
rect 8018 33504 8024 33516
rect 7979 33476 8024 33504
rect 8018 33464 8024 33476
rect 8076 33464 8082 33516
rect 8849 33507 8907 33513
rect 8849 33473 8861 33507
rect 8895 33504 8907 33507
rect 9674 33504 9680 33516
rect 8895 33476 9680 33504
rect 8895 33473 8907 33476
rect 8849 33467 8907 33473
rect 9674 33464 9680 33476
rect 9732 33464 9738 33516
rect 12526 33504 12532 33516
rect 12487 33476 12532 33504
rect 12526 33464 12532 33476
rect 12584 33464 12590 33516
rect 12802 33504 12808 33516
rect 12763 33476 12808 33504
rect 12802 33464 12808 33476
rect 12860 33464 12866 33516
rect 4706 33396 4712 33448
rect 4764 33445 4770 33448
rect 4764 33439 4802 33445
rect 4790 33405 4802 33439
rect 5258 33436 5264 33448
rect 5219 33408 5264 33436
rect 4764 33399 4802 33405
rect 4764 33396 4770 33399
rect 5258 33396 5264 33408
rect 5316 33396 5322 33448
rect 5788 33439 5846 33445
rect 5788 33405 5800 33439
rect 5834 33436 5846 33439
rect 9306 33436 9312 33448
rect 5834 33408 6316 33436
rect 9267 33408 9312 33436
rect 5834 33405 5846 33408
rect 5788 33399 5846 33405
rect 4724 33368 4752 33396
rect 5537 33371 5595 33377
rect 5537 33368 5549 33371
rect 4724 33340 5549 33368
rect 5537 33337 5549 33340
rect 5583 33368 5595 33371
rect 6086 33368 6092 33380
rect 5583 33340 6092 33368
rect 5583 33337 5595 33340
rect 5537 33331 5595 33337
rect 6086 33328 6092 33340
rect 6144 33328 6150 33380
rect 6288 33309 6316 33408
rect 9306 33396 9312 33408
rect 9364 33396 9370 33448
rect 11057 33439 11115 33445
rect 11057 33405 11069 33439
rect 11103 33436 11115 33439
rect 11146 33436 11152 33448
rect 11103 33408 11152 33436
rect 11103 33405 11115 33408
rect 11057 33399 11115 33405
rect 11146 33396 11152 33408
rect 11204 33436 11210 33448
rect 11609 33439 11667 33445
rect 11609 33436 11621 33439
rect 11204 33408 11621 33436
rect 11204 33396 11210 33408
rect 11609 33405 11621 33408
rect 11655 33436 11667 33439
rect 12250 33436 12256 33448
rect 11655 33408 12256 33436
rect 11655 33405 11667 33408
rect 11609 33399 11667 33405
rect 12250 33396 12256 33408
rect 12308 33396 12314 33448
rect 7193 33371 7251 33377
rect 7193 33337 7205 33371
rect 7239 33368 7251 33371
rect 7650 33368 7656 33380
rect 7239 33340 7656 33368
rect 7239 33337 7251 33340
rect 7193 33331 7251 33337
rect 7650 33328 7656 33340
rect 7708 33328 7714 33380
rect 9671 33371 9729 33377
rect 9671 33337 9683 33371
rect 9717 33337 9729 33371
rect 9671 33331 9729 33337
rect 6273 33303 6331 33309
rect 6273 33269 6285 33303
rect 6319 33300 6331 33303
rect 7282 33300 7288 33312
rect 6319 33272 7288 33300
rect 6319 33269 6331 33272
rect 6273 33263 6331 33269
rect 7282 33260 7288 33272
rect 7340 33260 7346 33312
rect 9217 33303 9275 33309
rect 9217 33269 9229 33303
rect 9263 33300 9275 33303
rect 9398 33300 9404 33312
rect 9263 33272 9404 33300
rect 9263 33269 9275 33272
rect 9217 33263 9275 33269
rect 9398 33260 9404 33272
rect 9456 33300 9462 33312
rect 9692 33300 9720 33331
rect 10870 33328 10876 33380
rect 10928 33368 10934 33380
rect 12161 33371 12219 33377
rect 12161 33368 12173 33371
rect 10928 33340 12173 33368
rect 10928 33328 10934 33340
rect 12161 33337 12173 33340
rect 12207 33368 12219 33371
rect 12621 33371 12679 33377
rect 12621 33368 12633 33371
rect 12207 33340 12633 33368
rect 12207 33337 12219 33340
rect 12161 33331 12219 33337
rect 12621 33337 12633 33340
rect 12667 33337 12679 33371
rect 12621 33331 12679 33337
rect 10042 33300 10048 33312
rect 9456 33272 10048 33300
rect 9456 33260 9462 33272
rect 10042 33260 10048 33272
rect 10100 33300 10106 33312
rect 10505 33303 10563 33309
rect 10505 33300 10517 33303
rect 10100 33272 10517 33300
rect 10100 33260 10106 33272
rect 10505 33269 10517 33272
rect 10551 33269 10563 33303
rect 10505 33263 10563 33269
rect 10965 33303 11023 33309
rect 10965 33269 10977 33303
rect 11011 33300 11023 33303
rect 11054 33300 11060 33312
rect 11011 33272 11060 33300
rect 11011 33269 11023 33272
rect 10965 33263 11023 33269
rect 11054 33260 11060 33272
rect 11112 33260 11118 33312
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 5859 33099 5917 33105
rect 5859 33065 5871 33099
rect 5905 33096 5917 33099
rect 6178 33096 6184 33108
rect 5905 33068 6184 33096
rect 5905 33065 5917 33068
rect 5859 33059 5917 33065
rect 6178 33056 6184 33068
rect 6236 33056 6242 33108
rect 7650 33096 7656 33108
rect 7611 33068 7656 33096
rect 7650 33056 7656 33068
rect 7708 33056 7714 33108
rect 7926 33096 7932 33108
rect 7887 33068 7932 33096
rect 7926 33056 7932 33068
rect 7984 33056 7990 33108
rect 8294 33096 8300 33108
rect 8255 33068 8300 33096
rect 8294 33056 8300 33068
rect 8352 33096 8358 33108
rect 8619 33099 8677 33105
rect 8619 33096 8631 33099
rect 8352 33068 8631 33096
rect 8352 33056 8358 33068
rect 8619 33065 8631 33068
rect 8665 33065 8677 33099
rect 8619 33059 8677 33065
rect 10410 33056 10416 33108
rect 10468 33096 10474 33108
rect 10597 33099 10655 33105
rect 10597 33096 10609 33099
rect 10468 33068 10609 33096
rect 10468 33056 10474 33068
rect 10597 33065 10609 33068
rect 10643 33096 10655 33099
rect 10870 33096 10876 33108
rect 10643 33068 10876 33096
rect 10643 33065 10655 33068
rect 10597 33059 10655 33065
rect 10870 33056 10876 33068
rect 10928 33056 10934 33108
rect 12526 33096 12532 33108
rect 12487 33068 12532 33096
rect 12526 33056 12532 33068
rect 12584 33056 12590 33108
rect 7095 33031 7153 33037
rect 7095 32997 7107 33031
rect 7141 33028 7153 33031
rect 7190 33028 7196 33040
rect 7141 33000 7196 33028
rect 7141 32997 7153 33000
rect 7095 32991 7153 32997
rect 7190 32988 7196 33000
rect 7248 32988 7254 33040
rect 9398 32988 9404 33040
rect 9456 33028 9462 33040
rect 9998 33031 10056 33037
rect 9998 33028 10010 33031
rect 9456 33000 10010 33028
rect 9456 32988 9462 33000
rect 9998 32997 10010 33000
rect 10044 32997 10056 33031
rect 9998 32991 10056 32997
rect 11054 32988 11060 33040
rect 11112 33028 11118 33040
rect 11609 33031 11667 33037
rect 11609 33028 11621 33031
rect 11112 33000 11621 33028
rect 11112 32988 11118 33000
rect 11609 32997 11621 33000
rect 11655 33028 11667 33031
rect 11698 33028 11704 33040
rect 11655 33000 11704 33028
rect 11655 32997 11667 33000
rect 11609 32991 11667 32997
rect 11698 32988 11704 33000
rect 11756 32988 11762 33040
rect 5788 32963 5846 32969
rect 5788 32929 5800 32963
rect 5834 32960 5846 32963
rect 5994 32960 6000 32972
rect 5834 32932 6000 32960
rect 5834 32929 5846 32932
rect 5788 32923 5846 32929
rect 5994 32920 6000 32932
rect 6052 32920 6058 32972
rect 8570 32969 8576 32972
rect 8548 32963 8576 32969
rect 8548 32929 8560 32963
rect 8548 32923 8576 32929
rect 8570 32920 8576 32923
rect 8628 32920 8634 32972
rect 13078 32969 13084 32972
rect 13056 32963 13084 32969
rect 13056 32929 13068 32963
rect 13056 32923 13084 32929
rect 13078 32920 13084 32923
rect 13136 32920 13142 32972
rect 6733 32895 6791 32901
rect 6733 32861 6745 32895
rect 6779 32892 6791 32895
rect 7466 32892 7472 32904
rect 6779 32864 7472 32892
rect 6779 32861 6791 32864
rect 6733 32855 6791 32861
rect 7466 32852 7472 32864
rect 7524 32852 7530 32904
rect 9677 32895 9735 32901
rect 9677 32861 9689 32895
rect 9723 32892 9735 32895
rect 10410 32892 10416 32904
rect 9723 32864 10416 32892
rect 9723 32861 9735 32864
rect 9677 32855 9735 32861
rect 10410 32852 10416 32864
rect 10468 32852 10474 32904
rect 11514 32892 11520 32904
rect 11475 32864 11520 32892
rect 11514 32852 11520 32864
rect 11572 32852 11578 32904
rect 11606 32852 11612 32904
rect 11664 32892 11670 32904
rect 11793 32895 11851 32901
rect 11793 32892 11805 32895
rect 11664 32864 11805 32892
rect 11664 32852 11670 32864
rect 11793 32861 11805 32864
rect 11839 32861 11851 32895
rect 11793 32855 11851 32861
rect 8754 32716 8760 32768
rect 8812 32756 8818 32768
rect 8941 32759 8999 32765
rect 8941 32756 8953 32759
rect 8812 32728 8953 32756
rect 8812 32716 8818 32728
rect 8941 32725 8953 32728
rect 8987 32725 8999 32759
rect 9306 32756 9312 32768
rect 9267 32728 9312 32756
rect 8941 32719 8999 32725
rect 9306 32716 9312 32728
rect 9364 32716 9370 32768
rect 11330 32756 11336 32768
rect 11243 32728 11336 32756
rect 11330 32716 11336 32728
rect 11388 32756 11394 32768
rect 13127 32759 13185 32765
rect 13127 32756 13139 32759
rect 11388 32728 13139 32756
rect 11388 32716 11394 32728
rect 13127 32725 13139 32728
rect 13173 32725 13185 32759
rect 13127 32719 13185 32725
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 7745 32555 7803 32561
rect 7745 32521 7757 32555
rect 7791 32552 7803 32555
rect 7926 32552 7932 32564
rect 7791 32524 7932 32552
rect 7791 32521 7803 32524
rect 7745 32515 7803 32521
rect 7926 32512 7932 32524
rect 7984 32512 7990 32564
rect 8570 32512 8576 32564
rect 8628 32512 8634 32564
rect 8662 32512 8668 32564
rect 8720 32552 8726 32564
rect 9493 32555 9551 32561
rect 9493 32552 9505 32555
rect 8720 32524 9505 32552
rect 8720 32512 8726 32524
rect 9493 32521 9505 32524
rect 9539 32521 9551 32555
rect 11698 32552 11704 32564
rect 11659 32524 11704 32552
rect 9493 32515 9551 32521
rect 11698 32512 11704 32524
rect 11756 32512 11762 32564
rect 12434 32512 12440 32564
rect 12492 32552 12498 32564
rect 12575 32555 12633 32561
rect 12575 32552 12587 32555
rect 12492 32524 12587 32552
rect 12492 32512 12498 32524
rect 12575 32521 12587 32524
rect 12621 32521 12633 32555
rect 12575 32515 12633 32521
rect 8481 32487 8539 32493
rect 8481 32453 8493 32487
rect 8527 32484 8539 32487
rect 8588 32484 8616 32512
rect 8938 32484 8944 32496
rect 8527 32456 8944 32484
rect 8527 32453 8539 32456
rect 8481 32447 8539 32453
rect 8938 32444 8944 32456
rect 8996 32444 9002 32496
rect 8573 32419 8631 32425
rect 8573 32385 8585 32419
rect 8619 32416 8631 32419
rect 8754 32416 8760 32428
rect 8619 32388 8760 32416
rect 8619 32385 8631 32388
rect 8573 32379 8631 32385
rect 8754 32376 8760 32388
rect 8812 32376 8818 32428
rect 6822 32348 6828 32360
rect 6783 32320 6828 32348
rect 6822 32308 6828 32320
rect 6880 32308 6886 32360
rect 10597 32351 10655 32357
rect 10597 32317 10609 32351
rect 10643 32348 10655 32351
rect 10686 32348 10692 32360
rect 10643 32320 10692 32348
rect 10643 32317 10655 32320
rect 10597 32311 10655 32317
rect 10686 32308 10692 32320
rect 10744 32308 10750 32360
rect 10781 32351 10839 32357
rect 10781 32317 10793 32351
rect 10827 32317 10839 32351
rect 12472 32351 12530 32357
rect 12472 32348 12484 32351
rect 10781 32311 10839 32317
rect 12176 32320 12484 32348
rect 7190 32289 7196 32292
rect 7187 32280 7196 32289
rect 6564 32252 7196 32280
rect 5813 32215 5871 32221
rect 5813 32181 5825 32215
rect 5859 32212 5871 32215
rect 5994 32212 6000 32224
rect 5859 32184 6000 32212
rect 5859 32181 5871 32184
rect 5813 32175 5871 32181
rect 5994 32172 6000 32184
rect 6052 32172 6058 32224
rect 6564 32221 6592 32252
rect 7187 32243 7196 32252
rect 7248 32280 7254 32292
rect 8113 32283 8171 32289
rect 8113 32280 8125 32283
rect 7248 32252 8125 32280
rect 7190 32240 7196 32243
rect 7248 32240 7254 32252
rect 8113 32249 8125 32252
rect 8159 32280 8171 32283
rect 8935 32283 8993 32289
rect 8935 32280 8947 32283
rect 8159 32252 8947 32280
rect 8159 32249 8171 32252
rect 8113 32243 8171 32249
rect 8935 32249 8947 32252
rect 8981 32280 8993 32283
rect 9398 32280 9404 32292
rect 8981 32252 9404 32280
rect 8981 32249 8993 32252
rect 8935 32243 8993 32249
rect 9398 32240 9404 32252
rect 9456 32280 9462 32292
rect 9769 32283 9827 32289
rect 9769 32280 9781 32283
rect 9456 32252 9781 32280
rect 9456 32240 9462 32252
rect 9769 32249 9781 32252
rect 9815 32249 9827 32283
rect 10226 32280 10232 32292
rect 10139 32252 10232 32280
rect 9769 32243 9827 32249
rect 10226 32240 10232 32252
rect 10284 32280 10290 32292
rect 10796 32280 10824 32311
rect 10284 32252 10824 32280
rect 10284 32240 10290 32252
rect 12176 32224 12204 32320
rect 12472 32317 12484 32320
rect 12518 32317 12530 32351
rect 12472 32311 12530 32317
rect 6273 32215 6331 32221
rect 6273 32181 6285 32215
rect 6319 32212 6331 32215
rect 6549 32215 6607 32221
rect 6549 32212 6561 32215
rect 6319 32184 6561 32212
rect 6319 32181 6331 32184
rect 6273 32175 6331 32181
rect 6549 32181 6561 32184
rect 6595 32181 6607 32215
rect 10410 32212 10416 32224
rect 10371 32184 10416 32212
rect 6549 32175 6607 32181
rect 10410 32172 10416 32184
rect 10468 32212 10474 32224
rect 11333 32215 11391 32221
rect 11333 32212 11345 32215
rect 10468 32184 11345 32212
rect 10468 32172 10474 32184
rect 11333 32181 11345 32184
rect 11379 32181 11391 32215
rect 12158 32212 12164 32224
rect 12119 32184 12164 32212
rect 11333 32175 11391 32181
rect 12158 32172 12164 32184
rect 12216 32172 12222 32224
rect 13078 32212 13084 32224
rect 13039 32184 13084 32212
rect 13078 32172 13084 32184
rect 13136 32172 13142 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 9674 31968 9680 32020
rect 9732 32008 9738 32020
rect 9769 32011 9827 32017
rect 9769 32008 9781 32011
rect 9732 31980 9781 32008
rect 9732 31968 9738 31980
rect 9769 31977 9781 31980
rect 9815 31977 9827 32011
rect 9769 31971 9827 31977
rect 11379 32011 11437 32017
rect 11379 31977 11391 32011
rect 11425 32008 11437 32011
rect 11514 32008 11520 32020
rect 11425 31980 11520 32008
rect 11425 31977 11437 31980
rect 11379 31971 11437 31977
rect 11514 31968 11520 31980
rect 11572 32008 11578 32020
rect 11701 32011 11759 32017
rect 11701 32008 11713 32011
rect 11572 31980 11713 32008
rect 11572 31968 11578 31980
rect 11701 31977 11713 31980
rect 11747 31977 11759 32011
rect 11701 31971 11759 31977
rect 6822 31940 6828 31952
rect 6735 31912 6828 31940
rect 6822 31900 6828 31912
rect 6880 31940 6886 31952
rect 7469 31943 7527 31949
rect 7469 31940 7481 31943
rect 6880 31912 7481 31940
rect 6880 31900 6886 31912
rect 7469 31909 7481 31912
rect 7515 31909 7527 31943
rect 7469 31903 7527 31909
rect 8389 31943 8447 31949
rect 8389 31909 8401 31943
rect 8435 31940 8447 31943
rect 8754 31940 8760 31952
rect 8435 31912 8760 31940
rect 8435 31909 8447 31912
rect 8389 31903 8447 31909
rect 8754 31900 8760 31912
rect 8812 31900 8818 31952
rect 10686 31940 10692 31952
rect 10647 31912 10692 31940
rect 10686 31900 10692 31912
rect 10744 31900 10750 31952
rect 5810 31832 5816 31884
rect 5868 31872 5874 31884
rect 6089 31875 6147 31881
rect 6089 31872 6101 31875
rect 5868 31844 6101 31872
rect 5868 31832 5874 31844
rect 6089 31841 6101 31844
rect 6135 31841 6147 31875
rect 6638 31872 6644 31884
rect 6599 31844 6644 31872
rect 6089 31835 6147 31841
rect 6638 31832 6644 31844
rect 6696 31832 6702 31884
rect 7929 31875 7987 31881
rect 7929 31841 7941 31875
rect 7975 31841 7987 31875
rect 8110 31872 8116 31884
rect 8071 31844 8116 31872
rect 7929 31835 7987 31841
rect 7742 31764 7748 31816
rect 7800 31804 7806 31816
rect 7944 31804 7972 31835
rect 8110 31832 8116 31844
rect 8168 31832 8174 31884
rect 9953 31875 10011 31881
rect 9953 31841 9965 31875
rect 9999 31841 10011 31875
rect 10226 31872 10232 31884
rect 10187 31844 10232 31872
rect 9953 31835 10011 31841
rect 9968 31804 9996 31835
rect 10226 31832 10232 31844
rect 10284 31832 10290 31884
rect 11238 31832 11244 31884
rect 11296 31881 11302 31884
rect 11296 31875 11334 31881
rect 11322 31841 11334 31875
rect 11296 31835 11334 31841
rect 11296 31832 11302 31835
rect 10134 31804 10140 31816
rect 7800 31776 10140 31804
rect 7800 31764 7806 31776
rect 10134 31764 10140 31776
rect 10192 31764 10198 31816
rect 7193 31671 7251 31677
rect 7193 31637 7205 31671
rect 7239 31668 7251 31671
rect 7374 31668 7380 31680
rect 7239 31640 7380 31668
rect 7239 31637 7251 31640
rect 7193 31631 7251 31637
rect 7374 31628 7380 31640
rect 7432 31628 7438 31680
rect 8662 31668 8668 31680
rect 8623 31640 8668 31668
rect 8662 31628 8668 31640
rect 8720 31628 8726 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 5810 31464 5816 31476
rect 5771 31436 5816 31464
rect 5810 31424 5816 31436
rect 5868 31424 5874 31476
rect 9769 31467 9827 31473
rect 9769 31433 9781 31467
rect 9815 31464 9827 31467
rect 10226 31464 10232 31476
rect 9815 31436 10232 31464
rect 9815 31433 9827 31436
rect 9769 31427 9827 31433
rect 7374 31328 7380 31340
rect 7335 31300 7380 31328
rect 7374 31288 7380 31300
rect 7432 31288 7438 31340
rect 9306 31328 9312 31340
rect 9267 31300 9312 31328
rect 9306 31288 9312 31300
rect 9364 31288 9370 31340
rect 6914 31260 6920 31272
rect 6875 31232 6920 31260
rect 6914 31220 6920 31232
rect 6972 31220 6978 31272
rect 7285 31263 7343 31269
rect 7285 31229 7297 31263
rect 7331 31229 7343 31263
rect 7285 31223 7343 31229
rect 6181 31127 6239 31133
rect 6181 31093 6193 31127
rect 6227 31124 6239 31127
rect 6638 31124 6644 31136
rect 6227 31096 6644 31124
rect 6227 31093 6239 31096
rect 6181 31087 6239 31093
rect 6638 31084 6644 31096
rect 6696 31124 6702 31136
rect 7300 31124 7328 31223
rect 8294 31220 8300 31272
rect 8352 31260 8358 31272
rect 8662 31260 8668 31272
rect 8352 31232 8668 31260
rect 8352 31220 8358 31232
rect 8662 31220 8668 31232
rect 8720 31220 8726 31272
rect 9217 31263 9275 31269
rect 9217 31229 9229 31263
rect 9263 31260 9275 31263
rect 9784 31260 9812 31427
rect 10226 31424 10232 31436
rect 10284 31424 10290 31476
rect 10689 31331 10747 31337
rect 10689 31297 10701 31331
rect 10735 31328 10747 31331
rect 10778 31328 10784 31340
rect 10735 31300 10784 31328
rect 10735 31297 10747 31300
rect 10689 31291 10747 31297
rect 10778 31288 10784 31300
rect 10836 31288 10842 31340
rect 10134 31260 10140 31272
rect 9263 31232 9812 31260
rect 10095 31232 10140 31260
rect 9263 31229 9275 31232
rect 9217 31223 9275 31229
rect 8573 31195 8631 31201
rect 8573 31161 8585 31195
rect 8619 31192 8631 31195
rect 9232 31192 9260 31223
rect 10134 31220 10140 31232
rect 10192 31220 10198 31272
rect 8619 31164 9260 31192
rect 10505 31195 10563 31201
rect 8619 31161 8631 31164
rect 8573 31155 8631 31161
rect 8680 31136 8708 31164
rect 10505 31161 10517 31195
rect 10551 31192 10563 31195
rect 10781 31195 10839 31201
rect 10781 31192 10793 31195
rect 10551 31164 10793 31192
rect 10551 31161 10563 31164
rect 10505 31155 10563 31161
rect 10781 31161 10793 31164
rect 10827 31192 10839 31195
rect 10962 31192 10968 31204
rect 10827 31164 10968 31192
rect 10827 31161 10839 31164
rect 10781 31155 10839 31161
rect 10962 31152 10968 31164
rect 11020 31152 11026 31204
rect 11333 31195 11391 31201
rect 11333 31161 11345 31195
rect 11379 31192 11391 31195
rect 12158 31192 12164 31204
rect 11379 31164 12164 31192
rect 11379 31161 11391 31164
rect 11333 31155 11391 31161
rect 12158 31152 12164 31164
rect 12216 31152 12222 31204
rect 7837 31127 7895 31133
rect 7837 31124 7849 31127
rect 6696 31096 7849 31124
rect 6696 31084 6702 31096
rect 7837 31093 7849 31096
rect 7883 31124 7895 31127
rect 8110 31124 8116 31136
rect 7883 31096 8116 31124
rect 7883 31093 7895 31096
rect 7837 31087 7895 31093
rect 8110 31084 8116 31096
rect 8168 31084 8174 31136
rect 8662 31084 8668 31136
rect 8720 31084 8726 31136
rect 11238 31084 11244 31136
rect 11296 31124 11302 31136
rect 11514 31124 11520 31136
rect 11296 31096 11520 31124
rect 11296 31084 11302 31096
rect 11514 31084 11520 31096
rect 11572 31124 11578 31136
rect 11609 31127 11667 31133
rect 11609 31124 11621 31127
rect 11572 31096 11621 31124
rect 11572 31084 11578 31096
rect 11609 31093 11621 31096
rect 11655 31093 11667 31127
rect 11609 31087 11667 31093
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 7742 30920 7748 30932
rect 7703 30892 7748 30920
rect 7742 30880 7748 30892
rect 7800 30880 7806 30932
rect 9490 30920 9496 30932
rect 9451 30892 9496 30920
rect 9490 30880 9496 30892
rect 9548 30920 9554 30932
rect 10778 30920 10784 30932
rect 9548 30892 9812 30920
rect 10739 30892 10784 30920
rect 9548 30880 9554 30892
rect 8202 30852 8208 30864
rect 8163 30824 8208 30852
rect 8202 30812 8208 30824
rect 8260 30812 8266 30864
rect 9784 30861 9812 30892
rect 10778 30880 10784 30892
rect 10836 30880 10842 30932
rect 9769 30855 9827 30861
rect 9769 30821 9781 30855
rect 9815 30821 9827 30855
rect 9769 30815 9827 30821
rect 9858 30812 9864 30864
rect 9916 30852 9922 30864
rect 11422 30852 11428 30864
rect 9916 30824 9961 30852
rect 11383 30824 11428 30852
rect 9916 30812 9922 30824
rect 11422 30812 11428 30824
rect 11480 30812 11486 30864
rect 7006 30716 7012 30728
rect 6967 30688 7012 30716
rect 7006 30676 7012 30688
rect 7064 30676 7070 30728
rect 7926 30676 7932 30728
rect 7984 30716 7990 30728
rect 8113 30719 8171 30725
rect 8113 30716 8125 30719
rect 7984 30688 8125 30716
rect 7984 30676 7990 30688
rect 8113 30685 8125 30688
rect 8159 30685 8171 30719
rect 8386 30716 8392 30728
rect 8347 30688 8392 30716
rect 8113 30679 8171 30685
rect 8386 30676 8392 30688
rect 8444 30716 8450 30728
rect 10045 30719 10103 30725
rect 10045 30716 10057 30719
rect 8444 30688 10057 30716
rect 8444 30676 8450 30688
rect 10045 30685 10057 30688
rect 10091 30685 10103 30719
rect 11330 30716 11336 30728
rect 11291 30688 11336 30716
rect 10045 30679 10103 30685
rect 11330 30676 11336 30688
rect 11388 30676 11394 30728
rect 11977 30719 12035 30725
rect 11977 30685 11989 30719
rect 12023 30716 12035 30719
rect 12158 30716 12164 30728
rect 12023 30688 12164 30716
rect 12023 30685 12035 30688
rect 11977 30679 12035 30685
rect 12158 30676 12164 30688
rect 12216 30676 12222 30728
rect 6914 30580 6920 30592
rect 6827 30552 6920 30580
rect 6914 30540 6920 30552
rect 6972 30580 6978 30592
rect 8386 30580 8392 30592
rect 6972 30552 8392 30580
rect 6972 30540 6978 30552
rect 8386 30540 8392 30552
rect 8444 30540 8450 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 11333 30379 11391 30385
rect 11333 30345 11345 30379
rect 11379 30376 11391 30379
rect 11422 30376 11428 30388
rect 11379 30348 11428 30376
rect 11379 30345 11391 30348
rect 11333 30339 11391 30345
rect 8478 30268 8484 30320
rect 8536 30308 8542 30320
rect 8987 30311 9045 30317
rect 8987 30308 8999 30311
rect 8536 30280 8999 30308
rect 8536 30268 8542 30280
rect 8987 30277 8999 30280
rect 9033 30277 9045 30311
rect 8987 30271 9045 30277
rect 10781 30311 10839 30317
rect 10781 30277 10793 30311
rect 10827 30308 10839 30311
rect 11348 30308 11376 30339
rect 11422 30336 11428 30348
rect 11480 30336 11486 30388
rect 10827 30280 11376 30308
rect 10827 30277 10839 30280
rect 10781 30271 10839 30277
rect 11330 30200 11336 30252
rect 11388 30240 11394 30252
rect 11609 30243 11667 30249
rect 11609 30240 11621 30243
rect 11388 30212 11621 30240
rect 11388 30200 11394 30212
rect 11609 30209 11621 30212
rect 11655 30209 11667 30243
rect 11609 30203 11667 30209
rect 7466 30172 7472 30184
rect 7427 30144 7472 30172
rect 7466 30132 7472 30144
rect 7524 30132 7530 30184
rect 7745 30175 7803 30181
rect 7745 30141 7757 30175
rect 7791 30141 7803 30175
rect 8754 30172 8760 30184
rect 8715 30144 8760 30172
rect 7745 30135 7803 30141
rect 7760 30104 7788 30135
rect 8754 30132 8760 30144
rect 8812 30172 8818 30184
rect 8884 30175 8942 30181
rect 8884 30172 8896 30175
rect 8812 30144 8896 30172
rect 8812 30132 8818 30144
rect 8884 30141 8896 30144
rect 8930 30141 8942 30175
rect 8884 30135 8942 30141
rect 9861 30175 9919 30181
rect 9861 30141 9873 30175
rect 9907 30172 9919 30175
rect 9950 30172 9956 30184
rect 9907 30144 9956 30172
rect 9907 30141 9919 30144
rect 9861 30135 9919 30141
rect 9950 30132 9956 30144
rect 10008 30132 10014 30184
rect 9766 30104 9772 30116
rect 7116 30076 7788 30104
rect 9324 30076 9772 30104
rect 6638 29996 6644 30048
rect 6696 30036 6702 30048
rect 7116 30045 7144 30076
rect 9324 30048 9352 30076
rect 9766 30064 9772 30076
rect 9824 30064 9830 30116
rect 10223 30107 10281 30113
rect 10223 30104 10235 30107
rect 9876 30076 10235 30104
rect 7101 30039 7159 30045
rect 7101 30036 7113 30039
rect 6696 30008 7113 30036
rect 6696 29996 6702 30008
rect 7101 30005 7113 30008
rect 7147 30005 7159 30039
rect 7558 30036 7564 30048
rect 7519 30008 7564 30036
rect 7101 29999 7159 30005
rect 7558 29996 7564 30008
rect 7616 29996 7622 30048
rect 8294 30036 8300 30048
rect 8255 30008 8300 30036
rect 8294 29996 8300 30008
rect 8352 29996 8358 30048
rect 9306 30036 9312 30048
rect 9267 30008 9312 30036
rect 9306 29996 9312 30008
rect 9364 29996 9370 30048
rect 9398 29996 9404 30048
rect 9456 30036 9462 30048
rect 9677 30039 9735 30045
rect 9677 30036 9689 30039
rect 9456 30008 9689 30036
rect 9456 29996 9462 30008
rect 9677 30005 9689 30008
rect 9723 30036 9735 30039
rect 9876 30036 9904 30076
rect 10223 30073 10235 30076
rect 10269 30104 10281 30107
rect 10410 30104 10416 30116
rect 10269 30076 10416 30104
rect 10269 30073 10281 30076
rect 10223 30067 10281 30073
rect 10410 30064 10416 30076
rect 10468 30104 10474 30116
rect 11054 30104 11060 30116
rect 10468 30076 11060 30104
rect 10468 30064 10474 30076
rect 11054 30064 11060 30076
rect 11112 30064 11118 30116
rect 9723 30008 9904 30036
rect 9723 30005 9735 30008
rect 9677 29999 9735 30005
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 7466 29832 7472 29844
rect 7427 29804 7472 29832
rect 7466 29792 7472 29804
rect 7524 29792 7530 29844
rect 7926 29832 7932 29844
rect 7887 29804 7932 29832
rect 7926 29792 7932 29804
rect 7984 29792 7990 29844
rect 10962 29832 10968 29844
rect 10923 29804 10968 29832
rect 10962 29792 10968 29804
rect 11020 29792 11026 29844
rect 7484 29764 7512 29792
rect 8386 29764 8392 29776
rect 7484 29736 8392 29764
rect 8386 29724 8392 29736
rect 8444 29724 8450 29776
rect 10410 29773 10416 29776
rect 10407 29764 10416 29773
rect 10371 29736 10416 29764
rect 10407 29727 10416 29736
rect 10410 29724 10416 29727
rect 10468 29724 10474 29776
rect 11974 29764 11980 29776
rect 11935 29736 11980 29764
rect 11974 29724 11980 29736
rect 12032 29724 12038 29776
rect 6549 29699 6607 29705
rect 6549 29665 6561 29699
rect 6595 29665 6607 29699
rect 6549 29659 6607 29665
rect 6564 29628 6592 29659
rect 6638 29656 6644 29708
rect 6696 29696 6702 29708
rect 6917 29699 6975 29705
rect 6917 29696 6929 29699
rect 6696 29668 6929 29696
rect 6696 29656 6702 29668
rect 6917 29665 6929 29668
rect 6963 29665 6975 29699
rect 8202 29696 8208 29708
rect 8163 29668 8208 29696
rect 6917 29659 6975 29665
rect 8202 29656 8208 29668
rect 8260 29656 8266 29708
rect 8573 29699 8631 29705
rect 8573 29665 8585 29699
rect 8619 29696 8631 29699
rect 8662 29696 8668 29708
rect 8619 29668 8668 29696
rect 8619 29665 8631 29668
rect 8573 29659 8631 29665
rect 8662 29656 8668 29668
rect 8720 29656 8726 29708
rect 6730 29628 6736 29640
rect 6564 29600 6736 29628
rect 6730 29588 6736 29600
rect 6788 29588 6794 29640
rect 7190 29628 7196 29640
rect 7151 29600 7196 29628
rect 7190 29588 7196 29600
rect 7248 29588 7254 29640
rect 8757 29631 8815 29637
rect 8757 29597 8769 29631
rect 8803 29628 8815 29631
rect 8846 29628 8852 29640
rect 8803 29600 8852 29628
rect 8803 29597 8815 29600
rect 8757 29591 8815 29597
rect 8846 29588 8852 29600
rect 8904 29628 8910 29640
rect 9125 29631 9183 29637
rect 9125 29628 9137 29631
rect 8904 29600 9137 29628
rect 8904 29588 8910 29600
rect 9125 29597 9137 29600
rect 9171 29597 9183 29631
rect 9125 29591 9183 29597
rect 10045 29631 10103 29637
rect 10045 29597 10057 29631
rect 10091 29628 10103 29631
rect 10686 29628 10692 29640
rect 10091 29600 10692 29628
rect 10091 29597 10103 29600
rect 10045 29591 10103 29597
rect 10686 29588 10692 29600
rect 10744 29588 10750 29640
rect 11882 29628 11888 29640
rect 11843 29600 11888 29628
rect 11882 29588 11888 29600
rect 11940 29588 11946 29640
rect 12158 29628 12164 29640
rect 12119 29600 12164 29628
rect 12158 29588 12164 29600
rect 12216 29588 12222 29640
rect 5261 29495 5319 29501
rect 5261 29461 5273 29495
rect 5307 29492 5319 29495
rect 5350 29492 5356 29504
rect 5307 29464 5356 29492
rect 5307 29461 5319 29464
rect 5261 29455 5319 29461
rect 5350 29452 5356 29464
rect 5408 29452 5414 29504
rect 9950 29492 9956 29504
rect 9911 29464 9956 29492
rect 9950 29452 9956 29464
rect 10008 29452 10014 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 8294 29288 8300 29300
rect 8255 29260 8300 29288
rect 8294 29248 8300 29260
rect 8352 29248 8358 29300
rect 8662 29288 8668 29300
rect 8623 29260 8668 29288
rect 8662 29248 8668 29260
rect 8720 29248 8726 29300
rect 9033 29291 9091 29297
rect 9033 29257 9045 29291
rect 9079 29288 9091 29291
rect 10410 29288 10416 29300
rect 9079 29260 10416 29288
rect 9079 29257 9091 29260
rect 9033 29251 9091 29257
rect 8570 29180 8576 29232
rect 8628 29180 8634 29232
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29152 5135 29155
rect 5258 29152 5264 29164
rect 5123 29124 5264 29152
rect 5123 29121 5135 29124
rect 5077 29115 5135 29121
rect 5258 29112 5264 29124
rect 5316 29112 5322 29164
rect 5902 29152 5908 29164
rect 5863 29124 5908 29152
rect 5902 29112 5908 29124
rect 5960 29112 5966 29164
rect 7190 29112 7196 29164
rect 7248 29152 7254 29164
rect 7377 29155 7435 29161
rect 7377 29152 7389 29155
rect 7248 29124 7389 29152
rect 7248 29112 7254 29124
rect 7377 29121 7389 29124
rect 7423 29121 7435 29155
rect 7377 29115 7435 29121
rect 8588 29096 8616 29180
rect 8846 29112 8852 29164
rect 8904 29152 8910 29164
rect 9125 29155 9183 29161
rect 9125 29152 9137 29155
rect 8904 29124 9137 29152
rect 8904 29112 8910 29124
rect 9125 29121 9137 29124
rect 9171 29121 9183 29155
rect 9125 29115 9183 29121
rect 6549 29087 6607 29093
rect 6549 29053 6561 29087
rect 6595 29084 6607 29087
rect 6638 29084 6644 29096
rect 6595 29056 6644 29084
rect 6595 29053 6607 29056
rect 6549 29047 6607 29053
rect 6638 29044 6644 29056
rect 6696 29084 6702 29096
rect 7926 29084 7932 29096
rect 6696 29056 7932 29084
rect 6696 29044 6702 29056
rect 7926 29044 7932 29056
rect 7984 29044 7990 29096
rect 8570 29044 8576 29096
rect 8628 29044 8634 29096
rect 4890 28976 4896 29028
rect 4948 29016 4954 29028
rect 4982 29016 4988 29028
rect 4948 28988 4988 29016
rect 4948 28976 4954 28988
rect 4982 28976 4988 28988
rect 5040 28976 5046 29028
rect 5350 29016 5356 29028
rect 5311 28988 5356 29016
rect 5350 28976 5356 28988
rect 5408 28976 5414 29028
rect 7285 29019 7343 29025
rect 7285 28985 7297 29019
rect 7331 29016 7343 29019
rect 7739 29019 7797 29025
rect 7739 29016 7751 29019
rect 7331 28988 7751 29016
rect 7331 28985 7343 28988
rect 7285 28979 7343 28985
rect 7739 28985 7751 28988
rect 7785 29016 7797 29019
rect 8110 29016 8116 29028
rect 7785 28988 8116 29016
rect 7785 28985 7797 28988
rect 7739 28979 7797 28985
rect 8110 28976 8116 28988
rect 8168 29016 8174 29028
rect 9508 29025 9536 29260
rect 10410 29248 10416 29260
rect 10468 29248 10474 29300
rect 11882 29288 11888 29300
rect 11843 29260 11888 29288
rect 11882 29248 11888 29260
rect 11940 29248 11946 29300
rect 10873 29155 10931 29161
rect 10873 29121 10885 29155
rect 10919 29152 10931 29155
rect 11900 29152 11928 29248
rect 10919 29124 11928 29152
rect 10919 29121 10931 29124
rect 10873 29115 10931 29121
rect 10045 29087 10103 29093
rect 10045 29053 10057 29087
rect 10091 29084 10103 29087
rect 11974 29084 11980 29096
rect 10091 29056 11980 29084
rect 10091 29053 10103 29056
rect 10045 29047 10103 29053
rect 11974 29044 11980 29056
rect 12032 29084 12038 29096
rect 12161 29087 12219 29093
rect 12161 29084 12173 29087
rect 12032 29056 12173 29084
rect 12032 29044 12038 29056
rect 12161 29053 12173 29056
rect 12207 29053 12219 29087
rect 12161 29047 12219 29053
rect 9487 29019 9545 29025
rect 9487 29016 9499 29019
rect 8168 28988 9499 29016
rect 8168 28976 8174 28988
rect 9487 28985 9499 28988
rect 9533 28985 9545 29019
rect 9487 28979 9545 28985
rect 9674 28976 9680 29028
rect 9732 29016 9738 29028
rect 10318 29016 10324 29028
rect 9732 28988 10324 29016
rect 9732 28976 9738 28988
rect 10318 28976 10324 28988
rect 10376 28976 10382 29028
rect 10686 28948 10692 28960
rect 10647 28920 10692 28948
rect 10686 28908 10692 28920
rect 10744 28908 10750 28960
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 7190 28704 7196 28756
rect 7248 28744 7254 28756
rect 7469 28747 7527 28753
rect 7469 28744 7481 28747
rect 7248 28716 7481 28744
rect 7248 28704 7254 28716
rect 7469 28713 7481 28716
rect 7515 28713 7527 28747
rect 7469 28707 7527 28713
rect 8573 28747 8631 28753
rect 8573 28713 8585 28747
rect 8619 28744 8631 28747
rect 9306 28744 9312 28756
rect 8619 28716 9312 28744
rect 8619 28713 8631 28716
rect 8573 28707 8631 28713
rect 9306 28704 9312 28716
rect 9364 28704 9370 28756
rect 9950 28744 9956 28756
rect 9911 28716 9956 28744
rect 9950 28704 9956 28716
rect 10008 28704 10014 28756
rect 11425 28747 11483 28753
rect 11425 28713 11437 28747
rect 11471 28713 11483 28747
rect 11425 28707 11483 28713
rect 8015 28679 8073 28685
rect 8015 28645 8027 28679
rect 8061 28676 8073 28679
rect 8110 28676 8116 28688
rect 8061 28648 8116 28676
rect 8061 28645 8073 28648
rect 8015 28639 8073 28645
rect 8110 28636 8116 28648
rect 8168 28636 8174 28688
rect 8662 28636 8668 28688
rect 8720 28676 8726 28688
rect 11440 28676 11468 28707
rect 8720 28648 11468 28676
rect 8720 28636 8726 28648
rect 4890 28617 4896 28620
rect 4868 28611 4896 28617
rect 4868 28577 4880 28611
rect 4868 28571 4896 28577
rect 4890 28568 4896 28571
rect 4948 28568 4954 28620
rect 6362 28608 6368 28620
rect 6323 28580 6368 28608
rect 6362 28568 6368 28580
rect 6420 28568 6426 28620
rect 6638 28608 6644 28620
rect 6599 28580 6644 28608
rect 6638 28568 6644 28580
rect 6696 28568 6702 28620
rect 7558 28568 7564 28620
rect 7616 28608 7622 28620
rect 7653 28611 7711 28617
rect 7653 28608 7665 28611
rect 7616 28580 7665 28608
rect 7616 28568 7622 28580
rect 7653 28577 7665 28580
rect 7699 28577 7711 28611
rect 7653 28571 7711 28577
rect 8294 28568 8300 28620
rect 8352 28608 8358 28620
rect 10152 28617 10180 28648
rect 8849 28611 8907 28617
rect 8849 28608 8861 28611
rect 8352 28580 8861 28608
rect 8352 28568 8358 28580
rect 8849 28577 8861 28580
rect 8895 28577 8907 28611
rect 8849 28571 8907 28577
rect 9677 28611 9735 28617
rect 9677 28577 9689 28611
rect 9723 28577 9735 28611
rect 9677 28571 9735 28577
rect 10137 28611 10195 28617
rect 10137 28577 10149 28611
rect 10183 28577 10195 28611
rect 11238 28608 11244 28620
rect 11199 28580 11244 28608
rect 10137 28571 10195 28577
rect 6822 28540 6828 28552
rect 6783 28512 6828 28540
rect 6822 28500 6828 28512
rect 6880 28500 6886 28552
rect 8386 28500 8392 28552
rect 8444 28540 8450 28552
rect 9692 28540 9720 28571
rect 11238 28568 11244 28580
rect 11296 28568 11302 28620
rect 10410 28540 10416 28552
rect 8444 28512 10416 28540
rect 8444 28500 8450 28512
rect 10410 28500 10416 28512
rect 10468 28500 10474 28552
rect 4798 28364 4804 28416
rect 4856 28404 4862 28416
rect 4939 28407 4997 28413
rect 4939 28404 4951 28407
rect 4856 28376 4951 28404
rect 4856 28364 4862 28376
rect 4939 28373 4951 28376
rect 4985 28373 4997 28407
rect 5258 28404 5264 28416
rect 5219 28376 5264 28404
rect 4939 28367 4997 28373
rect 5258 28364 5264 28376
rect 5316 28364 5322 28416
rect 5350 28364 5356 28416
rect 5408 28404 5414 28416
rect 5629 28407 5687 28413
rect 5629 28404 5641 28407
rect 5408 28376 5641 28404
rect 5408 28364 5414 28376
rect 5629 28373 5641 28376
rect 5675 28373 5687 28407
rect 5629 28367 5687 28373
rect 6730 28364 6736 28416
rect 6788 28404 6794 28416
rect 7193 28407 7251 28413
rect 7193 28404 7205 28407
rect 6788 28376 7205 28404
rect 6788 28364 6794 28376
rect 7193 28373 7205 28376
rect 7239 28404 7251 28407
rect 9398 28404 9404 28416
rect 7239 28376 9404 28404
rect 7239 28373 7251 28376
rect 7193 28367 7251 28373
rect 9398 28364 9404 28376
rect 9456 28364 9462 28416
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 6181 28203 6239 28209
rect 6181 28169 6193 28203
rect 6227 28200 6239 28203
rect 6638 28200 6644 28212
rect 6227 28172 6644 28200
rect 6227 28169 6239 28172
rect 6181 28163 6239 28169
rect 6638 28160 6644 28172
rect 6696 28160 6702 28212
rect 7558 28160 7564 28212
rect 7616 28200 7622 28212
rect 8389 28203 8447 28209
rect 8389 28200 8401 28203
rect 7616 28172 8401 28200
rect 7616 28160 7622 28172
rect 8389 28169 8401 28172
rect 8435 28169 8447 28203
rect 8389 28163 8447 28169
rect 8662 28160 8668 28212
rect 8720 28200 8726 28212
rect 9125 28203 9183 28209
rect 9125 28200 9137 28203
rect 8720 28172 9137 28200
rect 8720 28160 8726 28172
rect 9125 28169 9137 28172
rect 9171 28200 9183 28203
rect 10321 28203 10379 28209
rect 10321 28200 10333 28203
rect 9171 28172 10333 28200
rect 9171 28169 9183 28172
rect 9125 28163 9183 28169
rect 5626 28132 5632 28144
rect 4448 28104 5632 28132
rect 3234 27956 3240 28008
rect 3292 27996 3298 28008
rect 4448 28005 4476 28104
rect 5626 28092 5632 28104
rect 5684 28092 5690 28144
rect 7742 28132 7748 28144
rect 7703 28104 7748 28132
rect 7742 28092 7748 28104
rect 7800 28092 7806 28144
rect 8110 28132 8116 28144
rect 8071 28104 8116 28132
rect 8110 28092 8116 28104
rect 8168 28092 8174 28144
rect 5077 28067 5135 28073
rect 5077 28033 5089 28067
rect 5123 28064 5135 28067
rect 5350 28064 5356 28076
rect 5123 28036 5356 28064
rect 5123 28033 5135 28036
rect 5077 28027 5135 28033
rect 5350 28024 5356 28036
rect 5408 28024 5414 28076
rect 6822 28064 6828 28076
rect 6783 28036 6828 28064
rect 6822 28024 6828 28036
rect 6880 28024 6886 28076
rect 8386 28024 8392 28076
rect 8444 28064 8450 28076
rect 8757 28067 8815 28073
rect 8757 28064 8769 28067
rect 8444 28036 8769 28064
rect 8444 28024 8450 28036
rect 8757 28033 8769 28036
rect 8803 28033 8815 28067
rect 8757 28027 8815 28033
rect 4008 27999 4066 28005
rect 4008 27996 4020 27999
rect 3292 27968 4020 27996
rect 3292 27956 3298 27968
rect 4008 27965 4020 27968
rect 4054 27996 4066 27999
rect 4433 27999 4491 28005
rect 4433 27996 4445 27999
rect 4054 27968 4445 27996
rect 4054 27965 4066 27968
rect 4008 27959 4066 27965
rect 4433 27965 4445 27968
rect 4479 27965 4491 27999
rect 9398 27996 9404 28008
rect 9359 27968 9404 27996
rect 4433 27959 4491 27965
rect 9398 27956 9404 27968
rect 9456 27956 9462 28008
rect 9784 28005 9812 28172
rect 10321 28169 10333 28172
rect 10367 28169 10379 28203
rect 11054 28200 11060 28212
rect 11015 28172 11060 28200
rect 10321 28163 10379 28169
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 10045 28067 10103 28073
rect 10045 28033 10057 28067
rect 10091 28064 10103 28067
rect 10686 28064 10692 28076
rect 10091 28036 10692 28064
rect 10091 28033 10103 28036
rect 10045 28027 10103 28033
rect 10686 28024 10692 28036
rect 10744 28024 10750 28076
rect 9769 27999 9827 28005
rect 9769 27965 9781 27999
rect 9815 27965 9827 27999
rect 9769 27959 9827 27965
rect 10134 27956 10140 28008
rect 10192 27996 10198 28008
rect 10873 27999 10931 28005
rect 10873 27996 10885 27999
rect 10192 27968 10885 27996
rect 10192 27956 10198 27968
rect 10873 27965 10885 27968
rect 10919 27996 10931 27999
rect 11701 27999 11759 28005
rect 11701 27996 11713 27999
rect 10919 27968 11713 27996
rect 10919 27965 10931 27968
rect 10873 27959 10931 27965
rect 11701 27965 11713 27968
rect 11747 27965 11759 27999
rect 11701 27959 11759 27965
rect 5169 27931 5227 27937
rect 5169 27897 5181 27931
rect 5215 27928 5227 27931
rect 5258 27928 5264 27940
rect 5215 27900 5264 27928
rect 5215 27897 5227 27900
rect 5169 27891 5227 27897
rect 5258 27888 5264 27900
rect 5316 27888 5322 27940
rect 5718 27928 5724 27940
rect 5679 27900 5724 27928
rect 5718 27888 5724 27900
rect 5776 27888 5782 27940
rect 6641 27931 6699 27937
rect 6641 27897 6653 27931
rect 6687 27928 6699 27931
rect 7187 27931 7245 27937
rect 7187 27928 7199 27931
rect 6687 27900 7199 27928
rect 6687 27897 6699 27900
rect 6641 27891 6699 27897
rect 7187 27897 7199 27900
rect 7233 27928 7245 27931
rect 7926 27928 7932 27940
rect 7233 27900 7932 27928
rect 7233 27897 7245 27900
rect 7187 27891 7245 27897
rect 7926 27888 7932 27900
rect 7984 27928 7990 27940
rect 8110 27928 8116 27940
rect 7984 27900 8116 27928
rect 7984 27888 7990 27900
rect 8110 27888 8116 27900
rect 8168 27888 8174 27940
rect 4062 27820 4068 27872
rect 4120 27869 4126 27872
rect 4120 27863 4169 27869
rect 4120 27829 4123 27863
rect 4157 27829 4169 27863
rect 4890 27860 4896 27872
rect 4851 27832 4896 27860
rect 4120 27823 4169 27829
rect 4120 27820 4126 27823
rect 4890 27820 4896 27832
rect 4948 27820 4954 27872
rect 10318 27820 10324 27872
rect 10376 27860 10382 27872
rect 11238 27860 11244 27872
rect 10376 27832 11244 27860
rect 10376 27820 10382 27832
rect 11238 27820 11244 27832
rect 11296 27860 11302 27872
rect 11333 27863 11391 27869
rect 11333 27860 11345 27863
rect 11296 27832 11345 27860
rect 11296 27820 11302 27832
rect 11333 27829 11345 27832
rect 11379 27829 11391 27863
rect 11333 27823 11391 27829
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 4798 27656 4804 27668
rect 4759 27628 4804 27656
rect 4798 27616 4804 27628
rect 4856 27616 4862 27668
rect 5169 27659 5227 27665
rect 5169 27625 5181 27659
rect 5215 27656 5227 27659
rect 5258 27656 5264 27668
rect 5215 27628 5264 27656
rect 5215 27625 5227 27628
rect 5169 27619 5227 27625
rect 5258 27616 5264 27628
rect 5316 27616 5322 27668
rect 6178 27616 6184 27668
rect 6236 27656 6242 27668
rect 6365 27659 6423 27665
rect 6365 27656 6377 27659
rect 6236 27628 6377 27656
rect 6236 27616 6242 27628
rect 6365 27625 6377 27628
rect 6411 27625 6423 27659
rect 6365 27619 6423 27625
rect 6733 27659 6791 27665
rect 6733 27625 6745 27659
rect 6779 27656 6791 27659
rect 6822 27656 6828 27668
rect 6779 27628 6828 27656
rect 6779 27625 6791 27628
rect 6733 27619 6791 27625
rect 6822 27616 6828 27628
rect 6880 27616 6886 27668
rect 4387 27591 4445 27597
rect 4387 27557 4399 27591
rect 4433 27588 4445 27591
rect 5350 27588 5356 27600
rect 4433 27560 5356 27588
rect 4433 27557 4445 27560
rect 4387 27551 4445 27557
rect 5350 27548 5356 27560
rect 5408 27548 5414 27600
rect 5445 27591 5503 27597
rect 5445 27557 5457 27591
rect 5491 27588 5503 27591
rect 5626 27588 5632 27600
rect 5491 27560 5632 27588
rect 5491 27557 5503 27560
rect 5445 27551 5503 27557
rect 5626 27548 5632 27560
rect 5684 27588 5690 27600
rect 6270 27588 6276 27600
rect 5684 27560 6276 27588
rect 5684 27548 5690 27560
rect 6270 27548 6276 27560
rect 6328 27588 6334 27600
rect 7009 27591 7067 27597
rect 7009 27588 7021 27591
rect 6328 27560 7021 27588
rect 6328 27548 6334 27560
rect 7009 27557 7021 27560
rect 7055 27557 7067 27591
rect 7009 27551 7067 27557
rect 7098 27548 7104 27600
rect 7156 27588 7162 27600
rect 7374 27588 7380 27600
rect 7156 27560 7380 27588
rect 7156 27548 7162 27560
rect 7374 27548 7380 27560
rect 7432 27548 7438 27600
rect 9858 27588 9864 27600
rect 9819 27560 9864 27588
rect 9858 27548 9864 27560
rect 9916 27548 9922 27600
rect 11425 27591 11483 27597
rect 11425 27557 11437 27591
rect 11471 27588 11483 27591
rect 11974 27588 11980 27600
rect 11471 27560 11980 27588
rect 11471 27557 11483 27560
rect 11425 27551 11483 27557
rect 11974 27548 11980 27560
rect 12032 27548 12038 27600
rect 4300 27523 4358 27529
rect 4300 27489 4312 27523
rect 4346 27520 4358 27523
rect 4522 27520 4528 27532
rect 4346 27492 4528 27520
rect 4346 27489 4358 27492
rect 4300 27483 4358 27489
rect 4522 27480 4528 27492
rect 4580 27480 4586 27532
rect 8386 27480 8392 27532
rect 8444 27529 8450 27532
rect 8444 27523 8482 27529
rect 8470 27489 8482 27523
rect 8444 27483 8482 27489
rect 8444 27480 8450 27483
rect 12802 27480 12808 27532
rect 12860 27529 12866 27532
rect 12860 27523 12898 27529
rect 12886 27489 12898 27523
rect 12860 27483 12898 27489
rect 12860 27480 12866 27483
rect 5350 27452 5356 27464
rect 5311 27424 5356 27452
rect 5350 27412 5356 27424
rect 5408 27412 5414 27464
rect 5718 27452 5724 27464
rect 5679 27424 5724 27452
rect 5718 27412 5724 27424
rect 5776 27412 5782 27464
rect 6917 27455 6975 27461
rect 6917 27421 6929 27455
rect 6963 27452 6975 27455
rect 7834 27452 7840 27464
rect 6963 27424 7840 27452
rect 6963 27421 6975 27424
rect 6917 27415 6975 27421
rect 7834 27412 7840 27424
rect 7892 27412 7898 27464
rect 9766 27452 9772 27464
rect 9727 27424 9772 27452
rect 9766 27412 9772 27424
rect 9824 27412 9830 27464
rect 10226 27412 10232 27464
rect 10284 27452 10290 27464
rect 10413 27455 10471 27461
rect 10413 27452 10425 27455
rect 10284 27424 10425 27452
rect 10284 27412 10290 27424
rect 10413 27421 10425 27424
rect 10459 27452 10471 27455
rect 11333 27455 11391 27461
rect 11333 27452 11345 27455
rect 10459 27424 11345 27452
rect 10459 27421 10471 27424
rect 10413 27415 10471 27421
rect 11333 27421 11345 27424
rect 11379 27452 11391 27455
rect 11514 27452 11520 27464
rect 11379 27424 11520 27452
rect 11379 27421 11391 27424
rect 11333 27415 11391 27421
rect 11514 27412 11520 27424
rect 11572 27412 11578 27464
rect 11977 27455 12035 27461
rect 11977 27421 11989 27455
rect 12023 27452 12035 27455
rect 12066 27452 12072 27464
rect 12023 27424 12072 27452
rect 12023 27421 12035 27424
rect 11977 27415 12035 27421
rect 12066 27412 12072 27424
rect 12124 27412 12130 27464
rect 7006 27344 7012 27396
rect 7064 27384 7070 27396
rect 7469 27387 7527 27393
rect 7469 27384 7481 27387
rect 7064 27356 7481 27384
rect 7064 27344 7070 27356
rect 7469 27353 7481 27356
rect 7515 27353 7527 27387
rect 7469 27347 7527 27353
rect 5994 27276 6000 27328
rect 6052 27316 6058 27328
rect 6638 27316 6644 27328
rect 6052 27288 6644 27316
rect 6052 27276 6058 27288
rect 6638 27276 6644 27288
rect 6696 27276 6702 27328
rect 8527 27319 8585 27325
rect 8527 27285 8539 27319
rect 8573 27316 8585 27319
rect 8846 27316 8852 27328
rect 8573 27288 8852 27316
rect 8573 27285 8585 27288
rect 8527 27279 8585 27285
rect 8846 27276 8852 27288
rect 8904 27276 8910 27328
rect 9398 27316 9404 27328
rect 9359 27288 9404 27316
rect 9398 27276 9404 27288
rect 9456 27276 9462 27328
rect 12526 27276 12532 27328
rect 12584 27316 12590 27328
rect 12943 27319 13001 27325
rect 12943 27316 12955 27319
rect 12584 27288 12955 27316
rect 12584 27276 12590 27288
rect 12943 27285 12955 27288
rect 12989 27285 13001 27319
rect 12943 27279 13001 27285
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 3191 27115 3249 27121
rect 3191 27081 3203 27115
rect 3237 27112 3249 27115
rect 5350 27112 5356 27124
rect 3237 27084 5356 27112
rect 3237 27081 3249 27084
rect 3191 27075 3249 27081
rect 5350 27072 5356 27084
rect 5408 27072 5414 27124
rect 6270 27112 6276 27124
rect 6231 27084 6276 27112
rect 6270 27072 6276 27084
rect 6328 27072 6334 27124
rect 7834 27112 7840 27124
rect 7795 27084 7840 27112
rect 7834 27072 7840 27084
rect 7892 27112 7898 27124
rect 8527 27115 8585 27121
rect 8527 27112 8539 27115
rect 7892 27084 8539 27112
rect 7892 27072 7898 27084
rect 8527 27081 8539 27084
rect 8573 27081 8585 27115
rect 11974 27112 11980 27124
rect 11935 27084 11980 27112
rect 8527 27075 8585 27081
rect 11974 27072 11980 27084
rect 12032 27072 12038 27124
rect 12802 27072 12808 27124
rect 12860 27112 12866 27124
rect 13630 27121 13636 27124
rect 13265 27115 13323 27121
rect 13265 27112 13277 27115
rect 12860 27084 13277 27112
rect 12860 27072 12866 27084
rect 13265 27081 13277 27084
rect 13311 27081 13323 27115
rect 13265 27075 13323 27081
rect 13587 27115 13636 27121
rect 13587 27081 13599 27115
rect 13633 27081 13636 27115
rect 13587 27075 13636 27081
rect 13630 27072 13636 27075
rect 13688 27072 13694 27124
rect 4522 27044 4528 27056
rect 4483 27016 4528 27044
rect 4522 27004 4528 27016
rect 4580 27004 4586 27056
rect 5534 27044 5540 27056
rect 4724 27016 5540 27044
rect 4724 26976 4752 27016
rect 5534 27004 5540 27016
rect 5592 27004 5598 27056
rect 5721 27047 5779 27053
rect 5721 27013 5733 27047
rect 5767 27044 5779 27047
rect 5767 27016 7052 27044
rect 5767 27013 5779 27016
rect 5721 27007 5779 27013
rect 7024 26988 7052 27016
rect 8386 27004 8392 27056
rect 8444 27044 8450 27056
rect 8849 27047 8907 27053
rect 8849 27044 8861 27047
rect 8444 27016 8861 27044
rect 8444 27004 8450 27016
rect 8849 27013 8861 27016
rect 8895 27013 8907 27047
rect 10226 27044 10232 27056
rect 10187 27016 10232 27044
rect 8849 27007 8907 27013
rect 10226 27004 10232 27016
rect 10284 27004 10290 27056
rect 3528 26948 4752 26976
rect 2866 26868 2872 26920
rect 2924 26908 2930 26920
rect 3528 26917 3556 26948
rect 4798 26936 4804 26988
rect 4856 26976 4862 26988
rect 5169 26979 5227 26985
rect 5169 26976 5181 26979
rect 4856 26948 5181 26976
rect 4856 26936 4862 26948
rect 5169 26945 5181 26948
rect 5215 26945 5227 26979
rect 6914 26976 6920 26988
rect 6875 26948 6920 26976
rect 5169 26939 5227 26945
rect 6914 26936 6920 26948
rect 6972 26936 6978 26988
rect 7006 26936 7012 26988
rect 7064 26976 7070 26988
rect 7193 26979 7251 26985
rect 7193 26976 7205 26979
rect 7064 26948 7205 26976
rect 7064 26936 7070 26948
rect 7193 26945 7205 26948
rect 7239 26945 7251 26979
rect 7193 26939 7251 26945
rect 9858 26936 9864 26988
rect 9916 26976 9922 26988
rect 10965 26979 11023 26985
rect 10965 26976 10977 26979
rect 9916 26948 10977 26976
rect 9916 26936 9922 26948
rect 10965 26945 10977 26948
rect 11011 26945 11023 26979
rect 10965 26939 11023 26945
rect 11330 26936 11336 26988
rect 11388 26976 11394 26988
rect 12575 26979 12633 26985
rect 12575 26976 12587 26979
rect 11388 26948 12587 26976
rect 11388 26936 11394 26948
rect 12575 26945 12587 26948
rect 12621 26945 12633 26979
rect 12575 26939 12633 26945
rect 4154 26917 4160 26920
rect 3088 26911 3146 26917
rect 3088 26908 3100 26911
rect 2924 26880 3100 26908
rect 2924 26868 2930 26880
rect 3088 26877 3100 26880
rect 3134 26908 3146 26911
rect 3513 26911 3571 26917
rect 3513 26908 3525 26911
rect 3134 26880 3525 26908
rect 3134 26877 3146 26880
rect 3088 26871 3146 26877
rect 3513 26877 3525 26880
rect 3559 26877 3571 26911
rect 4132 26911 4160 26917
rect 4132 26908 4144 26911
rect 4067 26880 4144 26908
rect 3513 26871 3571 26877
rect 4132 26877 4144 26880
rect 4212 26908 4218 26920
rect 4212 26880 5028 26908
rect 4132 26871 4160 26877
rect 4154 26868 4160 26871
rect 4212 26868 4218 26880
rect 4203 26775 4261 26781
rect 4203 26741 4215 26775
rect 4249 26772 4261 26775
rect 4430 26772 4436 26784
rect 4249 26744 4436 26772
rect 4249 26741 4261 26744
rect 4203 26735 4261 26741
rect 4430 26732 4436 26744
rect 4488 26732 4494 26784
rect 5000 26781 5028 26880
rect 6178 26868 6184 26920
rect 6236 26908 6242 26920
rect 6549 26911 6607 26917
rect 6549 26908 6561 26911
rect 6236 26880 6561 26908
rect 6236 26868 6242 26880
rect 6549 26877 6561 26880
rect 6595 26877 6607 26911
rect 6549 26871 6607 26877
rect 5258 26840 5264 26852
rect 5219 26812 5264 26840
rect 5258 26800 5264 26812
rect 5316 26800 5322 26852
rect 4985 26775 5043 26781
rect 4985 26741 4997 26775
rect 5031 26772 5043 26775
rect 5166 26772 5172 26784
rect 5031 26744 5172 26772
rect 5031 26741 5043 26744
rect 4985 26735 5043 26741
rect 5166 26732 5172 26744
rect 5224 26732 5230 26784
rect 6564 26772 6592 26871
rect 8294 26868 8300 26920
rect 8352 26908 8358 26920
rect 8424 26911 8482 26917
rect 8424 26908 8436 26911
rect 8352 26880 8436 26908
rect 8352 26868 8358 26880
rect 8424 26877 8436 26880
rect 8470 26908 8482 26911
rect 9217 26911 9275 26917
rect 9217 26908 9229 26911
rect 8470 26880 9229 26908
rect 8470 26877 8482 26880
rect 8424 26871 8482 26877
rect 9217 26877 9229 26880
rect 9263 26877 9275 26911
rect 9217 26871 9275 26877
rect 11054 26868 11060 26920
rect 11112 26908 11118 26920
rect 11184 26911 11242 26917
rect 11184 26908 11196 26911
rect 11112 26880 11196 26908
rect 11112 26868 11118 26880
rect 11184 26877 11196 26880
rect 11230 26908 11242 26911
rect 11609 26911 11667 26917
rect 11609 26908 11621 26911
rect 11230 26880 11621 26908
rect 11230 26877 11242 26880
rect 11184 26871 11242 26877
rect 11609 26877 11621 26880
rect 11655 26877 11667 26911
rect 11609 26871 11667 26877
rect 12250 26868 12256 26920
rect 12308 26908 12314 26920
rect 12488 26911 12546 26917
rect 12488 26908 12500 26911
rect 12308 26880 12500 26908
rect 12308 26868 12314 26880
rect 12488 26877 12500 26880
rect 12534 26908 12546 26911
rect 12897 26911 12955 26917
rect 12897 26908 12909 26911
rect 12534 26880 12909 26908
rect 12534 26877 12546 26880
rect 12488 26871 12546 26877
rect 12897 26877 12909 26880
rect 12943 26877 12955 26911
rect 13516 26911 13574 26917
rect 13516 26908 13528 26911
rect 12897 26871 12955 26877
rect 13280 26880 13528 26908
rect 7009 26843 7067 26849
rect 7009 26809 7021 26843
rect 7055 26809 7067 26843
rect 9674 26840 9680 26852
rect 9635 26812 9680 26840
rect 7009 26803 7067 26809
rect 7024 26772 7052 26803
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 9766 26800 9772 26852
rect 9824 26840 9830 26852
rect 10597 26843 10655 26849
rect 10597 26840 10609 26843
rect 9824 26812 10609 26840
rect 9824 26800 9830 26812
rect 10597 26809 10609 26812
rect 10643 26809 10655 26843
rect 10597 26803 10655 26809
rect 12066 26800 12072 26852
rect 12124 26840 12130 26852
rect 13280 26840 13308 26880
rect 13516 26877 13528 26880
rect 13562 26908 13574 26911
rect 13909 26911 13967 26917
rect 13909 26908 13921 26911
rect 13562 26880 13921 26908
rect 13562 26877 13574 26880
rect 13516 26871 13574 26877
rect 13909 26877 13921 26880
rect 13955 26877 13967 26911
rect 13909 26871 13967 26877
rect 12124 26812 13308 26840
rect 12124 26800 12130 26812
rect 6564 26744 7052 26772
rect 11054 26732 11060 26784
rect 11112 26772 11118 26784
rect 11287 26775 11345 26781
rect 11287 26772 11299 26775
rect 11112 26744 11299 26772
rect 11112 26732 11118 26744
rect 11287 26741 11299 26744
rect 11333 26741 11345 26775
rect 11287 26735 11345 26741
rect 11974 26732 11980 26784
rect 12032 26772 12038 26784
rect 12710 26772 12716 26784
rect 12032 26744 12716 26772
rect 12032 26732 12038 26744
rect 12710 26732 12716 26744
rect 12768 26732 12774 26784
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 5261 26571 5319 26577
rect 5261 26537 5273 26571
rect 5307 26568 5319 26571
rect 5626 26568 5632 26580
rect 5307 26540 5632 26568
rect 5307 26537 5319 26540
rect 5261 26531 5319 26537
rect 5626 26528 5632 26540
rect 5684 26528 5690 26580
rect 6914 26528 6920 26580
rect 6972 26568 6978 26580
rect 7101 26571 7159 26577
rect 7101 26568 7113 26571
rect 6972 26540 7113 26568
rect 6972 26528 6978 26540
rect 7101 26537 7113 26540
rect 7147 26537 7159 26571
rect 7101 26531 7159 26537
rect 9493 26571 9551 26577
rect 9493 26537 9505 26571
rect 9539 26568 9551 26571
rect 9674 26568 9680 26580
rect 9539 26540 9680 26568
rect 9539 26537 9551 26540
rect 9493 26531 9551 26537
rect 9674 26528 9680 26540
rect 9732 26528 9738 26580
rect 11149 26571 11207 26577
rect 11149 26537 11161 26571
rect 11195 26568 11207 26571
rect 11514 26568 11520 26580
rect 11195 26540 11520 26568
rect 11195 26537 11207 26540
rect 11149 26531 11207 26537
rect 11514 26528 11520 26540
rect 11572 26568 11578 26580
rect 12618 26568 12624 26580
rect 11572 26540 12624 26568
rect 11572 26528 11578 26540
rect 12618 26528 12624 26540
rect 12676 26528 12682 26580
rect 12894 26568 12900 26580
rect 12855 26540 12900 26568
rect 12894 26528 12900 26540
rect 12952 26528 12958 26580
rect 4614 26460 4620 26512
rect 4672 26509 4678 26512
rect 4672 26503 4720 26509
rect 4672 26469 4674 26503
rect 4708 26469 4720 26503
rect 4672 26463 4720 26469
rect 4672 26460 4678 26463
rect 5350 26460 5356 26512
rect 5408 26500 5414 26512
rect 5905 26503 5963 26509
rect 5905 26500 5917 26503
rect 5408 26472 5917 26500
rect 5408 26460 5414 26472
rect 5905 26469 5917 26472
rect 5951 26469 5963 26503
rect 5905 26463 5963 26469
rect 6178 26460 6184 26512
rect 6236 26500 6242 26512
rect 6273 26503 6331 26509
rect 6273 26500 6285 26503
rect 6236 26472 6285 26500
rect 6236 26460 6242 26472
rect 6273 26469 6285 26472
rect 6319 26469 6331 26503
rect 6273 26463 6331 26469
rect 9125 26503 9183 26509
rect 9125 26469 9137 26503
rect 9171 26500 9183 26503
rect 9582 26500 9588 26512
rect 9171 26472 9588 26500
rect 9171 26469 9183 26472
rect 9125 26463 9183 26469
rect 9582 26460 9588 26472
rect 9640 26460 9646 26512
rect 9858 26500 9864 26512
rect 9819 26472 9864 26500
rect 9858 26460 9864 26472
rect 9916 26460 9922 26512
rect 11330 26500 11336 26512
rect 11291 26472 11336 26500
rect 11330 26460 11336 26472
rect 11388 26460 11394 26512
rect 11425 26503 11483 26509
rect 11425 26469 11437 26503
rect 11471 26500 11483 26503
rect 12434 26500 12440 26512
rect 11471 26472 12440 26500
rect 11471 26469 11483 26472
rect 11425 26463 11483 26469
rect 12434 26460 12440 26472
rect 12492 26500 12498 26512
rect 13354 26500 13360 26512
rect 12492 26472 12585 26500
rect 13096 26472 13360 26500
rect 12492 26460 12498 26472
rect 4430 26392 4436 26444
rect 4488 26432 4494 26444
rect 4488 26404 5672 26432
rect 4488 26392 4494 26404
rect 4341 26367 4399 26373
rect 4341 26333 4353 26367
rect 4387 26364 4399 26367
rect 5442 26364 5448 26376
rect 4387 26336 5448 26364
rect 4387 26333 4399 26336
rect 4341 26327 4399 26333
rect 5442 26324 5448 26336
rect 5500 26324 5506 26376
rect 5644 26364 5672 26404
rect 7558 26392 7564 26444
rect 7616 26432 7622 26444
rect 7837 26435 7895 26441
rect 7837 26432 7849 26435
rect 7616 26404 7849 26432
rect 7616 26392 7622 26404
rect 7837 26401 7849 26404
rect 7883 26401 7895 26435
rect 8294 26432 8300 26444
rect 8255 26404 8300 26432
rect 7837 26395 7895 26401
rect 8294 26392 8300 26404
rect 8352 26392 8358 26444
rect 13096 26441 13124 26472
rect 13354 26460 13360 26472
rect 13412 26460 13418 26512
rect 10413 26435 10471 26441
rect 10413 26401 10425 26435
rect 10459 26432 10471 26435
rect 13081 26435 13139 26441
rect 10459 26404 11192 26432
rect 10459 26401 10471 26404
rect 10413 26395 10471 26401
rect 11164 26376 11192 26404
rect 13081 26401 13093 26435
rect 13127 26401 13139 26435
rect 13081 26395 13139 26401
rect 13265 26435 13323 26441
rect 13265 26401 13277 26435
rect 13311 26401 13323 26435
rect 13265 26395 13323 26401
rect 6181 26367 6239 26373
rect 6181 26364 6193 26367
rect 5644 26336 6193 26364
rect 6181 26333 6193 26336
rect 6227 26364 6239 26367
rect 6454 26364 6460 26376
rect 6227 26336 6460 26364
rect 6227 26333 6239 26336
rect 6181 26327 6239 26333
rect 6454 26324 6460 26336
rect 6512 26324 6518 26376
rect 8386 26364 8392 26376
rect 8347 26336 8392 26364
rect 8386 26324 8392 26336
rect 8444 26324 8450 26376
rect 9769 26367 9827 26373
rect 9769 26333 9781 26367
rect 9815 26364 9827 26367
rect 9950 26364 9956 26376
rect 9815 26336 9956 26364
rect 9815 26333 9827 26336
rect 9769 26327 9827 26333
rect 9950 26324 9956 26336
rect 10008 26364 10014 26376
rect 11054 26364 11060 26376
rect 10008 26336 11060 26364
rect 10008 26324 10014 26336
rect 11054 26324 11060 26336
rect 11112 26324 11118 26376
rect 11146 26324 11152 26376
rect 11204 26364 11210 26376
rect 11609 26367 11667 26373
rect 11609 26364 11621 26367
rect 11204 26336 11621 26364
rect 11204 26324 11210 26336
rect 11609 26333 11621 26336
rect 11655 26333 11667 26367
rect 11609 26327 11667 26333
rect 11974 26324 11980 26376
rect 12032 26364 12038 26376
rect 12802 26364 12808 26376
rect 12032 26336 12808 26364
rect 12032 26324 12038 26336
rect 12802 26324 12808 26336
rect 12860 26364 12866 26376
rect 13280 26364 13308 26395
rect 12860 26336 13308 26364
rect 12860 26324 12866 26336
rect 5626 26256 5632 26308
rect 5684 26296 5690 26308
rect 6733 26299 6791 26305
rect 6733 26296 6745 26299
rect 5684 26268 6745 26296
rect 5684 26256 5690 26268
rect 6733 26265 6745 26268
rect 6779 26265 6791 26299
rect 6733 26259 6791 26265
rect 7561 26231 7619 26237
rect 7561 26197 7573 26231
rect 7607 26228 7619 26231
rect 7650 26228 7656 26240
rect 7607 26200 7656 26228
rect 7607 26197 7619 26200
rect 7561 26191 7619 26197
rect 7650 26188 7656 26200
rect 7708 26188 7714 26240
rect 10042 26188 10048 26240
rect 10100 26228 10106 26240
rect 10689 26231 10747 26237
rect 10689 26228 10701 26231
rect 10100 26200 10701 26228
rect 10100 26188 10106 26200
rect 10689 26197 10701 26200
rect 10735 26197 10747 26231
rect 10689 26191 10747 26197
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 5169 26027 5227 26033
rect 5169 25993 5181 26027
rect 5215 26024 5227 26027
rect 5258 26024 5264 26036
rect 5215 25996 5264 26024
rect 5215 25993 5227 25996
rect 5169 25987 5227 25993
rect 5258 25984 5264 25996
rect 5316 25984 5322 26036
rect 6454 26024 6460 26036
rect 6415 25996 6460 26024
rect 6454 25984 6460 25996
rect 6512 25984 6518 26036
rect 7469 26027 7527 26033
rect 7469 25993 7481 26027
rect 7515 26024 7527 26027
rect 8294 26024 8300 26036
rect 7515 25996 8300 26024
rect 7515 25993 7527 25996
rect 7469 25987 7527 25993
rect 8294 25984 8300 25996
rect 8352 25984 8358 26036
rect 9217 26027 9275 26033
rect 9217 25993 9229 26027
rect 9263 26024 9275 26027
rect 9306 26024 9312 26036
rect 9263 25996 9312 26024
rect 9263 25993 9275 25996
rect 9217 25987 9275 25993
rect 9306 25984 9312 25996
rect 9364 26024 9370 26036
rect 9490 26024 9496 26036
rect 9364 25996 9496 26024
rect 9364 25984 9370 25996
rect 9490 25984 9496 25996
rect 9548 25984 9554 26036
rect 9585 26027 9643 26033
rect 9585 25993 9597 26027
rect 9631 26024 9643 26027
rect 9858 26024 9864 26036
rect 9631 25996 9864 26024
rect 9631 25993 9643 25996
rect 9585 25987 9643 25993
rect 9858 25984 9864 25996
rect 9916 26024 9922 26036
rect 10965 26027 11023 26033
rect 10965 26024 10977 26027
rect 9916 25996 10977 26024
rect 9916 25984 9922 25996
rect 10965 25993 10977 25996
rect 11011 25993 11023 26027
rect 10965 25987 11023 25993
rect 11330 25984 11336 26036
rect 11388 26024 11394 26036
rect 11609 26027 11667 26033
rect 11609 26024 11621 26027
rect 11388 25996 11621 26024
rect 11388 25984 11394 25996
rect 11609 25993 11621 25996
rect 11655 25993 11667 26027
rect 11609 25987 11667 25993
rect 6914 25916 6920 25968
rect 6972 25965 6978 25968
rect 6972 25959 7021 25965
rect 6972 25925 6975 25959
rect 7009 25925 7021 25959
rect 6972 25919 7021 25925
rect 6972 25916 6978 25919
rect 7926 25916 7932 25968
rect 7984 25956 7990 25968
rect 8113 25959 8171 25965
rect 8113 25956 8125 25959
rect 7984 25928 8125 25956
rect 7984 25916 7990 25928
rect 8113 25925 8125 25928
rect 8159 25956 8171 25959
rect 9953 25959 10011 25965
rect 9953 25956 9965 25959
rect 8159 25928 9965 25956
rect 8159 25925 8171 25928
rect 8113 25919 8171 25925
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25888 8355 25891
rect 8386 25888 8392 25900
rect 8343 25860 8392 25888
rect 8343 25857 8355 25860
rect 8297 25851 8355 25857
rect 8386 25848 8392 25860
rect 8444 25848 8450 25900
rect 4249 25823 4307 25829
rect 4249 25820 4261 25823
rect 3988 25792 4261 25820
rect 3988 25696 4016 25792
rect 4249 25789 4261 25792
rect 4295 25789 4307 25823
rect 4249 25783 4307 25789
rect 6892 25823 6950 25829
rect 6892 25789 6904 25823
rect 6938 25820 6950 25823
rect 7650 25820 7656 25832
rect 6938 25792 7656 25820
rect 6938 25789 6950 25792
rect 6892 25783 6950 25789
rect 7650 25780 7656 25792
rect 7708 25780 7714 25832
rect 4614 25761 4620 25764
rect 4157 25755 4215 25761
rect 4157 25721 4169 25755
rect 4203 25752 4215 25755
rect 4611 25752 4620 25761
rect 4203 25724 4620 25752
rect 4203 25721 4215 25724
rect 4157 25715 4215 25721
rect 4611 25715 4620 25724
rect 4614 25712 4620 25715
rect 4672 25712 4678 25764
rect 8680 25761 8708 25928
rect 9953 25925 9965 25928
rect 9999 25925 10011 25959
rect 9953 25919 10011 25925
rect 9968 25888 9996 25919
rect 12526 25888 12532 25900
rect 9968 25860 10180 25888
rect 12487 25860 12532 25888
rect 10042 25820 10048 25832
rect 10003 25792 10048 25820
rect 10042 25780 10048 25792
rect 10100 25780 10106 25832
rect 8659 25755 8717 25761
rect 8659 25721 8671 25755
rect 8705 25721 8717 25755
rect 10152 25752 10180 25860
rect 12526 25848 12532 25860
rect 12584 25848 12590 25900
rect 12618 25848 12624 25900
rect 12676 25888 12682 25900
rect 12805 25891 12863 25897
rect 12805 25888 12817 25891
rect 12676 25860 12817 25888
rect 12676 25848 12682 25860
rect 12805 25857 12817 25860
rect 12851 25857 12863 25891
rect 12805 25851 12863 25857
rect 10962 25780 10968 25832
rect 11020 25820 11026 25832
rect 11333 25823 11391 25829
rect 11333 25820 11345 25823
rect 11020 25792 11345 25820
rect 11020 25780 11026 25792
rect 11333 25789 11345 25792
rect 11379 25820 11391 25823
rect 11379 25792 12296 25820
rect 11379 25789 11391 25792
rect 11333 25783 11391 25789
rect 10366 25755 10424 25761
rect 10366 25752 10378 25755
rect 10152 25724 10378 25752
rect 8659 25715 8717 25721
rect 10366 25721 10378 25724
rect 10412 25752 10424 25755
rect 10502 25752 10508 25764
rect 10412 25724 10508 25752
rect 10412 25721 10424 25724
rect 10366 25715 10424 25721
rect 10502 25712 10508 25724
rect 10560 25712 10566 25764
rect 3789 25687 3847 25693
rect 3789 25653 3801 25687
rect 3835 25684 3847 25687
rect 3970 25684 3976 25696
rect 3835 25656 3976 25684
rect 3835 25653 3847 25656
rect 3789 25647 3847 25653
rect 3970 25644 3976 25656
rect 4028 25644 4034 25696
rect 5534 25684 5540 25696
rect 5495 25656 5540 25684
rect 5534 25644 5540 25656
rect 5592 25644 5598 25696
rect 6086 25684 6092 25696
rect 6047 25656 6092 25684
rect 6086 25644 6092 25656
rect 6144 25644 6150 25696
rect 7558 25644 7564 25696
rect 7616 25684 7622 25696
rect 7745 25687 7803 25693
rect 7745 25684 7757 25687
rect 7616 25656 7757 25684
rect 7616 25644 7622 25656
rect 7745 25653 7757 25656
rect 7791 25653 7803 25687
rect 7745 25647 7803 25653
rect 11974 25644 11980 25696
rect 12032 25684 12038 25696
rect 12161 25687 12219 25693
rect 12161 25684 12173 25687
rect 12032 25656 12173 25684
rect 12032 25644 12038 25656
rect 12161 25653 12173 25656
rect 12207 25653 12219 25687
rect 12268 25684 12296 25792
rect 12621 25755 12679 25761
rect 12621 25721 12633 25755
rect 12667 25721 12679 25755
rect 12621 25715 12679 25721
rect 12434 25684 12440 25696
rect 12268 25656 12440 25684
rect 12161 25647 12219 25653
rect 12434 25644 12440 25656
rect 12492 25684 12498 25696
rect 12636 25684 12664 25715
rect 12492 25656 12664 25684
rect 12492 25644 12498 25656
rect 13354 25644 13360 25696
rect 13412 25684 13418 25696
rect 13449 25687 13507 25693
rect 13449 25684 13461 25687
rect 13412 25656 13461 25684
rect 13412 25644 13418 25656
rect 13449 25653 13461 25656
rect 13495 25653 13507 25687
rect 13449 25647 13507 25653
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 5813 25483 5871 25489
rect 5813 25449 5825 25483
rect 5859 25480 5871 25483
rect 6086 25480 6092 25492
rect 5859 25452 6092 25480
rect 5859 25449 5871 25452
rect 5813 25443 5871 25449
rect 6086 25440 6092 25452
rect 6144 25440 6150 25492
rect 8386 25480 8392 25492
rect 8347 25452 8392 25480
rect 8386 25440 8392 25452
rect 8444 25440 8450 25492
rect 8846 25440 8852 25492
rect 8904 25480 8910 25492
rect 8941 25483 8999 25489
rect 8941 25480 8953 25483
rect 8904 25452 8953 25480
rect 8904 25440 8910 25452
rect 8941 25449 8953 25452
rect 8987 25449 8999 25483
rect 9950 25480 9956 25492
rect 9911 25452 9956 25480
rect 8941 25443 8999 25449
rect 9950 25440 9956 25452
rect 10008 25440 10014 25492
rect 10962 25480 10968 25492
rect 10923 25452 10968 25480
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 11974 25440 11980 25492
rect 12032 25480 12038 25492
rect 12434 25480 12440 25492
rect 12032 25452 12440 25480
rect 12032 25440 12038 25452
rect 12434 25440 12440 25452
rect 12492 25440 12498 25492
rect 12526 25440 12532 25492
rect 12584 25480 12590 25492
rect 12989 25483 13047 25489
rect 12989 25480 13001 25483
rect 12584 25452 13001 25480
rect 12584 25440 12590 25452
rect 12989 25449 13001 25452
rect 13035 25449 13047 25483
rect 12989 25443 13047 25449
rect 13262 25440 13268 25492
rect 13320 25480 13326 25492
rect 13679 25483 13737 25489
rect 13679 25480 13691 25483
rect 13320 25452 13691 25480
rect 13320 25440 13326 25452
rect 13679 25449 13691 25452
rect 13725 25449 13737 25483
rect 13679 25443 13737 25449
rect 3142 25412 3148 25424
rect 3103 25384 3148 25412
rect 3142 25372 3148 25384
rect 3200 25372 3206 25424
rect 4341 25415 4399 25421
rect 4341 25381 4353 25415
rect 4387 25412 4399 25415
rect 4614 25412 4620 25424
rect 4387 25384 4620 25412
rect 4387 25381 4399 25384
rect 4341 25375 4399 25381
rect 4614 25372 4620 25384
rect 4672 25412 4678 25424
rect 5258 25421 5264 25424
rect 5255 25412 5264 25421
rect 4672 25384 5264 25412
rect 4672 25372 4678 25384
rect 5255 25375 5264 25384
rect 5258 25372 5264 25375
rect 5316 25372 5322 25424
rect 7098 25421 7104 25424
rect 7095 25412 7104 25421
rect 7011 25384 7104 25412
rect 7095 25375 7104 25384
rect 7156 25412 7162 25424
rect 7926 25412 7932 25424
rect 7156 25384 7932 25412
rect 7098 25372 7104 25375
rect 7156 25372 7162 25384
rect 7926 25372 7932 25384
rect 7984 25372 7990 25424
rect 10407 25415 10465 25421
rect 10407 25381 10419 25415
rect 10453 25412 10465 25415
rect 10502 25412 10508 25424
rect 10453 25384 10508 25412
rect 10453 25381 10465 25384
rect 10407 25375 10465 25381
rect 10502 25372 10508 25384
rect 10560 25412 10566 25424
rect 11790 25412 11796 25424
rect 10560 25384 11796 25412
rect 10560 25372 10566 25384
rect 11790 25372 11796 25384
rect 11848 25412 11854 25424
rect 12114 25415 12172 25421
rect 12114 25412 12126 25415
rect 11848 25384 12126 25412
rect 11848 25372 11854 25384
rect 12114 25381 12126 25384
rect 12160 25381 12172 25415
rect 12114 25375 12172 25381
rect 2682 25344 2688 25356
rect 2643 25316 2688 25344
rect 2682 25304 2688 25316
rect 2740 25304 2746 25356
rect 2958 25344 2964 25356
rect 2919 25316 2964 25344
rect 2958 25304 2964 25316
rect 3016 25304 3022 25356
rect 10045 25347 10103 25353
rect 10045 25313 10057 25347
rect 10091 25344 10103 25347
rect 10134 25344 10140 25356
rect 10091 25316 10140 25344
rect 10091 25313 10103 25316
rect 10045 25307 10103 25313
rect 10134 25304 10140 25316
rect 10192 25304 10198 25356
rect 12710 25344 12716 25356
rect 12671 25316 12716 25344
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 13446 25304 13452 25356
rect 13504 25344 13510 25356
rect 13576 25347 13634 25353
rect 13576 25344 13588 25347
rect 13504 25316 13588 25344
rect 13504 25304 13510 25316
rect 13576 25313 13588 25316
rect 13622 25313 13634 25347
rect 13576 25307 13634 25313
rect 4893 25279 4951 25285
rect 4893 25245 4905 25279
rect 4939 25245 4951 25279
rect 6733 25279 6791 25285
rect 6733 25276 6745 25279
rect 4893 25239 4951 25245
rect 6564 25248 6745 25276
rect 4154 25168 4160 25220
rect 4212 25208 4218 25220
rect 4709 25211 4767 25217
rect 4709 25208 4721 25211
rect 4212 25180 4721 25208
rect 4212 25168 4218 25180
rect 4709 25177 4721 25180
rect 4755 25208 4767 25211
rect 4908 25208 4936 25239
rect 4755 25180 4936 25208
rect 4755 25177 4767 25180
rect 4709 25171 4767 25177
rect 5902 25100 5908 25152
rect 5960 25140 5966 25152
rect 6564 25149 6592 25248
rect 6733 25245 6745 25248
rect 6779 25245 6791 25279
rect 8478 25276 8484 25288
rect 8439 25248 8484 25276
rect 6733 25239 6791 25245
rect 8478 25236 8484 25248
rect 8536 25236 8542 25288
rect 11793 25279 11851 25285
rect 11793 25245 11805 25279
rect 11839 25276 11851 25279
rect 11974 25276 11980 25288
rect 11839 25248 11980 25276
rect 11839 25245 11851 25248
rect 11793 25239 11851 25245
rect 11974 25236 11980 25248
rect 12032 25236 12038 25288
rect 6549 25143 6607 25149
rect 6549 25140 6561 25143
rect 5960 25112 6561 25140
rect 5960 25100 5966 25112
rect 6549 25109 6561 25112
rect 6595 25109 6607 25143
rect 6549 25103 6607 25109
rect 7282 25100 7288 25152
rect 7340 25140 7346 25152
rect 7653 25143 7711 25149
rect 7653 25140 7665 25143
rect 7340 25112 7665 25140
rect 7340 25100 7346 25112
rect 7653 25109 7665 25112
rect 7699 25140 7711 25143
rect 7929 25143 7987 25149
rect 7929 25140 7941 25143
rect 7699 25112 7941 25140
rect 7699 25109 7711 25112
rect 7653 25103 7711 25109
rect 7929 25109 7941 25112
rect 7975 25109 7987 25143
rect 7929 25103 7987 25109
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 2501 24939 2559 24945
rect 2501 24905 2513 24939
rect 2547 24936 2559 24939
rect 2682 24936 2688 24948
rect 2547 24908 2688 24936
rect 2547 24905 2559 24908
rect 2501 24899 2559 24905
rect 2682 24896 2688 24908
rect 2740 24896 2746 24948
rect 2869 24939 2927 24945
rect 2869 24905 2881 24939
rect 2915 24936 2927 24939
rect 2958 24936 2964 24948
rect 2915 24908 2964 24936
rect 2915 24905 2927 24908
rect 2869 24899 2927 24905
rect 2958 24896 2964 24908
rect 3016 24896 3022 24948
rect 8205 24939 8263 24945
rect 8205 24905 8217 24939
rect 8251 24936 8263 24939
rect 8478 24936 8484 24948
rect 8251 24908 8484 24936
rect 8251 24905 8263 24908
rect 8205 24899 8263 24905
rect 5902 24800 5908 24812
rect 5863 24772 5908 24800
rect 5902 24760 5908 24772
rect 5960 24760 5966 24812
rect 5994 24760 6000 24812
rect 6052 24800 6058 24812
rect 6181 24803 6239 24809
rect 6181 24800 6193 24803
rect 6052 24772 6193 24800
rect 6052 24760 6058 24772
rect 6181 24769 6193 24772
rect 6227 24800 6239 24803
rect 7006 24800 7012 24812
rect 6227 24772 7012 24800
rect 6227 24769 6239 24772
rect 6181 24763 6239 24769
rect 7006 24760 7012 24772
rect 7064 24760 7070 24812
rect 7193 24803 7251 24809
rect 7193 24769 7205 24803
rect 7239 24800 7251 24803
rect 8220 24800 8248 24899
rect 8478 24896 8484 24908
rect 8536 24896 8542 24948
rect 10042 24936 10048 24948
rect 9955 24908 10048 24936
rect 10042 24896 10048 24908
rect 10100 24936 10106 24948
rect 10321 24939 10379 24945
rect 10321 24936 10333 24939
rect 10100 24908 10333 24936
rect 10100 24896 10106 24908
rect 10321 24905 10333 24908
rect 10367 24936 10379 24939
rect 10502 24936 10508 24948
rect 10367 24908 10508 24936
rect 10367 24905 10379 24908
rect 10321 24899 10379 24905
rect 8846 24800 8852 24812
rect 7239 24772 8248 24800
rect 8807 24772 8852 24800
rect 7239 24769 7251 24772
rect 7193 24763 7251 24769
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 9490 24800 9496 24812
rect 9451 24772 9496 24800
rect 9490 24760 9496 24772
rect 9548 24760 9554 24812
rect 3605 24735 3663 24741
rect 3605 24732 3617 24735
rect 3436 24704 3617 24732
rect 3050 24556 3056 24608
rect 3108 24596 3114 24608
rect 3436 24605 3464 24704
rect 3605 24701 3617 24704
rect 3651 24701 3663 24735
rect 3605 24695 3663 24701
rect 4157 24735 4215 24741
rect 4157 24701 4169 24735
rect 4203 24732 4215 24735
rect 4246 24732 4252 24744
rect 4203 24704 4252 24732
rect 4203 24701 4215 24704
rect 4157 24695 4215 24701
rect 4246 24692 4252 24704
rect 4304 24692 4310 24744
rect 5445 24735 5503 24741
rect 5445 24701 5457 24735
rect 5491 24701 5503 24735
rect 5445 24695 5503 24701
rect 5460 24664 5488 24695
rect 5534 24692 5540 24744
rect 5592 24732 5598 24744
rect 5629 24735 5687 24741
rect 5629 24732 5641 24735
rect 5592 24704 5641 24732
rect 5592 24692 5598 24704
rect 5629 24701 5641 24704
rect 5675 24701 5687 24735
rect 5629 24695 5687 24701
rect 6012 24664 6040 24760
rect 5460 24636 6040 24664
rect 7282 24624 7288 24676
rect 7340 24664 7346 24676
rect 7340 24636 7385 24664
rect 7340 24624 7346 24636
rect 7650 24624 7656 24676
rect 7708 24664 7714 24676
rect 7837 24667 7895 24673
rect 7837 24664 7849 24667
rect 7708 24636 7849 24664
rect 7708 24624 7714 24636
rect 7837 24633 7849 24636
rect 7883 24633 7895 24667
rect 7837 24627 7895 24633
rect 8665 24667 8723 24673
rect 8665 24633 8677 24667
rect 8711 24664 8723 24667
rect 8941 24667 8999 24673
rect 8941 24664 8953 24667
rect 8711 24636 8953 24664
rect 8711 24633 8723 24636
rect 8665 24627 8723 24633
rect 8941 24633 8953 24636
rect 8987 24664 8999 24667
rect 9306 24664 9312 24676
rect 8987 24636 9312 24664
rect 8987 24633 8999 24636
rect 8941 24627 8999 24633
rect 9306 24624 9312 24636
rect 9364 24624 9370 24676
rect 10428 24664 10456 24908
rect 10502 24896 10508 24908
rect 10560 24896 10566 24948
rect 11790 24936 11796 24948
rect 11751 24908 11796 24936
rect 11790 24896 11796 24908
rect 11848 24896 11854 24948
rect 13446 24896 13452 24948
rect 13504 24936 13510 24948
rect 13541 24939 13599 24945
rect 13541 24936 13553 24939
rect 13504 24908 13553 24936
rect 13504 24896 13510 24908
rect 13541 24905 13553 24908
rect 13587 24905 13599 24939
rect 13541 24899 13599 24905
rect 12526 24868 12532 24880
rect 12176 24840 12532 24868
rect 10778 24760 10784 24812
rect 10836 24800 10842 24812
rect 12176 24809 12204 24840
rect 12526 24828 12532 24840
rect 12584 24868 12590 24880
rect 13354 24868 13360 24880
rect 12584 24840 13360 24868
rect 12584 24828 12590 24840
rect 13354 24828 13360 24840
rect 13412 24828 13418 24880
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 10836 24772 12173 24800
rect 10836 24760 10842 24772
rect 12161 24769 12173 24772
rect 12207 24769 12219 24803
rect 12161 24763 12219 24769
rect 10505 24735 10563 24741
rect 10505 24701 10517 24735
rect 10551 24732 10563 24735
rect 10962 24732 10968 24744
rect 10551 24704 10968 24732
rect 10551 24701 10563 24704
rect 10505 24695 10563 24701
rect 10962 24692 10968 24704
rect 11020 24692 11026 24744
rect 12526 24732 12532 24744
rect 12487 24704 12532 24732
rect 12526 24692 12532 24704
rect 12584 24692 12590 24744
rect 12894 24732 12900 24744
rect 12855 24704 12900 24732
rect 12894 24692 12900 24704
rect 12952 24692 12958 24744
rect 10826 24667 10884 24673
rect 10826 24664 10838 24667
rect 10428 24636 10838 24664
rect 10826 24633 10838 24636
rect 10872 24633 10884 24667
rect 10826 24627 10884 24633
rect 3421 24599 3479 24605
rect 3421 24596 3433 24599
rect 3108 24568 3433 24596
rect 3108 24556 3114 24568
rect 3421 24565 3433 24568
rect 3467 24565 3479 24599
rect 3421 24559 3479 24565
rect 3881 24599 3939 24605
rect 3881 24565 3893 24599
rect 3927 24596 3939 24599
rect 3970 24596 3976 24608
rect 3927 24568 3976 24596
rect 3927 24565 3939 24568
rect 3881 24559 3939 24565
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 4985 24599 5043 24605
rect 4985 24565 4997 24599
rect 5031 24596 5043 24599
rect 5258 24596 5264 24608
rect 5031 24568 5264 24596
rect 5031 24565 5043 24568
rect 4985 24559 5043 24565
rect 5258 24556 5264 24568
rect 5316 24596 5322 24608
rect 6638 24596 6644 24608
rect 5316 24568 6644 24596
rect 5316 24556 5322 24568
rect 6638 24556 6644 24568
rect 6696 24596 6702 24608
rect 7098 24596 7104 24608
rect 6696 24568 7104 24596
rect 6696 24556 6702 24568
rect 7098 24556 7104 24568
rect 7156 24556 7162 24608
rect 11238 24556 11244 24608
rect 11296 24596 11302 24608
rect 11425 24599 11483 24605
rect 11425 24596 11437 24599
rect 11296 24568 11437 24596
rect 11296 24556 11302 24568
rect 11425 24565 11437 24568
rect 11471 24565 11483 24599
rect 12526 24596 12532 24608
rect 12487 24568 12532 24596
rect 11425 24559 11483 24565
rect 12526 24556 12532 24568
rect 12584 24556 12590 24608
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 8754 24392 8760 24404
rect 8715 24364 8760 24392
rect 8754 24352 8760 24364
rect 8812 24352 8818 24404
rect 10134 24352 10140 24404
rect 10192 24392 10198 24404
rect 10505 24395 10563 24401
rect 10505 24392 10517 24395
rect 10192 24364 10517 24392
rect 10192 24352 10198 24364
rect 10505 24361 10517 24364
rect 10551 24361 10563 24395
rect 10505 24355 10563 24361
rect 12529 24395 12587 24401
rect 12529 24361 12541 24395
rect 12575 24392 12587 24395
rect 12894 24392 12900 24404
rect 12575 24364 12900 24392
rect 12575 24361 12587 24364
rect 12529 24355 12587 24361
rect 12894 24352 12900 24364
rect 12952 24352 12958 24404
rect 4801 24327 4859 24333
rect 4801 24293 4813 24327
rect 4847 24324 4859 24327
rect 5442 24324 5448 24336
rect 4847 24296 5448 24324
rect 4847 24293 4859 24296
rect 4801 24287 4859 24293
rect 5442 24284 5448 24296
rect 5500 24284 5506 24336
rect 6549 24327 6607 24333
rect 6549 24293 6561 24327
rect 6595 24324 6607 24327
rect 7193 24327 7251 24333
rect 7193 24324 7205 24327
rect 6595 24296 7205 24324
rect 6595 24293 6607 24296
rect 6549 24287 6607 24293
rect 7193 24293 7205 24296
rect 7239 24324 7251 24327
rect 7282 24324 7288 24336
rect 7239 24296 7288 24324
rect 7239 24293 7251 24296
rect 7193 24287 7251 24293
rect 7282 24284 7288 24296
rect 7340 24284 7346 24336
rect 10229 24327 10287 24333
rect 10229 24293 10241 24327
rect 10275 24324 10287 24327
rect 10410 24324 10416 24336
rect 10275 24296 10416 24324
rect 10275 24293 10287 24296
rect 10229 24287 10287 24293
rect 10410 24284 10416 24296
rect 10468 24284 10474 24336
rect 10962 24324 10968 24336
rect 10923 24296 10968 24324
rect 10962 24284 10968 24296
rect 11020 24284 11026 24336
rect 11238 24324 11244 24336
rect 11199 24296 11244 24324
rect 11238 24284 11244 24296
rect 11296 24284 11302 24336
rect 12759 24327 12817 24333
rect 12759 24293 12771 24327
rect 12805 24324 12817 24327
rect 12986 24324 12992 24336
rect 12805 24296 12992 24324
rect 12805 24293 12817 24296
rect 12759 24287 12817 24293
rect 12986 24284 12992 24296
rect 13044 24284 13050 24336
rect 2961 24259 3019 24265
rect 2961 24225 2973 24259
rect 3007 24256 3019 24259
rect 3142 24256 3148 24268
rect 3007 24228 3148 24256
rect 3007 24225 3019 24228
rect 2961 24219 3019 24225
rect 3142 24216 3148 24228
rect 3200 24216 3206 24268
rect 4065 24259 4123 24265
rect 4065 24225 4077 24259
rect 4111 24225 4123 24259
rect 4065 24219 4123 24225
rect 4080 24188 4108 24219
rect 4246 24216 4252 24268
rect 4304 24256 4310 24268
rect 4525 24259 4583 24265
rect 4525 24256 4537 24259
rect 4304 24228 4537 24256
rect 4304 24216 4310 24228
rect 4525 24225 4537 24228
rect 4571 24225 4583 24259
rect 4525 24219 4583 24225
rect 5997 24259 6055 24265
rect 5997 24225 6009 24259
rect 6043 24256 6055 24259
rect 6270 24256 6276 24268
rect 6043 24228 6276 24256
rect 6043 24225 6055 24228
rect 5997 24219 6055 24225
rect 6270 24216 6276 24228
rect 6328 24216 6334 24268
rect 8386 24216 8392 24268
rect 8444 24256 8450 24268
rect 8573 24259 8631 24265
rect 8573 24256 8585 24259
rect 8444 24228 8585 24256
rect 8444 24216 8450 24228
rect 8573 24225 8585 24228
rect 8619 24225 8631 24259
rect 9674 24256 9680 24268
rect 9635 24228 9680 24256
rect 8573 24219 8631 24225
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 12618 24216 12624 24268
rect 12676 24265 12682 24268
rect 12676 24259 12714 24265
rect 12702 24225 12714 24259
rect 12676 24219 12714 24225
rect 12676 24216 12682 24219
rect 4706 24188 4712 24200
rect 4080 24160 4712 24188
rect 4706 24148 4712 24160
rect 4764 24148 4770 24200
rect 7101 24191 7159 24197
rect 7101 24157 7113 24191
rect 7147 24188 7159 24191
rect 7926 24188 7932 24200
rect 7147 24160 7932 24188
rect 7147 24157 7159 24160
rect 7101 24151 7159 24157
rect 7926 24148 7932 24160
rect 7984 24148 7990 24200
rect 11146 24188 11152 24200
rect 11107 24160 11152 24188
rect 11146 24148 11152 24160
rect 11204 24148 11210 24200
rect 11514 24188 11520 24200
rect 11475 24160 11520 24188
rect 11514 24148 11520 24160
rect 11572 24188 11578 24200
rect 12066 24188 12072 24200
rect 11572 24160 12072 24188
rect 11572 24148 11578 24160
rect 12066 24148 12072 24160
rect 12124 24148 12130 24200
rect 5442 24080 5448 24132
rect 5500 24120 5506 24132
rect 6181 24123 6239 24129
rect 6181 24120 6193 24123
rect 5500 24092 6193 24120
rect 5500 24080 5506 24092
rect 6181 24089 6193 24092
rect 6227 24089 6239 24123
rect 7650 24120 7656 24132
rect 7611 24092 7656 24120
rect 6181 24083 6239 24089
rect 7650 24080 7656 24092
rect 7708 24080 7714 24132
rect 8662 24080 8668 24132
rect 8720 24120 8726 24132
rect 9033 24123 9091 24129
rect 9033 24120 9045 24123
rect 8720 24092 9045 24120
rect 8720 24080 8726 24092
rect 9033 24089 9045 24092
rect 9079 24089 9091 24123
rect 9858 24120 9864 24132
rect 9819 24092 9864 24120
rect 9033 24083 9091 24089
rect 9858 24080 9864 24092
rect 9916 24080 9922 24132
rect 3050 24012 3056 24064
rect 3108 24052 3114 24064
rect 3145 24055 3203 24061
rect 3145 24052 3157 24055
rect 3108 24024 3157 24052
rect 3108 24012 3114 24024
rect 3145 24021 3157 24024
rect 3191 24021 3203 24055
rect 3145 24015 3203 24021
rect 3697 24055 3755 24061
rect 3697 24021 3709 24055
rect 3743 24052 3755 24055
rect 4246 24052 4252 24064
rect 3743 24024 4252 24052
rect 3743 24021 3755 24024
rect 3697 24015 3755 24021
rect 4246 24012 4252 24024
rect 4304 24012 4310 24064
rect 5261 24055 5319 24061
rect 5261 24021 5273 24055
rect 5307 24052 5319 24055
rect 5534 24052 5540 24064
rect 5307 24024 5540 24052
rect 5307 24021 5319 24024
rect 5261 24015 5319 24021
rect 5534 24012 5540 24024
rect 5592 24012 5598 24064
rect 6822 24052 6828 24064
rect 6783 24024 6828 24052
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 10870 24012 10876 24064
rect 10928 24052 10934 24064
rect 11974 24052 11980 24064
rect 10928 24024 11980 24052
rect 10928 24012 10934 24024
rect 11974 24012 11980 24024
rect 12032 24052 12038 24064
rect 12069 24055 12127 24061
rect 12069 24052 12081 24055
rect 12032 24024 12081 24052
rect 12032 24012 12038 24024
rect 12069 24021 12081 24024
rect 12115 24021 12127 24055
rect 12069 24015 12127 24021
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 2501 23851 2559 23857
rect 2501 23817 2513 23851
rect 2547 23848 2559 23851
rect 3142 23848 3148 23860
rect 2547 23820 3148 23848
rect 2547 23817 2559 23820
rect 2501 23811 2559 23817
rect 3142 23808 3148 23820
rect 3200 23808 3206 23860
rect 6638 23848 6644 23860
rect 6599 23820 6644 23848
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 11238 23848 11244 23860
rect 11199 23820 11244 23848
rect 11238 23808 11244 23820
rect 11296 23808 11302 23860
rect 2777 23783 2835 23789
rect 2777 23749 2789 23783
rect 2823 23780 2835 23783
rect 4706 23780 4712 23792
rect 2823 23752 4712 23780
rect 2823 23749 2835 23752
rect 2777 23743 2835 23749
rect 4706 23740 4712 23752
rect 4764 23740 4770 23792
rect 11146 23740 11152 23792
rect 11204 23780 11210 23792
rect 11517 23783 11575 23789
rect 11517 23780 11529 23783
rect 11204 23752 11529 23780
rect 11204 23740 11210 23752
rect 11517 23749 11529 23752
rect 11563 23749 11575 23783
rect 11517 23743 11575 23749
rect 7650 23672 7656 23724
rect 7708 23712 7714 23724
rect 8941 23715 8999 23721
rect 8941 23712 8953 23715
rect 7708 23684 8953 23712
rect 7708 23672 7714 23684
rect 8941 23681 8953 23684
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 10410 23672 10416 23724
rect 10468 23672 10474 23724
rect 10870 23712 10876 23724
rect 10831 23684 10876 23712
rect 10870 23672 10876 23684
rect 10928 23672 10934 23724
rect 2593 23647 2651 23653
rect 2593 23613 2605 23647
rect 2639 23613 2651 23647
rect 3605 23647 3663 23653
rect 3605 23644 3617 23647
rect 2593 23607 2651 23613
rect 3436 23616 3617 23644
rect 2608 23576 2636 23607
rect 3053 23579 3111 23585
rect 3053 23576 3065 23579
rect 2608 23548 3065 23576
rect 3053 23545 3065 23548
rect 3099 23576 3111 23579
rect 3142 23576 3148 23588
rect 3099 23548 3148 23576
rect 3099 23545 3111 23548
rect 3053 23539 3111 23545
rect 3142 23536 3148 23548
rect 3200 23536 3206 23588
rect 3326 23468 3332 23520
rect 3384 23508 3390 23520
rect 3436 23517 3464 23616
rect 3605 23613 3617 23616
rect 3651 23613 3663 23647
rect 3605 23607 3663 23613
rect 4157 23647 4215 23653
rect 4157 23613 4169 23647
rect 4203 23644 4215 23647
rect 4246 23644 4252 23656
rect 4203 23616 4252 23644
rect 4203 23613 4215 23616
rect 4157 23607 4215 23613
rect 4246 23604 4252 23616
rect 4304 23604 4310 23656
rect 5074 23644 5080 23656
rect 4987 23616 5080 23644
rect 5074 23604 5080 23616
rect 5132 23644 5138 23656
rect 5442 23644 5448 23656
rect 5132 23616 5448 23644
rect 5132 23604 5138 23616
rect 5442 23604 5448 23616
rect 5500 23604 5506 23656
rect 5534 23604 5540 23656
rect 5592 23644 5598 23656
rect 5629 23647 5687 23653
rect 5629 23644 5641 23647
rect 5592 23616 5641 23644
rect 5592 23604 5598 23616
rect 5629 23613 5641 23616
rect 5675 23613 5687 23647
rect 6270 23644 6276 23656
rect 6231 23616 6276 23644
rect 5629 23607 5687 23613
rect 6270 23604 6276 23616
rect 6328 23604 6334 23656
rect 6822 23644 6828 23656
rect 6783 23616 6828 23644
rect 6822 23604 6828 23616
rect 6880 23604 6886 23656
rect 9861 23647 9919 23653
rect 9861 23613 9873 23647
rect 9907 23644 9919 23647
rect 10137 23647 10195 23653
rect 10137 23644 10149 23647
rect 9907 23616 10149 23644
rect 9907 23613 9919 23616
rect 9861 23607 9919 23613
rect 10137 23613 10149 23616
rect 10183 23613 10195 23647
rect 10137 23607 10195 23613
rect 10226 23604 10232 23656
rect 10284 23644 10290 23656
rect 10428 23644 10456 23672
rect 10597 23647 10655 23653
rect 10597 23644 10609 23647
rect 10284 23616 10609 23644
rect 10284 23604 10290 23616
rect 10597 23613 10609 23616
rect 10643 23613 10655 23647
rect 12618 23644 12624 23656
rect 12579 23616 12624 23644
rect 10597 23607 10655 23613
rect 12618 23604 12624 23616
rect 12676 23604 12682 23656
rect 5902 23576 5908 23588
rect 5863 23548 5908 23576
rect 5902 23536 5908 23548
rect 5960 23536 5966 23588
rect 6638 23536 6644 23588
rect 6696 23576 6702 23588
rect 7146 23579 7204 23585
rect 7146 23576 7158 23579
rect 6696 23548 7158 23576
rect 6696 23536 6702 23548
rect 7146 23545 7158 23548
rect 7192 23545 7204 23579
rect 8662 23576 8668 23588
rect 7146 23539 7204 23545
rect 8036 23548 8524 23576
rect 8623 23548 8668 23576
rect 3421 23511 3479 23517
rect 3421 23508 3433 23511
rect 3384 23480 3433 23508
rect 3384 23468 3390 23480
rect 3421 23477 3433 23480
rect 3467 23477 3479 23511
rect 3421 23471 3479 23477
rect 3881 23511 3939 23517
rect 3881 23477 3893 23511
rect 3927 23508 3939 23511
rect 4062 23508 4068 23520
rect 3927 23480 4068 23508
rect 3927 23477 3939 23480
rect 3881 23471 3939 23477
rect 4062 23468 4068 23480
rect 4120 23468 4126 23520
rect 4706 23508 4712 23520
rect 4619 23480 4712 23508
rect 4706 23468 4712 23480
rect 4764 23508 4770 23520
rect 5258 23508 5264 23520
rect 4764 23480 5264 23508
rect 4764 23468 4770 23480
rect 5258 23468 5264 23480
rect 5316 23468 5322 23520
rect 8036 23517 8064 23548
rect 7745 23511 7803 23517
rect 7745 23477 7757 23511
rect 7791 23508 7803 23511
rect 8021 23511 8079 23517
rect 8021 23508 8033 23511
rect 7791 23480 8033 23508
rect 7791 23477 7803 23480
rect 7745 23471 7803 23477
rect 8021 23477 8033 23480
rect 8067 23477 8079 23511
rect 8386 23508 8392 23520
rect 8347 23480 8392 23508
rect 8021 23471 8079 23477
rect 8386 23468 8392 23480
rect 8444 23468 8450 23520
rect 8496 23508 8524 23548
rect 8662 23536 8668 23548
rect 8720 23536 8726 23588
rect 8757 23579 8815 23585
rect 8757 23545 8769 23579
rect 8803 23545 8815 23579
rect 9674 23576 9680 23588
rect 9587 23548 9680 23576
rect 8757 23539 8815 23545
rect 8772 23508 8800 23539
rect 9674 23536 9680 23548
rect 9732 23576 9738 23588
rect 10410 23576 10416 23588
rect 9732 23548 10416 23576
rect 9732 23536 9738 23548
rect 10410 23536 10416 23548
rect 10468 23536 10474 23588
rect 11606 23536 11612 23588
rect 11664 23536 11670 23588
rect 9858 23508 9864 23520
rect 8496 23480 8800 23508
rect 9771 23480 9864 23508
rect 9858 23468 9864 23480
rect 9916 23508 9922 23520
rect 10045 23511 10103 23517
rect 10045 23508 10057 23511
rect 9916 23480 10057 23508
rect 9916 23468 9922 23480
rect 10045 23477 10057 23480
rect 10091 23508 10103 23511
rect 10502 23508 10508 23520
rect 10091 23480 10508 23508
rect 10091 23477 10103 23480
rect 10045 23471 10103 23477
rect 10502 23468 10508 23480
rect 10560 23508 10566 23520
rect 10778 23508 10784 23520
rect 10560 23480 10784 23508
rect 10560 23468 10566 23480
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 11624 23508 11652 23536
rect 12158 23508 12164 23520
rect 11624 23480 12164 23508
rect 12158 23468 12164 23480
rect 12216 23468 12222 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 5902 23264 5908 23316
rect 5960 23304 5966 23316
rect 6181 23307 6239 23313
rect 6181 23304 6193 23307
rect 5960 23276 6193 23304
rect 5960 23264 5966 23276
rect 6181 23273 6193 23276
rect 6227 23273 6239 23307
rect 7282 23304 7288 23316
rect 7243 23276 7288 23304
rect 6181 23267 6239 23273
rect 4982 23236 4988 23248
rect 4943 23208 4988 23236
rect 4982 23196 4988 23208
rect 5040 23196 5046 23248
rect 2958 23168 2964 23180
rect 2919 23140 2964 23168
rect 2958 23128 2964 23140
rect 3016 23128 3022 23180
rect 6196 23168 6224 23267
rect 7282 23264 7288 23276
rect 7340 23264 7346 23316
rect 7926 23304 7932 23316
rect 7887 23276 7932 23304
rect 7926 23264 7932 23276
rect 7984 23264 7990 23316
rect 8938 23304 8944 23316
rect 8899 23276 8944 23304
rect 8938 23264 8944 23276
rect 8996 23264 9002 23316
rect 9861 23307 9919 23313
rect 9861 23273 9873 23307
rect 9907 23304 9919 23307
rect 10226 23304 10232 23316
rect 9907 23276 10232 23304
rect 9907 23273 9919 23276
rect 9861 23267 9919 23273
rect 10226 23264 10232 23276
rect 10284 23264 10290 23316
rect 11422 23304 11428 23316
rect 11164 23276 11428 23304
rect 6638 23196 6644 23248
rect 6696 23245 6702 23248
rect 11164 23245 11192 23276
rect 11422 23264 11428 23276
rect 11480 23304 11486 23316
rect 12621 23307 12679 23313
rect 12621 23304 12633 23307
rect 11480 23276 12633 23304
rect 11480 23264 11486 23276
rect 12621 23273 12633 23276
rect 12667 23273 12679 23307
rect 12621 23267 12679 23273
rect 6696 23239 6744 23245
rect 6696 23205 6698 23239
rect 6732 23205 6744 23239
rect 6696 23199 6744 23205
rect 11149 23239 11207 23245
rect 11149 23205 11161 23239
rect 11195 23205 11207 23239
rect 11149 23199 11207 23205
rect 6696 23196 6702 23199
rect 11238 23196 11244 23248
rect 11296 23236 11302 23248
rect 11296 23208 11341 23236
rect 11296 23196 11302 23208
rect 6365 23171 6423 23177
rect 6365 23168 6377 23171
rect 6196 23140 6377 23168
rect 6365 23137 6377 23140
rect 6411 23137 6423 23171
rect 6365 23131 6423 23137
rect 7006 23128 7012 23180
rect 7064 23168 7070 23180
rect 8110 23168 8116 23180
rect 7064 23140 8116 23168
rect 7064 23128 7070 23140
rect 8110 23128 8116 23140
rect 8168 23128 8174 23180
rect 9674 23168 9680 23180
rect 9635 23140 9680 23168
rect 9674 23128 9680 23140
rect 9732 23168 9738 23180
rect 10137 23171 10195 23177
rect 10137 23168 10149 23171
rect 9732 23140 10149 23168
rect 9732 23128 9738 23140
rect 10137 23137 10149 23140
rect 10183 23137 10195 23171
rect 10137 23131 10195 23137
rect 3510 23060 3516 23112
rect 3568 23100 3574 23112
rect 4893 23103 4951 23109
rect 4893 23100 4905 23103
rect 3568 23072 4905 23100
rect 3568 23060 3574 23072
rect 4893 23069 4905 23072
rect 4939 23100 4951 23103
rect 5626 23100 5632 23112
rect 4939 23072 5632 23100
rect 4939 23069 4951 23072
rect 4893 23063 4951 23069
rect 5626 23060 5632 23072
rect 5684 23060 5690 23112
rect 11514 23100 11520 23112
rect 11475 23072 11520 23100
rect 11514 23060 11520 23072
rect 11572 23060 11578 23112
rect 5442 23032 5448 23044
rect 5403 23004 5448 23032
rect 5442 22992 5448 23004
rect 5500 22992 5506 23044
rect 3145 22967 3203 22973
rect 3145 22933 3157 22967
rect 3191 22964 3203 22967
rect 3326 22964 3332 22976
rect 3191 22936 3332 22964
rect 3191 22933 3203 22936
rect 3145 22927 3203 22933
rect 3326 22924 3332 22936
rect 3384 22924 3390 22976
rect 3697 22967 3755 22973
rect 3697 22933 3709 22967
rect 3743 22964 3755 22967
rect 4246 22964 4252 22976
rect 3743 22936 4252 22964
rect 3743 22933 3755 22936
rect 3697 22927 3755 22933
rect 4246 22924 4252 22936
rect 4304 22924 4310 22976
rect 4614 22964 4620 22976
rect 4575 22936 4620 22964
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 7374 22924 7380 22976
rect 7432 22964 7438 22976
rect 7561 22967 7619 22973
rect 7561 22964 7573 22967
rect 7432 22936 7573 22964
rect 7432 22924 7438 22936
rect 7561 22933 7573 22936
rect 7607 22933 7619 22967
rect 7561 22927 7619 22933
rect 8297 22967 8355 22973
rect 8297 22933 8309 22967
rect 8343 22964 8355 22967
rect 8478 22964 8484 22976
rect 8343 22936 8484 22964
rect 8343 22933 8355 22936
rect 8297 22927 8355 22933
rect 8478 22924 8484 22936
rect 8536 22964 8542 22976
rect 8573 22967 8631 22973
rect 8573 22964 8585 22967
rect 8536 22936 8585 22964
rect 8536 22924 8542 22936
rect 8573 22933 8585 22936
rect 8619 22933 8631 22967
rect 8573 22927 8631 22933
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 2958 22760 2964 22772
rect 2919 22732 2964 22760
rect 2958 22720 2964 22732
rect 3016 22720 3022 22772
rect 3510 22760 3516 22772
rect 3471 22732 3516 22760
rect 3510 22720 3516 22732
rect 3568 22720 3574 22772
rect 4982 22720 4988 22772
rect 5040 22760 5046 22772
rect 5442 22760 5448 22772
rect 5040 22732 5448 22760
rect 5040 22720 5046 22732
rect 5442 22720 5448 22732
rect 5500 22760 5506 22772
rect 5813 22763 5871 22769
rect 5813 22760 5825 22763
rect 5500 22732 5825 22760
rect 5500 22720 5506 22732
rect 5813 22729 5825 22732
rect 5859 22729 5871 22763
rect 5813 22723 5871 22729
rect 6457 22763 6515 22769
rect 6457 22729 6469 22763
rect 6503 22760 6515 22763
rect 6638 22760 6644 22772
rect 6503 22732 6644 22760
rect 6503 22729 6515 22732
rect 6457 22723 6515 22729
rect 3789 22695 3847 22701
rect 3789 22661 3801 22695
rect 3835 22692 3847 22695
rect 4430 22692 4436 22704
rect 3835 22664 4436 22692
rect 3835 22661 3847 22664
rect 3789 22655 3847 22661
rect 4430 22652 4436 22664
rect 4488 22652 4494 22704
rect 4614 22624 4620 22636
rect 4575 22596 4620 22624
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 4982 22584 4988 22636
rect 5040 22624 5046 22636
rect 6472 22624 6500 22723
rect 6638 22720 6644 22732
rect 6696 22720 6702 22772
rect 8110 22760 8116 22772
rect 8071 22732 8116 22760
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 11422 22760 11428 22772
rect 11383 22732 11428 22760
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 12526 22720 12532 22772
rect 12584 22760 12590 22772
rect 12621 22763 12679 22769
rect 12621 22760 12633 22763
rect 12584 22732 12633 22760
rect 12584 22720 12590 22732
rect 12621 22729 12633 22732
rect 12667 22729 12679 22763
rect 12621 22723 12679 22729
rect 10594 22652 10600 22704
rect 10652 22692 10658 22704
rect 13633 22695 13691 22701
rect 13633 22692 13645 22695
rect 10652 22664 13645 22692
rect 10652 22652 10658 22664
rect 13633 22661 13645 22664
rect 13679 22661 13691 22695
rect 13633 22655 13691 22661
rect 7190 22624 7196 22636
rect 5040 22596 6500 22624
rect 7151 22596 7196 22624
rect 5040 22584 5046 22596
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 9858 22624 9864 22636
rect 9771 22596 9864 22624
rect 9858 22584 9864 22596
rect 9916 22624 9922 22636
rect 10045 22627 10103 22633
rect 10045 22624 10057 22627
rect 9916 22596 10057 22624
rect 9916 22584 9922 22596
rect 10045 22593 10057 22596
rect 10091 22593 10103 22627
rect 10410 22624 10416 22636
rect 10371 22596 10416 22624
rect 10045 22587 10103 22593
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 3605 22559 3663 22565
rect 3605 22525 3617 22559
rect 3651 22556 3663 22559
rect 4065 22559 4123 22565
rect 4065 22556 4077 22559
rect 3651 22528 4077 22556
rect 3651 22525 3663 22528
rect 3605 22519 3663 22525
rect 4065 22525 4077 22528
rect 4111 22556 4123 22559
rect 4338 22556 4344 22568
rect 4111 22528 4344 22556
rect 4111 22525 4123 22528
rect 4065 22519 4123 22525
rect 4338 22516 4344 22528
rect 4396 22516 4402 22568
rect 5537 22559 5595 22565
rect 5537 22525 5549 22559
rect 5583 22556 5595 22559
rect 8478 22556 8484 22568
rect 5583 22528 6776 22556
rect 8439 22528 8484 22556
rect 5583 22525 5595 22528
rect 5537 22519 5595 22525
rect 4982 22497 4988 22500
rect 4525 22491 4583 22497
rect 4525 22457 4537 22491
rect 4571 22488 4583 22491
rect 4979 22488 4988 22497
rect 4571 22460 4988 22488
rect 4571 22457 4583 22460
rect 4525 22451 4583 22457
rect 4979 22451 4988 22460
rect 4982 22448 4988 22451
rect 5040 22448 5046 22500
rect 6748 22420 6776 22528
rect 8478 22516 8484 22528
rect 8536 22516 8542 22568
rect 8846 22556 8852 22568
rect 8807 22528 8852 22556
rect 8846 22516 8852 22528
rect 8904 22516 8910 22568
rect 9493 22559 9551 22565
rect 9493 22525 9505 22559
rect 9539 22556 9551 22559
rect 9674 22556 9680 22568
rect 9539 22528 9680 22556
rect 9539 22525 9551 22528
rect 9493 22519 9551 22525
rect 9674 22516 9680 22528
rect 9732 22556 9738 22568
rect 9953 22559 10011 22565
rect 9953 22556 9965 22559
rect 9732 22528 9965 22556
rect 9732 22516 9738 22528
rect 9953 22525 9965 22528
rect 9999 22525 10011 22559
rect 10226 22556 10232 22568
rect 10187 22528 10232 22556
rect 9953 22519 10011 22525
rect 10226 22516 10232 22528
rect 10284 22516 10290 22568
rect 12437 22559 12495 22565
rect 12437 22525 12449 22559
rect 12483 22556 12495 22559
rect 12526 22556 12532 22568
rect 12483 22528 12532 22556
rect 12483 22525 12495 22528
rect 12437 22519 12495 22525
rect 12526 22516 12532 22528
rect 12584 22556 12590 22568
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12584 22528 12909 22556
rect 12584 22516 12590 22528
rect 12897 22525 12909 22528
rect 12943 22525 12955 22559
rect 13446 22556 13452 22568
rect 13407 22528 13452 22556
rect 12897 22519 12955 22525
rect 13446 22516 13452 22528
rect 13504 22556 13510 22568
rect 13909 22559 13967 22565
rect 13909 22556 13921 22559
rect 13504 22528 13921 22556
rect 13504 22516 13510 22528
rect 13909 22525 13921 22528
rect 13955 22525 13967 22559
rect 13909 22519 13967 22525
rect 6914 22488 6920 22500
rect 6875 22460 6920 22488
rect 6914 22448 6920 22460
rect 6972 22448 6978 22500
rect 7009 22491 7067 22497
rect 7009 22457 7021 22491
rect 7055 22488 7067 22491
rect 7374 22488 7380 22500
rect 7055 22460 7380 22488
rect 7055 22457 7067 22460
rect 7009 22451 7067 22457
rect 7024 22420 7052 22451
rect 7374 22448 7380 22460
rect 7432 22448 7438 22500
rect 9122 22488 9128 22500
rect 9083 22460 9128 22488
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 10962 22420 10968 22432
rect 6748 22392 7052 22420
rect 10923 22392 10968 22420
rect 10962 22380 10968 22392
rect 11020 22380 11026 22432
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 11238 22420 11244 22432
rect 11112 22392 11244 22420
rect 11112 22380 11118 22392
rect 11238 22380 11244 22392
rect 11296 22420 11302 22432
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 11296 22392 11713 22420
rect 11296 22380 11302 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 11701 22383 11759 22389
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 5442 22216 5448 22228
rect 5403 22188 5448 22216
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 6549 22219 6607 22225
rect 6549 22185 6561 22219
rect 6595 22216 6607 22219
rect 6822 22216 6828 22228
rect 6595 22188 6828 22216
rect 6595 22185 6607 22188
rect 6549 22179 6607 22185
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 7653 22219 7711 22225
rect 7653 22216 7665 22219
rect 6972 22188 7665 22216
rect 6972 22176 6978 22188
rect 7653 22185 7665 22188
rect 7699 22185 7711 22219
rect 7653 22179 7711 22185
rect 9122 22176 9128 22228
rect 9180 22216 9186 22228
rect 9401 22219 9459 22225
rect 9401 22216 9413 22219
rect 9180 22188 9413 22216
rect 9180 22176 9186 22188
rect 9401 22185 9413 22188
rect 9447 22185 9459 22219
rect 9401 22179 9459 22185
rect 4887 22151 4945 22157
rect 4887 22117 4899 22151
rect 4933 22148 4945 22151
rect 4982 22148 4988 22160
rect 4933 22120 4988 22148
rect 4933 22117 4945 22120
rect 4887 22111 4945 22117
rect 4982 22108 4988 22120
rect 5040 22108 5046 22160
rect 5994 22040 6000 22092
rect 6052 22080 6058 22092
rect 6273 22083 6331 22089
rect 6273 22080 6285 22083
rect 6052 22052 6285 22080
rect 6052 22040 6058 22052
rect 6273 22049 6285 22052
rect 6319 22049 6331 22083
rect 6822 22080 6828 22092
rect 6783 22052 6828 22080
rect 6273 22043 6331 22049
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 8665 22083 8723 22089
rect 8665 22049 8677 22083
rect 8711 22080 8723 22083
rect 9416 22080 9444 22179
rect 10042 22176 10048 22228
rect 10100 22176 10106 22228
rect 10226 22176 10232 22228
rect 10284 22216 10290 22228
rect 10962 22216 10968 22228
rect 10284 22188 10968 22216
rect 10284 22176 10290 22188
rect 10962 22176 10968 22188
rect 11020 22216 11026 22228
rect 12066 22216 12072 22228
rect 11020 22188 12072 22216
rect 11020 22176 11026 22188
rect 12066 22176 12072 22188
rect 12124 22176 12130 22228
rect 10060 22148 10088 22176
rect 10366 22151 10424 22157
rect 10366 22148 10378 22151
rect 10060 22120 10378 22148
rect 10366 22117 10378 22120
rect 10412 22148 10424 22151
rect 12526 22148 12532 22160
rect 10412 22120 11192 22148
rect 12487 22120 12532 22148
rect 10412 22117 10424 22120
rect 10366 22111 10424 22117
rect 10045 22083 10103 22089
rect 10045 22080 10057 22083
rect 8711 22052 9352 22080
rect 9416 22052 10057 22080
rect 8711 22049 8723 22052
rect 8665 22043 8723 22049
rect 4522 22012 4528 22024
rect 4483 21984 4528 22012
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 5534 21972 5540 22024
rect 5592 22012 5598 22024
rect 6840 22012 6868 22040
rect 5592 21984 6868 22012
rect 5592 21972 5598 21984
rect 6914 21972 6920 22024
rect 6972 22012 6978 22024
rect 7377 22015 7435 22021
rect 7377 22012 7389 22015
rect 6972 21984 7389 22012
rect 6972 21972 6978 21984
rect 7377 21981 7389 21984
rect 7423 22012 7435 22015
rect 8754 22012 8760 22024
rect 7423 21984 8760 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 8754 21972 8760 21984
rect 8812 21972 8818 22024
rect 9324 22012 9352 22052
rect 10045 22049 10057 22052
rect 10091 22049 10103 22083
rect 10045 22043 10103 22049
rect 11164 22024 11192 22120
rect 12526 22108 12532 22120
rect 12584 22108 12590 22160
rect 11422 22040 11428 22092
rect 11480 22080 11486 22092
rect 11793 22083 11851 22089
rect 11793 22080 11805 22083
rect 11480 22052 11805 22080
rect 11480 22040 11486 22052
rect 11793 22049 11805 22052
rect 11839 22049 11851 22083
rect 12066 22080 12072 22092
rect 12027 22052 12072 22080
rect 11793 22043 11851 22049
rect 12066 22040 12072 22052
rect 12124 22040 12130 22092
rect 9490 22012 9496 22024
rect 9324 21984 9496 22012
rect 9490 21972 9496 21984
rect 9548 21972 9554 22024
rect 11146 21972 11152 22024
rect 11204 21972 11210 22024
rect 10962 21944 10968 21956
rect 10923 21916 10968 21944
rect 10962 21904 10968 21916
rect 11020 21904 11026 21956
rect 11882 21944 11888 21956
rect 11843 21916 11888 21944
rect 11882 21904 11888 21916
rect 11940 21904 11946 21956
rect 4246 21836 4252 21888
rect 4304 21876 4310 21888
rect 4341 21879 4399 21885
rect 4341 21876 4353 21879
rect 4304 21848 4353 21876
rect 4304 21836 4310 21848
rect 4341 21845 4353 21848
rect 4387 21876 4399 21879
rect 4614 21876 4620 21888
rect 4387 21848 4620 21876
rect 4387 21845 4399 21848
rect 4341 21839 4399 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 9674 21836 9680 21888
rect 9732 21876 9738 21888
rect 9861 21879 9919 21885
rect 9861 21876 9873 21879
rect 9732 21848 9873 21876
rect 9732 21836 9738 21848
rect 9861 21845 9873 21848
rect 9907 21845 9919 21879
rect 9861 21839 9919 21845
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 4982 21632 4988 21684
rect 5040 21672 5046 21684
rect 5261 21675 5319 21681
rect 5261 21672 5273 21675
rect 5040 21644 5273 21672
rect 5040 21632 5046 21644
rect 5261 21641 5273 21644
rect 5307 21672 5319 21675
rect 5442 21672 5448 21684
rect 5307 21644 5448 21672
rect 5307 21641 5319 21644
rect 5261 21635 5319 21641
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 9490 21672 9496 21684
rect 8496 21644 9496 21672
rect 6914 21604 6920 21616
rect 6875 21576 6920 21604
rect 6914 21564 6920 21576
rect 6972 21564 6978 21616
rect 8496 21613 8524 21644
rect 9490 21632 9496 21644
rect 9548 21632 9554 21684
rect 11057 21675 11115 21681
rect 11057 21641 11069 21675
rect 11103 21672 11115 21675
rect 11146 21672 11152 21684
rect 11103 21644 11152 21672
rect 11103 21641 11115 21644
rect 11057 21635 11115 21641
rect 11146 21632 11152 21644
rect 11204 21632 11210 21684
rect 8481 21607 8539 21613
rect 8481 21573 8493 21607
rect 8527 21573 8539 21607
rect 8481 21567 8539 21573
rect 8754 21564 8760 21616
rect 8812 21604 8818 21616
rect 10045 21607 10103 21613
rect 10045 21604 10057 21607
rect 8812 21576 10057 21604
rect 8812 21564 8818 21576
rect 10045 21573 10057 21576
rect 10091 21604 10103 21607
rect 11333 21607 11391 21613
rect 11333 21604 11345 21607
rect 10091 21576 11345 21604
rect 10091 21573 10103 21576
rect 10045 21567 10103 21573
rect 11333 21573 11345 21576
rect 11379 21573 11391 21607
rect 12618 21604 12624 21616
rect 12579 21576 12624 21604
rect 11333 21567 11391 21573
rect 12618 21564 12624 21576
rect 12676 21564 12682 21616
rect 4798 21536 4804 21548
rect 4759 21508 4804 21536
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 7558 21536 7564 21548
rect 7519 21508 7564 21536
rect 7558 21496 7564 21508
rect 7616 21496 7622 21548
rect 9125 21539 9183 21545
rect 9125 21505 9137 21539
rect 9171 21536 9183 21539
rect 9582 21536 9588 21548
rect 9171 21508 9588 21536
rect 9171 21505 9183 21508
rect 9125 21499 9183 21505
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 4341 21471 4399 21477
rect 4341 21437 4353 21471
rect 4387 21437 4399 21471
rect 4341 21431 4399 21437
rect 4356 21400 4384 21431
rect 4614 21428 4620 21480
rect 4672 21468 4678 21480
rect 4709 21471 4767 21477
rect 4709 21468 4721 21471
rect 4672 21440 4721 21468
rect 4672 21428 4678 21440
rect 4709 21437 4721 21440
rect 4755 21437 4767 21471
rect 4709 21431 4767 21437
rect 6641 21471 6699 21477
rect 6641 21437 6653 21471
rect 6687 21468 6699 21471
rect 6730 21468 6736 21480
rect 6687 21440 6736 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 6730 21428 6736 21440
rect 6788 21468 6794 21480
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6788 21440 6837 21468
rect 6788 21428 6794 21440
rect 6825 21437 6837 21440
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 7101 21471 7159 21477
rect 7101 21437 7113 21471
rect 7147 21437 7159 21471
rect 7101 21431 7159 21437
rect 5074 21400 5080 21412
rect 4356 21372 5080 21400
rect 4356 21344 4384 21372
rect 5074 21360 5080 21372
rect 5132 21360 5138 21412
rect 6273 21403 6331 21409
rect 6273 21369 6285 21403
rect 6319 21400 6331 21403
rect 7116 21400 7144 21431
rect 8294 21428 8300 21480
rect 8352 21468 8358 21480
rect 8389 21471 8447 21477
rect 8389 21468 8401 21471
rect 8352 21440 8401 21468
rect 8352 21428 8358 21440
rect 8389 21437 8401 21440
rect 8435 21437 8447 21471
rect 8389 21431 8447 21437
rect 8665 21471 8723 21477
rect 8665 21437 8677 21471
rect 8711 21437 8723 21471
rect 8665 21431 8723 21437
rect 7929 21403 7987 21409
rect 7929 21400 7941 21403
rect 6319 21372 7941 21400
rect 6319 21369 6331 21372
rect 6273 21363 6331 21369
rect 7929 21369 7941 21372
rect 7975 21400 7987 21403
rect 8680 21400 8708 21431
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 9953 21471 10011 21477
rect 9953 21468 9965 21471
rect 9732 21440 9965 21468
rect 9732 21428 9738 21440
rect 9953 21437 9965 21440
rect 9999 21437 10011 21471
rect 9953 21431 10011 21437
rect 10229 21471 10287 21477
rect 10229 21437 10241 21471
rect 10275 21437 10287 21471
rect 10229 21431 10287 21437
rect 10689 21471 10747 21477
rect 10689 21437 10701 21471
rect 10735 21468 10747 21471
rect 12437 21471 12495 21477
rect 12437 21468 12449 21471
rect 10735 21440 12449 21468
rect 10735 21437 10747 21440
rect 10689 21431 10747 21437
rect 12437 21437 12449 21440
rect 12483 21468 12495 21471
rect 12897 21471 12955 21477
rect 12897 21468 12909 21471
rect 12483 21440 12909 21468
rect 12483 21437 12495 21440
rect 12437 21431 12495 21437
rect 12897 21437 12909 21440
rect 12943 21437 12955 21471
rect 12897 21431 12955 21437
rect 7975 21372 9812 21400
rect 7975 21369 7987 21372
rect 7929 21363 7987 21369
rect 9784 21344 9812 21372
rect 3786 21332 3792 21344
rect 3747 21304 3792 21332
rect 3786 21292 3792 21304
rect 3844 21292 3850 21344
rect 4157 21335 4215 21341
rect 4157 21301 4169 21335
rect 4203 21332 4215 21335
rect 4338 21332 4344 21344
rect 4203 21304 4344 21332
rect 4203 21301 4215 21304
rect 4157 21295 4215 21301
rect 4338 21292 4344 21304
rect 4396 21292 4402 21344
rect 4430 21292 4436 21344
rect 4488 21332 4494 21344
rect 5813 21335 5871 21341
rect 5813 21332 5825 21335
rect 4488 21304 5825 21332
rect 4488 21292 4494 21304
rect 5813 21301 5825 21304
rect 5859 21332 5871 21335
rect 5994 21332 6000 21344
rect 5859 21304 6000 21332
rect 5859 21301 5871 21304
rect 5813 21295 5871 21301
rect 5994 21292 6000 21304
rect 6052 21292 6058 21344
rect 8294 21332 8300 21344
rect 8255 21304 8300 21332
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 9766 21332 9772 21344
rect 9727 21304 9772 21332
rect 9766 21292 9772 21304
rect 9824 21332 9830 21344
rect 10244 21332 10272 21431
rect 11514 21360 11520 21412
rect 11572 21400 11578 21412
rect 11882 21400 11888 21412
rect 11572 21372 11888 21400
rect 11572 21360 11578 21372
rect 11882 21360 11888 21372
rect 11940 21400 11946 21412
rect 12161 21403 12219 21409
rect 12161 21400 12173 21403
rect 11940 21372 12173 21400
rect 11940 21360 11946 21372
rect 12161 21369 12173 21372
rect 12207 21369 12219 21403
rect 12161 21363 12219 21369
rect 9824 21304 10272 21332
rect 9824 21292 9830 21304
rect 11422 21292 11428 21344
rect 11480 21332 11486 21344
rect 11793 21335 11851 21341
rect 11793 21332 11805 21335
rect 11480 21304 11805 21332
rect 11480 21292 11486 21304
rect 11793 21301 11805 21304
rect 11839 21301 11851 21335
rect 11793 21295 11851 21301
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 3786 21088 3792 21140
rect 3844 21128 3850 21140
rect 4249 21131 4307 21137
rect 4249 21128 4261 21131
rect 3844 21100 4261 21128
rect 3844 21088 3850 21100
rect 4249 21097 4261 21100
rect 4295 21128 4307 21131
rect 4522 21128 4528 21140
rect 4295 21100 4528 21128
rect 4295 21097 4307 21100
rect 4249 21091 4307 21097
rect 4522 21088 4528 21100
rect 4580 21088 4586 21140
rect 5626 21088 5632 21140
rect 5684 21128 5690 21140
rect 6365 21131 6423 21137
rect 6365 21128 6377 21131
rect 5684 21100 6377 21128
rect 5684 21088 5690 21100
rect 6365 21097 6377 21100
rect 6411 21128 6423 21131
rect 6822 21128 6828 21140
rect 6411 21100 6828 21128
rect 6411 21097 6423 21100
rect 6365 21091 6423 21097
rect 6822 21088 6828 21100
rect 6880 21088 6886 21140
rect 8665 21131 8723 21137
rect 8665 21097 8677 21131
rect 8711 21128 8723 21131
rect 9490 21128 9496 21140
rect 8711 21100 9496 21128
rect 8711 21097 8723 21100
rect 8665 21091 8723 21097
rect 9490 21088 9496 21100
rect 9548 21088 9554 21140
rect 10137 21131 10195 21137
rect 10137 21097 10149 21131
rect 10183 21128 10195 21131
rect 10226 21128 10232 21140
rect 10183 21100 10232 21128
rect 10183 21097 10195 21100
rect 10137 21091 10195 21097
rect 10226 21088 10232 21100
rect 10284 21088 10290 21140
rect 11146 21088 11152 21140
rect 11204 21128 11210 21140
rect 11701 21131 11759 21137
rect 11701 21128 11713 21131
rect 11204 21100 11713 21128
rect 11204 21088 11210 21100
rect 11701 21097 11713 21100
rect 11747 21097 11759 21131
rect 11701 21091 11759 21097
rect 12066 21088 12072 21140
rect 12124 21128 12130 21140
rect 12253 21131 12311 21137
rect 12253 21128 12265 21131
rect 12124 21100 12265 21128
rect 12124 21088 12130 21100
rect 12253 21097 12265 21100
rect 12299 21097 12311 21131
rect 12253 21091 12311 21097
rect 6638 21020 6644 21072
rect 6696 21060 6702 21072
rect 6733 21063 6791 21069
rect 6733 21060 6745 21063
rect 6696 21032 6745 21060
rect 6696 21020 6702 21032
rect 6733 21029 6745 21032
rect 6779 21029 6791 21063
rect 6733 21023 6791 21029
rect 10410 21020 10416 21072
rect 10468 21060 10474 21072
rect 10781 21063 10839 21069
rect 10781 21060 10793 21063
rect 10468 21032 10793 21060
rect 10468 21020 10474 21032
rect 10781 21029 10793 21032
rect 10827 21060 10839 21063
rect 11974 21060 11980 21072
rect 10827 21032 11980 21060
rect 10827 21029 10839 21032
rect 10781 21023 10839 21029
rect 11974 21020 11980 21032
rect 12032 21020 12038 21072
rect 4430 20992 4436 21004
rect 4391 20964 4436 20992
rect 4430 20952 4436 20964
rect 4488 20952 4494 21004
rect 4614 20992 4620 21004
rect 4527 20964 4620 20992
rect 4614 20952 4620 20964
rect 4672 20952 4678 21004
rect 7742 20952 7748 21004
rect 7800 20992 7806 21004
rect 8148 20995 8206 21001
rect 8148 20992 8160 20995
rect 7800 20964 8160 20992
rect 7800 20952 7806 20964
rect 8148 20961 8160 20964
rect 8194 20992 8206 20995
rect 8570 20992 8576 21004
rect 8194 20964 8576 20992
rect 8194 20961 8206 20964
rect 8148 20955 8206 20961
rect 8570 20952 8576 20964
rect 8628 20952 8634 21004
rect 10321 20995 10379 21001
rect 10321 20961 10333 20995
rect 10367 20992 10379 20995
rect 10367 20964 10548 20992
rect 10367 20961 10379 20964
rect 10321 20955 10379 20961
rect 3970 20884 3976 20936
rect 4028 20924 4034 20936
rect 4632 20924 4660 20952
rect 4028 20896 4660 20924
rect 4028 20884 4034 20896
rect 6270 20884 6276 20936
rect 6328 20924 6334 20936
rect 6641 20927 6699 20933
rect 6641 20924 6653 20927
rect 6328 20896 6653 20924
rect 6328 20884 6334 20896
rect 6641 20893 6653 20896
rect 6687 20924 6699 20927
rect 8251 20927 8309 20933
rect 8251 20924 8263 20927
rect 6687 20896 8263 20924
rect 6687 20893 6699 20896
rect 6641 20887 6699 20893
rect 8251 20893 8263 20896
rect 8297 20893 8309 20927
rect 8251 20887 8309 20893
rect 7190 20856 7196 20868
rect 7103 20828 7196 20856
rect 7190 20816 7196 20828
rect 7248 20856 7254 20868
rect 7374 20856 7380 20868
rect 7248 20828 7380 20856
rect 7248 20816 7254 20828
rect 7374 20816 7380 20828
rect 7432 20816 7438 20868
rect 6914 20748 6920 20800
rect 6972 20788 6978 20800
rect 7561 20791 7619 20797
rect 7561 20788 7573 20791
rect 6972 20760 7573 20788
rect 6972 20748 6978 20760
rect 7561 20757 7573 20760
rect 7607 20757 7619 20791
rect 7561 20751 7619 20757
rect 9493 20791 9551 20797
rect 9493 20757 9505 20791
rect 9539 20788 9551 20791
rect 9674 20788 9680 20800
rect 9539 20760 9680 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 9766 20748 9772 20800
rect 9824 20788 9830 20800
rect 10520 20788 10548 20964
rect 11146 20952 11152 21004
rect 11204 20992 11210 21004
rect 11241 20995 11299 21001
rect 11241 20992 11253 20995
rect 11204 20964 11253 20992
rect 11204 20952 11210 20964
rect 11241 20961 11253 20964
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 11517 20995 11575 21001
rect 11517 20961 11529 20995
rect 11563 20992 11575 20995
rect 11606 20992 11612 21004
rect 11563 20964 11612 20992
rect 11563 20961 11575 20964
rect 11517 20955 11575 20961
rect 11606 20952 11612 20964
rect 11664 20952 11670 21004
rect 11333 20859 11391 20865
rect 11333 20825 11345 20859
rect 11379 20856 11391 20859
rect 11514 20856 11520 20868
rect 11379 20828 11520 20856
rect 11379 20825 11391 20828
rect 11333 20819 11391 20825
rect 11514 20816 11520 20828
rect 11572 20856 11578 20868
rect 12066 20856 12072 20868
rect 11572 20828 12072 20856
rect 11572 20816 11578 20828
rect 12066 20816 12072 20828
rect 12124 20816 12130 20868
rect 11606 20788 11612 20800
rect 9824 20760 11612 20788
rect 9824 20748 9830 20760
rect 11606 20748 11612 20760
rect 11664 20748 11670 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 6270 20584 6276 20596
rect 6231 20556 6276 20584
rect 6270 20544 6276 20556
rect 6328 20544 6334 20596
rect 9766 20584 9772 20596
rect 9727 20556 9772 20584
rect 9766 20544 9772 20556
rect 9824 20544 9830 20596
rect 11974 20584 11980 20596
rect 11935 20556 11980 20584
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 5350 20516 5356 20528
rect 5311 20488 5356 20516
rect 5350 20476 5356 20488
rect 5408 20476 5414 20528
rect 10045 20519 10103 20525
rect 10045 20485 10057 20519
rect 10091 20516 10103 20519
rect 10870 20516 10876 20528
rect 10091 20488 10876 20516
rect 10091 20485 10103 20488
rect 10045 20479 10103 20485
rect 10870 20476 10876 20488
rect 10928 20476 10934 20528
rect 7374 20448 7380 20460
rect 7335 20420 7380 20448
rect 7374 20408 7380 20420
rect 7432 20408 7438 20460
rect 3764 20383 3822 20389
rect 3764 20349 3776 20383
rect 3810 20380 3822 20383
rect 8294 20380 8300 20392
rect 3810 20352 4292 20380
rect 8207 20352 8300 20380
rect 3810 20349 3822 20352
rect 3764 20343 3822 20349
rect 3605 20315 3663 20321
rect 3605 20281 3617 20315
rect 3651 20312 3663 20315
rect 3970 20312 3976 20324
rect 3651 20284 3976 20312
rect 3651 20281 3663 20284
rect 3605 20275 3663 20281
rect 3970 20272 3976 20284
rect 4028 20272 4034 20324
rect 4264 20256 4292 20352
rect 8294 20340 8300 20352
rect 8352 20380 8358 20392
rect 8754 20380 8760 20392
rect 8352 20352 8760 20380
rect 8352 20340 8358 20352
rect 8754 20340 8760 20352
rect 8812 20340 8818 20392
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 9953 20383 10011 20389
rect 9953 20380 9965 20383
rect 9732 20352 9965 20380
rect 9732 20340 9738 20352
rect 9953 20349 9965 20352
rect 9999 20349 10011 20383
rect 9953 20343 10011 20349
rect 10229 20383 10287 20389
rect 10229 20349 10241 20383
rect 10275 20380 10287 20383
rect 10410 20380 10416 20392
rect 10275 20352 10416 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 4798 20312 4804 20324
rect 4759 20284 4804 20312
rect 4798 20272 4804 20284
rect 4856 20272 4862 20324
rect 4890 20272 4896 20324
rect 4948 20312 4954 20324
rect 6914 20312 6920 20324
rect 4948 20284 4993 20312
rect 6875 20284 6920 20312
rect 4948 20272 4954 20284
rect 6914 20272 6920 20284
rect 6972 20272 6978 20324
rect 7006 20272 7012 20324
rect 7064 20312 7070 20324
rect 10686 20312 10692 20324
rect 7064 20284 7109 20312
rect 10647 20284 10692 20312
rect 7064 20272 7070 20284
rect 10686 20272 10692 20284
rect 10744 20272 10750 20324
rect 11333 20315 11391 20321
rect 11333 20281 11345 20315
rect 11379 20312 11391 20315
rect 11606 20312 11612 20324
rect 11379 20284 11612 20312
rect 11379 20281 11391 20284
rect 11333 20275 11391 20281
rect 11606 20272 11612 20284
rect 11664 20312 11670 20324
rect 11974 20312 11980 20324
rect 11664 20284 11980 20312
rect 11664 20272 11670 20284
rect 11974 20272 11980 20284
rect 12032 20272 12038 20324
rect 3878 20253 3884 20256
rect 3835 20247 3884 20253
rect 3835 20213 3847 20247
rect 3881 20213 3884 20247
rect 3835 20207 3884 20213
rect 3878 20204 3884 20207
rect 3936 20204 3942 20256
rect 4246 20244 4252 20256
rect 4207 20216 4252 20244
rect 4246 20204 4252 20216
rect 4304 20204 4310 20256
rect 4430 20204 4436 20256
rect 4488 20244 4494 20256
rect 4614 20244 4620 20256
rect 4488 20216 4620 20244
rect 4488 20204 4494 20216
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 6638 20244 6644 20256
rect 6599 20216 6644 20244
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 7742 20204 7748 20256
rect 7800 20244 7806 20256
rect 7837 20247 7895 20253
rect 7837 20244 7849 20247
rect 7800 20216 7849 20244
rect 7800 20204 7806 20216
rect 7837 20213 7849 20216
rect 7883 20213 7895 20247
rect 7837 20207 7895 20213
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 8665 20247 8723 20253
rect 8665 20244 8677 20247
rect 8536 20216 8677 20244
rect 8536 20204 8542 20216
rect 8665 20213 8677 20216
rect 8711 20244 8723 20247
rect 9582 20244 9588 20256
rect 8711 20216 9588 20244
rect 8711 20213 8723 20216
rect 8665 20207 8723 20213
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 11701 20247 11759 20253
rect 11701 20213 11713 20247
rect 11747 20244 11759 20247
rect 12066 20244 12072 20256
rect 11747 20216 12072 20244
rect 11747 20213 11759 20216
rect 11701 20207 11759 20213
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4387 20043 4445 20049
rect 4387 20040 4399 20043
rect 4212 20012 4399 20040
rect 4212 20000 4218 20012
rect 4387 20009 4399 20012
rect 4433 20009 4445 20043
rect 4387 20003 4445 20009
rect 4890 20000 4896 20052
rect 4948 20040 4954 20052
rect 5077 20043 5135 20049
rect 5077 20040 5089 20043
rect 4948 20012 5089 20040
rect 4948 20000 4954 20012
rect 5077 20009 5089 20012
rect 5123 20009 5135 20043
rect 5077 20003 5135 20009
rect 6457 20043 6515 20049
rect 6457 20009 6469 20043
rect 6503 20009 6515 20043
rect 6457 20003 6515 20009
rect 9493 20043 9551 20049
rect 9493 20009 9505 20043
rect 9539 20040 9551 20043
rect 10870 20040 10876 20052
rect 9539 20012 10876 20040
rect 9539 20009 9551 20012
rect 9493 20003 9551 20009
rect 2961 19975 3019 19981
rect 2961 19941 2973 19975
rect 3007 19972 3019 19975
rect 4709 19975 4767 19981
rect 4709 19972 4721 19975
rect 3007 19944 4721 19972
rect 3007 19941 3019 19944
rect 2961 19935 3019 19941
rect 4709 19941 4721 19944
rect 4755 19972 4767 19975
rect 4798 19972 4804 19984
rect 4755 19944 4804 19972
rect 4755 19941 4767 19944
rect 4709 19935 4767 19941
rect 4798 19932 4804 19944
rect 4856 19932 4862 19984
rect 5534 19932 5540 19984
rect 5592 19972 5598 19984
rect 5718 19972 5724 19984
rect 5592 19944 5724 19972
rect 5592 19932 5598 19944
rect 5718 19932 5724 19944
rect 5776 19972 5782 19984
rect 5858 19975 5916 19981
rect 5858 19972 5870 19975
rect 5776 19944 5870 19972
rect 5776 19932 5782 19944
rect 5858 19941 5870 19944
rect 5904 19941 5916 19975
rect 6472 19972 6500 20003
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 6638 19972 6644 19984
rect 6472 19944 6644 19972
rect 5858 19935 5916 19941
rect 6638 19932 6644 19944
rect 6696 19972 6702 19984
rect 7469 19975 7527 19981
rect 7469 19972 7481 19975
rect 6696 19944 7481 19972
rect 6696 19932 6702 19944
rect 7469 19941 7481 19944
rect 7515 19972 7527 19975
rect 7834 19972 7840 19984
rect 7515 19944 7840 19972
rect 7515 19941 7527 19944
rect 7469 19935 7527 19941
rect 7834 19932 7840 19944
rect 7892 19932 7898 19984
rect 4062 19864 4068 19916
rect 4120 19904 4126 19916
rect 4316 19907 4374 19913
rect 4316 19904 4328 19907
rect 4120 19876 4328 19904
rect 4120 19864 4126 19876
rect 4316 19873 4328 19876
rect 4362 19904 4374 19907
rect 5350 19904 5356 19916
rect 4362 19876 5356 19904
rect 4362 19873 4374 19876
rect 4316 19867 4374 19873
rect 5350 19864 5356 19876
rect 5408 19864 5414 19916
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 9861 19907 9919 19913
rect 9861 19904 9873 19907
rect 9732 19876 9873 19904
rect 9732 19864 9738 19876
rect 9861 19873 9873 19876
rect 9907 19904 9919 19907
rect 10042 19904 10048 19916
rect 9907 19876 10048 19904
rect 9907 19873 9919 19876
rect 9861 19867 9919 19873
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19904 10195 19907
rect 10410 19904 10416 19916
rect 10183 19876 10416 19904
rect 10183 19873 10195 19876
rect 10137 19867 10195 19873
rect 10410 19864 10416 19876
rect 10468 19864 10474 19916
rect 10686 19864 10692 19916
rect 10744 19904 10750 19916
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 10744 19876 11437 19904
rect 10744 19864 10750 19876
rect 11425 19873 11437 19876
rect 11471 19904 11483 19907
rect 11514 19904 11520 19916
rect 11471 19876 11520 19904
rect 11471 19873 11483 19876
rect 11425 19867 11483 19873
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 5534 19836 5540 19848
rect 5495 19808 5540 19836
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 7190 19796 7196 19848
rect 7248 19836 7254 19848
rect 7377 19839 7435 19845
rect 7377 19836 7389 19839
rect 7248 19808 7389 19836
rect 7248 19796 7254 19808
rect 7377 19805 7389 19808
rect 7423 19836 7435 19839
rect 8294 19836 8300 19848
rect 7423 19808 8300 19836
rect 7423 19805 7435 19808
rect 7377 19799 7435 19805
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 10318 19836 10324 19848
rect 10279 19808 10324 19836
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 7926 19768 7932 19780
rect 7887 19740 7932 19768
rect 7926 19728 7932 19740
rect 7984 19728 7990 19780
rect 9950 19768 9956 19780
rect 9911 19740 9956 19768
rect 9950 19728 9956 19740
rect 10008 19728 10014 19780
rect 10502 19728 10508 19780
rect 10560 19768 10566 19780
rect 11609 19771 11667 19777
rect 11609 19768 11621 19771
rect 10560 19740 11621 19768
rect 10560 19728 10566 19740
rect 11609 19737 11621 19740
rect 11655 19737 11667 19771
rect 11609 19731 11667 19737
rect 6914 19700 6920 19712
rect 6875 19672 6920 19700
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 8386 19700 8392 19712
rect 8347 19672 8392 19700
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 4890 19456 4896 19508
rect 4948 19496 4954 19508
rect 5169 19499 5227 19505
rect 5169 19496 5181 19499
rect 4948 19468 5181 19496
rect 4948 19456 4954 19468
rect 5169 19465 5181 19468
rect 5215 19465 5227 19499
rect 5169 19459 5227 19465
rect 5629 19499 5687 19505
rect 5629 19465 5641 19499
rect 5675 19496 5687 19499
rect 5718 19496 5724 19508
rect 5675 19468 5724 19496
rect 5675 19465 5687 19468
rect 5629 19459 5687 19465
rect 5718 19456 5724 19468
rect 5776 19456 5782 19508
rect 7834 19496 7840 19508
rect 7795 19468 7840 19496
rect 7834 19456 7840 19468
rect 7892 19456 7898 19508
rect 9677 19499 9735 19505
rect 9677 19465 9689 19499
rect 9723 19496 9735 19499
rect 10410 19496 10416 19508
rect 9723 19468 10416 19496
rect 9723 19465 9735 19468
rect 9677 19459 9735 19465
rect 10410 19456 10416 19468
rect 10468 19456 10474 19508
rect 10870 19496 10876 19508
rect 10831 19468 10876 19496
rect 10870 19456 10876 19468
rect 10928 19456 10934 19508
rect 11514 19496 11520 19508
rect 11475 19468 11520 19496
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 6917 19363 6975 19369
rect 6917 19329 6929 19363
rect 6963 19360 6975 19363
rect 7006 19360 7012 19372
rect 6963 19332 7012 19360
rect 6963 19329 6975 19332
rect 6917 19323 6975 19329
rect 7006 19320 7012 19332
rect 7064 19320 7070 19372
rect 7561 19363 7619 19369
rect 7561 19329 7573 19363
rect 7607 19360 7619 19363
rect 7926 19360 7932 19372
rect 7607 19332 7932 19360
rect 7607 19329 7619 19332
rect 7561 19323 7619 19329
rect 7926 19320 7932 19332
rect 7984 19320 7990 19372
rect 8386 19360 8392 19372
rect 8220 19332 8392 19360
rect 2685 19295 2743 19301
rect 2685 19292 2697 19295
rect 2516 19264 2697 19292
rect 2516 19224 2544 19264
rect 2685 19261 2697 19264
rect 2731 19261 2743 19295
rect 2685 19255 2743 19261
rect 3234 19252 3240 19304
rect 3292 19292 3298 19304
rect 3789 19295 3847 19301
rect 3292 19264 3337 19292
rect 3292 19252 3298 19264
rect 3789 19261 3801 19295
rect 3835 19292 3847 19295
rect 4062 19292 4068 19304
rect 3835 19264 4068 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4249 19295 4307 19301
rect 4249 19292 4261 19295
rect 4212 19264 4261 19292
rect 4212 19252 4218 19264
rect 4249 19261 4261 19264
rect 4295 19261 4307 19295
rect 5534 19292 5540 19304
rect 4249 19255 4307 19261
rect 4448 19264 5540 19292
rect 3050 19224 3056 19236
rect 2516 19196 3056 19224
rect 2406 19116 2412 19168
rect 2464 19156 2470 19168
rect 2516 19165 2544 19196
rect 3050 19184 3056 19196
rect 3108 19184 3114 19236
rect 3421 19227 3479 19233
rect 3421 19193 3433 19227
rect 3467 19224 3479 19227
rect 4448 19224 4476 19264
rect 5534 19252 5540 19264
rect 5592 19292 5598 19304
rect 5905 19295 5963 19301
rect 5905 19292 5917 19295
rect 5592 19264 5917 19292
rect 5592 19252 5598 19264
rect 5905 19261 5917 19264
rect 5951 19261 5963 19295
rect 5905 19255 5963 19261
rect 4611 19227 4669 19233
rect 4611 19224 4623 19227
rect 3467 19196 4476 19224
rect 4540 19196 4623 19224
rect 3467 19193 3479 19196
rect 3421 19187 3479 19193
rect 2501 19159 2559 19165
rect 2501 19156 2513 19159
rect 2464 19128 2513 19156
rect 2464 19116 2470 19128
rect 2501 19125 2513 19128
rect 2547 19125 2559 19159
rect 2501 19119 2559 19125
rect 4157 19159 4215 19165
rect 4157 19125 4169 19159
rect 4203 19156 4215 19159
rect 4540 19156 4568 19196
rect 4611 19193 4623 19196
rect 4657 19224 4669 19227
rect 5718 19224 5724 19236
rect 4657 19196 5724 19224
rect 4657 19193 4669 19196
rect 4611 19187 4669 19193
rect 5718 19184 5724 19196
rect 5776 19184 5782 19236
rect 7009 19227 7067 19233
rect 7009 19193 7021 19227
rect 7055 19193 7067 19227
rect 7009 19187 7067 19193
rect 6638 19156 6644 19168
rect 4203 19128 4568 19156
rect 6551 19128 6644 19156
rect 4203 19125 4215 19128
rect 4157 19119 4215 19125
rect 6638 19116 6644 19128
rect 6696 19156 6702 19168
rect 7024 19156 7052 19187
rect 7098 19184 7104 19236
rect 7156 19224 7162 19236
rect 8220 19224 8248 19332
rect 8386 19320 8392 19332
rect 8444 19320 8450 19372
rect 8938 19360 8944 19372
rect 8899 19332 8944 19360
rect 8938 19320 8944 19332
rect 8996 19320 9002 19372
rect 8573 19295 8631 19301
rect 8573 19261 8585 19295
rect 8619 19292 8631 19295
rect 9214 19292 9220 19304
rect 8619 19264 9220 19292
rect 8619 19261 8631 19264
rect 8573 19255 8631 19261
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 9858 19252 9864 19304
rect 9916 19292 9922 19304
rect 10413 19295 10471 19301
rect 10413 19292 10425 19295
rect 9916 19264 10425 19292
rect 9916 19252 9922 19264
rect 10413 19261 10425 19264
rect 10459 19292 10471 19295
rect 10870 19292 10876 19304
rect 10459 19264 10876 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 10870 19252 10876 19264
rect 10928 19252 10934 19304
rect 7156 19196 8248 19224
rect 8297 19227 8355 19233
rect 7156 19184 7162 19196
rect 8297 19193 8309 19227
rect 8343 19224 8355 19227
rect 8386 19224 8392 19236
rect 8343 19196 8392 19224
rect 8343 19193 8355 19196
rect 8297 19187 8355 19193
rect 8386 19184 8392 19196
rect 8444 19184 8450 19236
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10505 19227 10563 19233
rect 10505 19224 10517 19227
rect 10008 19196 10517 19224
rect 10008 19184 10014 19196
rect 10505 19193 10517 19196
rect 10551 19224 10563 19227
rect 11149 19227 11207 19233
rect 11149 19224 11161 19227
rect 10551 19196 11161 19224
rect 10551 19193 10563 19196
rect 10505 19187 10563 19193
rect 11149 19193 11161 19196
rect 11195 19193 11207 19227
rect 11149 19187 11207 19193
rect 6696 19128 7052 19156
rect 6696 19116 6702 19128
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 2774 18952 2780 18964
rect 2735 18924 2780 18952
rect 2774 18912 2780 18924
rect 2832 18912 2838 18964
rect 3099 18955 3157 18961
rect 3099 18921 3111 18955
rect 3145 18952 3157 18955
rect 3418 18952 3424 18964
rect 3145 18924 3424 18952
rect 3145 18921 3157 18924
rect 3099 18915 3157 18921
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18921 6515 18955
rect 8294 18952 8300 18964
rect 8255 18924 8300 18952
rect 6457 18915 6515 18921
rect 5718 18844 5724 18896
rect 5776 18884 5782 18896
rect 5858 18887 5916 18893
rect 5858 18884 5870 18887
rect 5776 18856 5870 18884
rect 5776 18844 5782 18856
rect 5858 18853 5870 18856
rect 5904 18853 5916 18887
rect 6472 18884 6500 18915
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 9401 18955 9459 18961
rect 9401 18921 9413 18955
rect 9447 18952 9459 18955
rect 9582 18952 9588 18964
rect 9447 18924 9588 18952
rect 9447 18921 9459 18924
rect 9401 18915 9459 18921
rect 9582 18912 9588 18924
rect 9640 18952 9646 18964
rect 9950 18952 9956 18964
rect 9640 18924 9956 18952
rect 9640 18912 9646 18924
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 10594 18952 10600 18964
rect 10100 18924 10600 18952
rect 10100 18912 10106 18924
rect 10594 18912 10600 18924
rect 10652 18952 10658 18964
rect 10689 18955 10747 18961
rect 10689 18952 10701 18955
rect 10652 18924 10701 18952
rect 10652 18912 10658 18924
rect 10689 18921 10701 18924
rect 10735 18921 10747 18955
rect 10689 18915 10747 18921
rect 6914 18884 6920 18896
rect 6472 18856 6920 18884
rect 5858 18847 5916 18853
rect 6914 18844 6920 18856
rect 6972 18884 6978 18896
rect 7469 18887 7527 18893
rect 7469 18884 7481 18887
rect 6972 18856 7481 18884
rect 6972 18844 6978 18856
rect 7469 18853 7481 18856
rect 7515 18884 7527 18887
rect 8018 18884 8024 18896
rect 7515 18856 8024 18884
rect 7515 18853 7527 18856
rect 7469 18847 7527 18853
rect 8018 18844 8024 18856
rect 8076 18844 8082 18896
rect 10410 18884 10416 18896
rect 9968 18856 10416 18884
rect 2038 18825 2044 18828
rect 2016 18819 2044 18825
rect 2016 18785 2028 18819
rect 2016 18779 2044 18785
rect 2038 18776 2044 18779
rect 2096 18776 2102 18828
rect 3028 18819 3086 18825
rect 3028 18785 3040 18819
rect 3074 18816 3086 18819
rect 3142 18816 3148 18828
rect 3074 18788 3148 18816
rect 3074 18785 3086 18788
rect 3028 18779 3086 18785
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 4430 18776 4436 18828
rect 4488 18816 4494 18828
rect 4560 18819 4618 18825
rect 4560 18816 4572 18819
rect 4488 18788 4572 18816
rect 4488 18776 4494 18788
rect 4560 18785 4572 18788
rect 4606 18785 4618 18819
rect 9033 18819 9091 18825
rect 4560 18779 4618 18785
rect 4678 18788 5856 18816
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 3513 18751 3571 18757
rect 3513 18748 3525 18751
rect 3476 18720 3525 18748
rect 3476 18708 3482 18720
rect 3513 18717 3525 18720
rect 3559 18748 3571 18751
rect 4678 18748 4706 18788
rect 3559 18720 4706 18748
rect 5537 18751 5595 18757
rect 3559 18717 3571 18720
rect 3513 18711 3571 18717
rect 5537 18717 5549 18751
rect 5583 18748 5595 18751
rect 5718 18748 5724 18760
rect 5583 18720 5724 18748
rect 5583 18717 5595 18720
rect 5537 18711 5595 18717
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 4663 18683 4721 18689
rect 4663 18649 4675 18683
rect 4709 18680 4721 18683
rect 5626 18680 5632 18692
rect 4709 18652 5632 18680
rect 4709 18649 4721 18652
rect 4663 18643 4721 18649
rect 5626 18640 5632 18652
rect 5684 18640 5690 18692
rect 5828 18680 5856 18788
rect 9033 18785 9045 18819
rect 9079 18816 9091 18819
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 9079 18788 9689 18816
rect 9079 18785 9091 18788
rect 9033 18779 9091 18785
rect 9677 18785 9689 18788
rect 9723 18816 9735 18819
rect 9766 18816 9772 18828
rect 9723 18788 9772 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 9766 18776 9772 18788
rect 9824 18776 9830 18828
rect 9968 18825 9996 18856
rect 10410 18844 10416 18856
rect 10468 18844 10474 18896
rect 9953 18819 10011 18825
rect 9953 18785 9965 18819
rect 9999 18785 10011 18819
rect 9953 18779 10011 18785
rect 11238 18776 11244 18828
rect 11296 18816 11302 18828
rect 11333 18819 11391 18825
rect 11333 18816 11345 18819
rect 11296 18788 11345 18816
rect 11296 18776 11302 18788
rect 11333 18785 11345 18788
rect 11379 18816 11391 18819
rect 13078 18816 13084 18828
rect 11379 18788 13084 18816
rect 11379 18785 11391 18788
rect 11333 18779 11391 18785
rect 13078 18776 13084 18788
rect 13136 18776 13142 18828
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 7377 18751 7435 18757
rect 7377 18748 7389 18751
rect 6236 18720 7389 18748
rect 6236 18708 6242 18720
rect 7377 18717 7389 18720
rect 7423 18717 7435 18751
rect 8570 18748 8576 18760
rect 7377 18711 7435 18717
rect 7484 18720 8576 18748
rect 7484 18680 7512 18720
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 10410 18748 10416 18760
rect 10371 18720 10416 18748
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 7926 18680 7932 18692
rect 5828 18652 7512 18680
rect 7887 18652 7932 18680
rect 7926 18640 7932 18652
rect 7984 18640 7990 18692
rect 9769 18683 9827 18689
rect 9769 18649 9781 18683
rect 9815 18680 9827 18683
rect 9858 18680 9864 18692
rect 9815 18652 9864 18680
rect 9815 18649 9827 18652
rect 9769 18643 9827 18649
rect 9858 18640 9864 18652
rect 9916 18640 9922 18692
rect 11422 18640 11428 18692
rect 11480 18680 11486 18692
rect 12250 18680 12256 18692
rect 11480 18652 12256 18680
rect 11480 18640 11486 18652
rect 12250 18640 12256 18652
rect 12308 18640 12314 18692
rect 2087 18615 2145 18621
rect 2087 18581 2099 18615
rect 2133 18612 2145 18615
rect 3234 18612 3240 18624
rect 2133 18584 3240 18612
rect 2133 18581 2145 18584
rect 2087 18575 2145 18581
rect 3234 18572 3240 18584
rect 3292 18572 3298 18624
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 4249 18615 4307 18621
rect 4249 18612 4261 18615
rect 4212 18584 4261 18612
rect 4212 18572 4218 18584
rect 4249 18581 4261 18584
rect 4295 18581 4307 18615
rect 4249 18575 4307 18581
rect 4890 18572 4896 18624
rect 4948 18612 4954 18624
rect 4985 18615 5043 18621
rect 4985 18612 4997 18615
rect 4948 18584 4997 18612
rect 4948 18572 4954 18584
rect 4985 18581 4997 18584
rect 5031 18612 5043 18615
rect 5258 18612 5264 18624
rect 5031 18584 5264 18612
rect 5031 18581 5043 18584
rect 4985 18575 5043 18581
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 5445 18615 5503 18621
rect 5445 18581 5457 18615
rect 5491 18612 5503 18615
rect 5534 18612 5540 18624
rect 5491 18584 5540 18612
rect 5491 18581 5503 18584
rect 5445 18575 5503 18581
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 6822 18612 6828 18624
rect 6783 18584 6828 18612
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 11517 18615 11575 18621
rect 11517 18612 11529 18615
rect 11204 18584 11529 18612
rect 11204 18572 11210 18584
rect 11517 18581 11529 18584
rect 11563 18581 11575 18615
rect 11517 18575 11575 18581
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 2593 18411 2651 18417
rect 2593 18377 2605 18411
rect 2639 18408 2651 18411
rect 2774 18408 2780 18420
rect 2639 18380 2780 18408
rect 2639 18377 2651 18380
rect 2593 18371 2651 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 3053 18411 3111 18417
rect 3053 18377 3065 18411
rect 3099 18408 3111 18411
rect 3142 18408 3148 18420
rect 3099 18380 3148 18408
rect 3099 18377 3111 18380
rect 3053 18371 3111 18377
rect 3142 18368 3148 18380
rect 3200 18368 3206 18420
rect 5258 18368 5264 18420
rect 5316 18408 5322 18420
rect 5810 18408 5816 18420
rect 5316 18380 5816 18408
rect 5316 18368 5322 18380
rect 5810 18368 5816 18380
rect 5868 18408 5874 18420
rect 5997 18411 6055 18417
rect 5997 18408 6009 18411
rect 5868 18380 6009 18408
rect 5868 18368 5874 18380
rect 5997 18377 6009 18380
rect 6043 18408 6055 18411
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6043 18380 6561 18408
rect 6043 18377 6055 18380
rect 5997 18371 6055 18377
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 8018 18408 8024 18420
rect 7979 18380 8024 18408
rect 6549 18371 6607 18377
rect 4154 18272 4160 18284
rect 4115 18244 4160 18272
rect 4154 18232 4160 18244
rect 4212 18232 4218 18284
rect 6564 18272 6592 18371
rect 8018 18368 8024 18380
rect 8076 18368 8082 18420
rect 8478 18408 8484 18420
rect 8439 18380 8484 18408
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 9582 18408 9588 18420
rect 9543 18380 9588 18408
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 9953 18411 10011 18417
rect 9953 18377 9965 18411
rect 9999 18408 10011 18411
rect 10134 18408 10140 18420
rect 9999 18380 10140 18408
rect 9999 18377 10011 18380
rect 9953 18371 10011 18377
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 10413 18411 10471 18417
rect 10413 18377 10425 18411
rect 10459 18408 10471 18411
rect 10502 18408 10508 18420
rect 10459 18380 10508 18408
rect 10459 18377 10471 18380
rect 10413 18371 10471 18377
rect 6638 18300 6644 18352
rect 6696 18340 6702 18352
rect 7745 18343 7803 18349
rect 7745 18340 7757 18343
rect 6696 18312 7757 18340
rect 6696 18300 6702 18312
rect 7745 18309 7757 18312
rect 7791 18309 7803 18343
rect 7745 18303 7803 18309
rect 8849 18343 8907 18349
rect 8849 18309 8861 18343
rect 8895 18340 8907 18343
rect 9858 18340 9864 18352
rect 8895 18312 9864 18340
rect 8895 18309 8907 18312
rect 8849 18303 8907 18309
rect 9858 18300 9864 18312
rect 9916 18300 9922 18352
rect 9217 18275 9275 18281
rect 6564 18244 6960 18272
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 2498 18204 2504 18216
rect 2455 18176 2504 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 2498 18164 2504 18176
rect 2556 18164 2562 18216
rect 3418 18204 3424 18216
rect 3379 18176 3424 18204
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 3878 18204 3884 18216
rect 3839 18176 3884 18204
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 4890 18164 4896 18216
rect 4948 18204 4954 18216
rect 4985 18207 5043 18213
rect 4985 18204 4997 18207
rect 4948 18176 4997 18204
rect 4948 18164 4954 18176
rect 4985 18173 4997 18176
rect 5031 18173 5043 18207
rect 5534 18204 5540 18216
rect 5495 18176 5540 18204
rect 4985 18167 5043 18173
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 5810 18164 5816 18216
rect 5868 18204 5874 18216
rect 6822 18204 6828 18216
rect 5868 18176 6828 18204
rect 5868 18164 5874 18176
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 2038 18136 2044 18148
rect 1951 18108 2044 18136
rect 2038 18096 2044 18108
rect 2096 18136 2102 18148
rect 5350 18136 5356 18148
rect 2096 18108 5356 18136
rect 2096 18096 2102 18108
rect 5350 18096 5356 18108
rect 5408 18096 5414 18148
rect 5718 18136 5724 18148
rect 5679 18108 5724 18136
rect 5718 18096 5724 18108
rect 5776 18096 5782 18148
rect 6932 18136 6960 18244
rect 9217 18241 9229 18275
rect 9263 18272 9275 18275
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9263 18244 9689 18272
rect 9263 18241 9275 18244
rect 9217 18235 9275 18241
rect 9677 18241 9689 18244
rect 9723 18272 9735 18275
rect 10428 18272 10456 18371
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 11238 18368 11244 18420
rect 11296 18408 11302 18420
rect 11333 18411 11391 18417
rect 11333 18408 11345 18411
rect 11296 18380 11345 18408
rect 11296 18368 11302 18380
rect 11333 18377 11345 18380
rect 11379 18377 11391 18411
rect 11333 18371 11391 18377
rect 11514 18272 11520 18284
rect 9723 18244 11520 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 9456 18207 9514 18213
rect 9456 18173 9468 18207
rect 9502 18204 9514 18207
rect 9766 18204 9772 18216
rect 9502 18176 9772 18204
rect 9502 18173 9514 18176
rect 9456 18167 9514 18173
rect 9766 18164 9772 18176
rect 9824 18164 9830 18216
rect 10410 18164 10416 18216
rect 10468 18204 10474 18216
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 10468 18176 10885 18204
rect 10468 18164 10474 18176
rect 10873 18173 10885 18176
rect 10919 18204 10931 18207
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 10919 18176 11713 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 12434 18204 12440 18216
rect 12395 18176 12440 18204
rect 11701 18167 11759 18173
rect 12434 18164 12440 18176
rect 12492 18204 12498 18216
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12492 18176 12909 18204
rect 12492 18164 12498 18176
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 12897 18167 12955 18173
rect 7146 18139 7204 18145
rect 7146 18136 7158 18139
rect 6932 18108 7158 18136
rect 7146 18105 7158 18108
rect 7192 18105 7204 18139
rect 7146 18099 7204 18105
rect 9309 18139 9367 18145
rect 9309 18105 9321 18139
rect 9355 18136 9367 18139
rect 9582 18136 9588 18148
rect 9355 18108 9588 18136
rect 9355 18105 9367 18108
rect 9309 18099 9367 18105
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 4430 18028 4436 18080
rect 4488 18068 4494 18080
rect 4525 18071 4583 18077
rect 4525 18068 4537 18071
rect 4488 18040 4537 18068
rect 4488 18028 4494 18040
rect 4525 18037 4537 18040
rect 4571 18037 4583 18071
rect 10686 18068 10692 18080
rect 10647 18040 10692 18068
rect 4525 18031 4583 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 11054 18068 11060 18080
rect 11015 18040 11060 18068
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 12618 18068 12624 18080
rect 12579 18040 12624 18068
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 3145 17867 3203 17873
rect 3145 17833 3157 17867
rect 3191 17864 3203 17867
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 3191 17836 3433 17864
rect 3191 17833 3203 17836
rect 3145 17827 3203 17833
rect 3421 17833 3433 17836
rect 3467 17864 3479 17867
rect 3878 17864 3884 17876
rect 3467 17836 3884 17864
rect 3467 17833 3479 17836
rect 3421 17827 3479 17833
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 4203 17867 4261 17873
rect 4203 17833 4215 17867
rect 4249 17864 4261 17867
rect 4798 17864 4804 17876
rect 4249 17836 4804 17864
rect 4249 17833 4261 17836
rect 4203 17827 4261 17833
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 5718 17824 5724 17876
rect 5776 17864 5782 17876
rect 6089 17867 6147 17873
rect 6089 17864 6101 17867
rect 5776 17836 6101 17864
rect 5776 17824 5782 17836
rect 6089 17833 6101 17836
rect 6135 17833 6147 17867
rect 6089 17827 6147 17833
rect 6549 17867 6607 17873
rect 6549 17833 6561 17867
rect 6595 17864 6607 17867
rect 6638 17864 6644 17876
rect 6595 17836 6644 17864
rect 6595 17833 6607 17836
rect 6549 17827 6607 17833
rect 6638 17824 6644 17836
rect 6696 17864 6702 17876
rect 9401 17867 9459 17873
rect 9401 17864 9413 17867
rect 6696 17836 6868 17864
rect 6696 17824 6702 17836
rect 3234 17756 3240 17808
rect 3292 17796 3298 17808
rect 4893 17799 4951 17805
rect 4893 17796 4905 17799
rect 3292 17768 4905 17796
rect 3292 17756 3298 17768
rect 4893 17765 4905 17768
rect 4939 17796 4951 17799
rect 5810 17796 5816 17808
rect 4939 17768 5672 17796
rect 5771 17768 5816 17796
rect 4939 17765 4951 17768
rect 4893 17759 4951 17765
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 3050 17728 3056 17740
rect 3007 17700 3056 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 3050 17688 3056 17700
rect 3108 17688 3114 17740
rect 4154 17737 4160 17740
rect 4132 17731 4160 17737
rect 4132 17697 4144 17731
rect 4132 17691 4160 17697
rect 4154 17688 4160 17691
rect 4212 17688 4218 17740
rect 5074 17728 5080 17740
rect 5035 17700 5080 17728
rect 5074 17688 5080 17700
rect 5132 17688 5138 17740
rect 5534 17728 5540 17740
rect 5495 17700 5540 17728
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 5644 17728 5672 17768
rect 5810 17756 5816 17768
rect 5868 17756 5874 17808
rect 6840 17805 6868 17836
rect 8220 17836 9413 17864
rect 6825 17799 6883 17805
rect 6825 17765 6837 17799
rect 6871 17765 6883 17799
rect 7374 17796 7380 17808
rect 7335 17768 7380 17796
rect 6825 17759 6883 17765
rect 7374 17756 7380 17768
rect 7432 17756 7438 17808
rect 8220 17805 8248 17836
rect 9401 17833 9413 17836
rect 9447 17864 9459 17867
rect 9582 17864 9588 17876
rect 9447 17836 9588 17864
rect 9447 17833 9459 17836
rect 9401 17827 9459 17833
rect 9582 17824 9588 17836
rect 9640 17824 9646 17876
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 10652 17836 13277 17864
rect 10652 17824 10658 17836
rect 13265 17833 13277 17836
rect 13311 17833 13323 17867
rect 13265 17827 13323 17833
rect 8113 17799 8171 17805
rect 8113 17765 8125 17799
rect 8159 17796 8171 17799
rect 8205 17799 8263 17805
rect 8205 17796 8217 17799
rect 8159 17768 8217 17796
rect 8159 17765 8171 17768
rect 8113 17759 8171 17765
rect 8205 17765 8217 17768
rect 8251 17765 8263 17799
rect 9766 17796 9772 17808
rect 9679 17768 9772 17796
rect 8205 17759 8263 17765
rect 6178 17728 6184 17740
rect 5644 17700 6184 17728
rect 6178 17688 6184 17700
rect 6236 17688 6242 17740
rect 9692 17737 9720 17768
rect 9766 17756 9772 17768
rect 9824 17796 9830 17808
rect 10686 17796 10692 17808
rect 9824 17768 10692 17796
rect 9824 17756 9830 17768
rect 10686 17756 10692 17768
rect 10744 17796 10750 17808
rect 10781 17799 10839 17805
rect 10781 17796 10793 17799
rect 10744 17768 10793 17796
rect 10744 17756 10750 17768
rect 10781 17765 10793 17768
rect 10827 17796 10839 17799
rect 10827 17768 12848 17796
rect 10827 17765 10839 17768
rect 10781 17759 10839 17765
rect 12820 17740 12848 17768
rect 8389 17731 8447 17737
rect 8389 17697 8401 17731
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 9953 17731 10011 17737
rect 9953 17697 9965 17731
rect 9999 17728 10011 17731
rect 11514 17728 11520 17740
rect 9999 17700 11284 17728
rect 11475 17700 11520 17728
rect 9999 17697 10011 17700
rect 9953 17691 10011 17697
rect 5626 17620 5632 17672
rect 5684 17660 5690 17672
rect 6733 17663 6791 17669
rect 6733 17660 6745 17663
rect 5684 17632 6745 17660
rect 5684 17620 5690 17632
rect 6733 17629 6745 17632
rect 6779 17629 6791 17663
rect 6733 17623 6791 17629
rect 8294 17620 8300 17672
rect 8352 17660 8358 17672
rect 8404 17660 8432 17691
rect 11256 17672 11284 17700
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 12802 17728 12808 17740
rect 12763 17700 12808 17728
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 13078 17728 13084 17740
rect 13039 17700 13084 17728
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 8352 17632 10149 17660
rect 8352 17620 8358 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 11238 17660 11244 17672
rect 11199 17632 11244 17660
rect 10137 17623 10195 17629
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 7745 17595 7803 17601
rect 7745 17561 7757 17595
rect 7791 17592 7803 17595
rect 8846 17592 8852 17604
rect 7791 17564 8852 17592
rect 7791 17561 7803 17564
rect 7745 17555 7803 17561
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 9769 17595 9827 17601
rect 9769 17561 9781 17595
rect 9815 17592 9827 17595
rect 9858 17592 9864 17604
rect 9815 17564 9864 17592
rect 9815 17561 9827 17564
rect 9769 17555 9827 17561
rect 9858 17552 9864 17564
rect 9916 17552 9922 17604
rect 12894 17592 12900 17604
rect 12855 17564 12900 17592
rect 12894 17552 12900 17564
rect 12952 17552 12958 17604
rect 2498 17524 2504 17536
rect 2459 17496 2504 17524
rect 2498 17484 2504 17496
rect 2556 17484 2562 17536
rect 4617 17527 4675 17533
rect 4617 17493 4629 17527
rect 4663 17524 4675 17527
rect 4706 17524 4712 17536
rect 4663 17496 4712 17524
rect 4663 17493 4675 17496
rect 4617 17487 4675 17493
rect 4706 17484 4712 17496
rect 4764 17484 4770 17536
rect 8478 17524 8484 17536
rect 8439 17496 8484 17524
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 10962 17524 10968 17536
rect 9732 17496 10968 17524
rect 9732 17484 9738 17496
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 4154 17320 4160 17332
rect 4115 17292 4160 17320
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5261 17323 5319 17329
rect 5261 17320 5273 17323
rect 5132 17292 5273 17320
rect 5132 17280 5138 17292
rect 5261 17289 5273 17292
rect 5307 17289 5319 17323
rect 5261 17283 5319 17289
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 5592 17292 5641 17320
rect 5592 17280 5598 17292
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 8294 17320 8300 17332
rect 8255 17292 8300 17320
rect 5629 17283 5687 17289
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 10045 17323 10103 17329
rect 10045 17320 10057 17323
rect 9916 17292 10057 17320
rect 9916 17280 9922 17292
rect 10045 17289 10057 17292
rect 10091 17320 10103 17323
rect 10413 17323 10471 17329
rect 10413 17320 10425 17323
rect 10091 17292 10425 17320
rect 10091 17289 10103 17292
rect 10045 17283 10103 17289
rect 10413 17289 10425 17292
rect 10459 17320 10471 17323
rect 10459 17292 10732 17320
rect 10459 17289 10471 17292
rect 10413 17283 10471 17289
rect 3050 17252 3056 17264
rect 3011 17224 3056 17252
rect 3050 17212 3056 17224
rect 3108 17212 3114 17264
rect 10704 17261 10732 17292
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11572 17292 11621 17320
rect 11572 17280 11578 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 12802 17280 12808 17332
rect 12860 17320 12866 17332
rect 13541 17323 13599 17329
rect 13541 17320 13553 17323
rect 12860 17292 13553 17320
rect 12860 17280 12866 17292
rect 13541 17289 13553 17292
rect 13587 17289 13599 17323
rect 13541 17283 13599 17289
rect 6273 17255 6331 17261
rect 6273 17221 6285 17255
rect 6319 17252 6331 17255
rect 10689 17255 10747 17261
rect 6319 17224 7696 17252
rect 6319 17221 6331 17224
rect 6273 17215 6331 17221
rect 3789 17187 3847 17193
rect 3789 17153 3801 17187
rect 3835 17184 3847 17187
rect 4614 17184 4620 17196
rect 3835 17156 4620 17184
rect 3835 17153 3847 17156
rect 3789 17147 3847 17153
rect 4540 17125 4568 17156
rect 4614 17144 4620 17156
rect 4672 17184 4678 17196
rect 5074 17184 5080 17196
rect 4672 17156 5080 17184
rect 4672 17144 4678 17156
rect 5074 17144 5080 17156
rect 5132 17144 5138 17196
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 6972 17156 7573 17184
rect 6972 17144 6978 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17085 4583 17119
rect 4706 17116 4712 17128
rect 4667 17088 4712 17116
rect 4525 17079 4583 17085
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 7101 17119 7159 17125
rect 7101 17085 7113 17119
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 4982 17048 4988 17060
rect 4943 17020 4988 17048
rect 4982 17008 4988 17020
rect 5040 17008 5046 17060
rect 6641 17051 6699 17057
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 7116 17048 7144 17079
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7377 17119 7435 17125
rect 7248 17088 7293 17116
rect 7248 17076 7254 17088
rect 7377 17085 7389 17119
rect 7423 17116 7435 17119
rect 7668 17116 7696 17224
rect 10689 17221 10701 17255
rect 10735 17221 10747 17255
rect 10689 17215 10747 17221
rect 13078 17212 13084 17264
rect 13136 17252 13142 17264
rect 13173 17255 13231 17261
rect 13173 17252 13185 17255
rect 13136 17224 13185 17252
rect 13136 17212 13142 17224
rect 13173 17221 13185 17224
rect 13219 17221 13231 17255
rect 13173 17215 13231 17221
rect 8570 17144 8576 17196
rect 8628 17184 8634 17196
rect 8628 17156 9076 17184
rect 8628 17144 8634 17156
rect 7742 17116 7748 17128
rect 7423 17088 7748 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8941 17119 8999 17125
rect 8941 17085 8953 17119
rect 8987 17085 8999 17119
rect 9048 17116 9076 17156
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 9582 17184 9588 17196
rect 9180 17156 9588 17184
rect 9180 17144 9186 17156
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 9048 17088 9505 17116
rect 8941 17079 8999 17085
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 10594 17116 10600 17128
rect 10555 17088 10600 17116
rect 9493 17079 9551 17085
rect 7558 17048 7564 17060
rect 6687 17020 7564 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 7558 17008 7564 17020
rect 7616 17048 7622 17060
rect 8294 17048 8300 17060
rect 7616 17020 8300 17048
rect 7616 17008 7622 17020
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 8846 17008 8852 17060
rect 8904 17048 8910 17060
rect 8956 17048 8984 17079
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10870 17116 10876 17128
rect 10783 17088 10876 17116
rect 10870 17076 10876 17088
rect 10928 17116 10934 17128
rect 11238 17116 11244 17128
rect 10928 17088 11244 17116
rect 10928 17076 10934 17088
rect 11238 17076 11244 17088
rect 11296 17076 11302 17128
rect 9674 17048 9680 17060
rect 8904 17020 9680 17048
rect 8904 17008 8910 17020
rect 9674 17008 9680 17020
rect 9732 17008 9738 17060
rect 9582 16980 9588 16992
rect 9543 16952 9588 16980
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 11054 16980 11060 16992
rect 11015 16952 11060 16980
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 4982 16736 4988 16788
rect 5040 16776 5046 16788
rect 5261 16779 5319 16785
rect 5261 16776 5273 16779
rect 5040 16748 5273 16776
rect 5040 16736 5046 16748
rect 5261 16745 5273 16748
rect 5307 16745 5319 16779
rect 5261 16739 5319 16745
rect 5626 16736 5632 16788
rect 5684 16776 5690 16788
rect 5813 16779 5871 16785
rect 5813 16776 5825 16779
rect 5684 16748 5825 16776
rect 5684 16736 5690 16748
rect 5813 16745 5825 16748
rect 5859 16745 5871 16779
rect 7190 16776 7196 16788
rect 7151 16748 7196 16776
rect 5813 16739 5871 16745
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 9122 16776 9128 16788
rect 8803 16748 9128 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 9122 16736 9128 16748
rect 9180 16776 9186 16788
rect 9398 16776 9404 16788
rect 9180 16748 9404 16776
rect 9180 16736 9186 16748
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 10781 16779 10839 16785
rect 10781 16745 10793 16779
rect 10827 16776 10839 16779
rect 10870 16776 10876 16788
rect 10827 16748 10876 16776
rect 10827 16745 10839 16748
rect 10781 16739 10839 16745
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16609 4307 16643
rect 4706 16640 4712 16652
rect 4667 16612 4712 16640
rect 4249 16603 4307 16609
rect 4264 16572 4292 16603
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 6086 16600 6092 16652
rect 6144 16640 6150 16652
rect 6641 16643 6699 16649
rect 6641 16640 6653 16643
rect 6144 16612 6653 16640
rect 6144 16600 6150 16612
rect 6641 16609 6653 16612
rect 6687 16640 6699 16643
rect 7208 16640 7236 16736
rect 9493 16711 9551 16717
rect 9493 16677 9505 16711
rect 9539 16708 9551 16711
rect 10796 16708 10824 16739
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 13679 16779 13737 16785
rect 13679 16776 13691 16779
rect 12492 16748 13691 16776
rect 12492 16736 12498 16748
rect 13679 16745 13691 16748
rect 13725 16745 13737 16779
rect 13679 16739 13737 16745
rect 9539 16680 10824 16708
rect 11977 16711 12035 16717
rect 9539 16677 9551 16680
rect 9493 16671 9551 16677
rect 11977 16677 11989 16711
rect 12023 16708 12035 16711
rect 12802 16708 12808 16720
rect 12023 16680 12808 16708
rect 12023 16677 12035 16680
rect 11977 16671 12035 16677
rect 12802 16668 12808 16680
rect 12860 16668 12866 16720
rect 7558 16640 7564 16652
rect 6687 16612 7236 16640
rect 7519 16612 7564 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 7742 16600 7748 16652
rect 7800 16640 7806 16652
rect 7837 16643 7895 16649
rect 7837 16640 7849 16643
rect 7800 16612 7849 16640
rect 7800 16600 7806 16612
rect 7837 16609 7849 16612
rect 7883 16640 7895 16643
rect 8018 16640 8024 16652
rect 7883 16612 8024 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 9950 16640 9956 16652
rect 9911 16612 9956 16640
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10594 16600 10600 16652
rect 10652 16640 10658 16652
rect 11057 16643 11115 16649
rect 11057 16640 11069 16643
rect 10652 16612 11069 16640
rect 10652 16600 10658 16612
rect 11057 16609 11069 16612
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 12434 16640 12440 16652
rect 11931 16612 12440 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 13538 16600 13544 16652
rect 13596 16649 13602 16652
rect 13596 16643 13634 16649
rect 13622 16609 13634 16643
rect 13596 16603 13634 16609
rect 13596 16600 13602 16603
rect 4430 16572 4436 16584
rect 4264 16544 4436 16572
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 4798 16572 4804 16584
rect 4759 16544 4804 16572
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16572 6791 16575
rect 7653 16575 7711 16581
rect 7653 16572 7665 16575
rect 6779 16544 7665 16572
rect 6779 16541 6791 16544
rect 6733 16535 6791 16541
rect 7653 16541 7665 16544
rect 7699 16572 7711 16575
rect 8202 16572 8208 16584
rect 7699 16544 8208 16572
rect 7699 16541 7711 16544
rect 7653 16535 7711 16541
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 10410 16572 10416 16584
rect 10371 16544 10416 16572
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 9766 16504 9772 16516
rect 9727 16476 9772 16504
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 3234 16192 3240 16244
rect 3292 16232 3298 16244
rect 3743 16235 3801 16241
rect 3743 16232 3755 16235
rect 3292 16204 3755 16232
rect 3292 16192 3298 16204
rect 3743 16201 3755 16204
rect 3789 16201 3801 16235
rect 3743 16195 3801 16201
rect 4525 16235 4583 16241
rect 4525 16201 4537 16235
rect 4571 16232 4583 16235
rect 5258 16232 5264 16244
rect 4571 16204 5264 16232
rect 4571 16201 4583 16204
rect 4525 16195 4583 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6086 16232 6092 16244
rect 6047 16204 6092 16232
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 7929 16235 7987 16241
rect 7929 16201 7941 16235
rect 7975 16232 7987 16235
rect 8202 16232 8208 16244
rect 7975 16204 8208 16232
rect 7975 16201 7987 16204
rect 7929 16195 7987 16201
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 10137 16235 10195 16241
rect 10137 16232 10149 16235
rect 9824 16204 10149 16232
rect 9824 16192 9830 16204
rect 10137 16201 10149 16204
rect 10183 16232 10195 16235
rect 10962 16232 10968 16244
rect 10183 16204 10968 16232
rect 10183 16201 10195 16204
rect 10137 16195 10195 16201
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 13538 16232 13544 16244
rect 13499 16204 13544 16232
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 6549 16167 6607 16173
rect 6549 16164 6561 16167
rect 4448 16136 6561 16164
rect 4448 16108 4476 16136
rect 6549 16133 6561 16136
rect 6595 16133 6607 16167
rect 6549 16127 6607 16133
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16096 4215 16099
rect 4430 16096 4436 16108
rect 4203 16068 4436 16096
rect 4203 16065 4215 16068
rect 4157 16059 4215 16065
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16096 4675 16099
rect 4982 16096 4988 16108
rect 4663 16068 4988 16096
rect 4663 16065 4675 16068
rect 4617 16059 4675 16065
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 3513 16031 3571 16037
rect 3513 15997 3525 16031
rect 3559 16028 3571 16031
rect 3640 16031 3698 16037
rect 3640 16028 3652 16031
rect 3559 16000 3652 16028
rect 3559 15997 3571 16000
rect 3513 15991 3571 15997
rect 3640 15997 3652 16000
rect 3686 16028 3698 16031
rect 4246 16028 4252 16040
rect 3686 16000 4252 16028
rect 3686 15997 3698 16000
rect 3640 15991 3698 15997
rect 4246 15988 4252 16000
rect 4304 15988 4310 16040
rect 6564 16028 6592 16127
rect 11238 16124 11244 16176
rect 11296 16164 11302 16176
rect 11974 16164 11980 16176
rect 11296 16136 11980 16164
rect 11296 16124 11302 16136
rect 11974 16124 11980 16136
rect 12032 16124 12038 16176
rect 9398 16096 9404 16108
rect 9359 16068 9404 16096
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16096 10931 16099
rect 11146 16096 11152 16108
rect 10919 16068 11152 16096
rect 10919 16065 10931 16068
rect 10873 16059 10931 16065
rect 11146 16056 11152 16068
rect 11204 16096 11210 16108
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 11204 16068 12449 16096
rect 11204 16056 11210 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6564 16000 6837 16028
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 7374 16028 7380 16040
rect 7335 16000 7380 16028
rect 6825 15991 6883 15997
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 8846 16028 8852 16040
rect 8807 16000 8852 16028
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 4979 15963 5037 15969
rect 4979 15929 4991 15963
rect 5025 15960 5037 15963
rect 5258 15960 5264 15972
rect 5025 15932 5264 15960
rect 5025 15929 5037 15932
rect 4979 15923 5037 15929
rect 5258 15920 5264 15932
rect 5316 15920 5322 15972
rect 8573 15963 8631 15969
rect 8573 15929 8585 15963
rect 8619 15960 8631 15963
rect 8754 15960 8760 15972
rect 8619 15932 8760 15960
rect 8619 15929 8631 15932
rect 8573 15923 8631 15929
rect 8754 15920 8760 15932
rect 8812 15960 8818 15972
rect 9398 15960 9404 15972
rect 8812 15932 9404 15960
rect 8812 15920 8818 15932
rect 9398 15920 9404 15932
rect 9456 15960 9462 15972
rect 9508 15960 9536 15991
rect 9456 15932 9536 15960
rect 9456 15920 9462 15932
rect 10962 15920 10968 15972
rect 11020 15960 11026 15972
rect 11517 15963 11575 15969
rect 11020 15932 11065 15960
rect 11020 15920 11026 15932
rect 11517 15929 11529 15963
rect 11563 15960 11575 15963
rect 11974 15960 11980 15972
rect 11563 15932 11980 15960
rect 11563 15929 11575 15932
rect 11517 15923 11575 15929
rect 11974 15920 11980 15932
rect 12032 15920 12038 15972
rect 5537 15895 5595 15901
rect 5537 15861 5549 15895
rect 5583 15892 5595 15895
rect 5902 15892 5908 15904
rect 5583 15864 5908 15892
rect 5583 15861 5595 15864
rect 5537 15855 5595 15861
rect 5902 15852 5908 15864
rect 5960 15852 5966 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 9582 15892 9588 15904
rect 9543 15864 9588 15892
rect 9582 15852 9588 15864
rect 9640 15852 9646 15904
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 10980 15892 11008 15920
rect 10735 15864 11008 15892
rect 11885 15895 11943 15901
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 11885 15861 11897 15895
rect 11931 15892 11943 15895
rect 12434 15892 12440 15904
rect 11931 15864 12440 15892
rect 11931 15861 11943 15864
rect 11885 15855 11943 15861
rect 12434 15852 12440 15864
rect 12492 15852 12498 15904
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 4341 15691 4399 15697
rect 4341 15657 4353 15691
rect 4387 15688 4399 15691
rect 4706 15688 4712 15700
rect 4387 15660 4712 15688
rect 4387 15657 4399 15660
rect 4341 15651 4399 15657
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 7745 15691 7803 15697
rect 7745 15688 7757 15691
rect 7616 15660 7757 15688
rect 7616 15648 7622 15660
rect 7745 15657 7757 15660
rect 7791 15657 7803 15691
rect 7745 15651 7803 15657
rect 9033 15691 9091 15697
rect 9033 15657 9045 15691
rect 9079 15688 9091 15691
rect 9490 15688 9496 15700
rect 9079 15660 9496 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 4979 15623 5037 15629
rect 4979 15589 4991 15623
rect 5025 15620 5037 15623
rect 5258 15620 5264 15632
rect 5025 15592 5264 15620
rect 5025 15589 5037 15592
rect 4979 15583 5037 15589
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 5902 15580 5908 15632
rect 5960 15620 5966 15632
rect 6546 15620 6552 15632
rect 5960 15592 6552 15620
rect 5960 15580 5966 15592
rect 6546 15580 6552 15592
rect 6604 15580 6610 15632
rect 8846 15620 8852 15632
rect 7944 15592 8852 15620
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4798 15552 4804 15564
rect 4663 15524 4804 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4798 15512 4804 15524
rect 4856 15552 4862 15564
rect 5534 15552 5540 15564
rect 4856 15524 5540 15552
rect 4856 15512 4862 15524
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 7944 15561 7972 15592
rect 8846 15580 8852 15592
rect 8904 15580 8910 15632
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 8018 15512 8024 15564
rect 8076 15552 8082 15564
rect 8205 15555 8263 15561
rect 8205 15552 8217 15555
rect 8076 15524 8217 15552
rect 8076 15512 8082 15524
rect 8205 15521 8217 15524
rect 8251 15552 8263 15555
rect 9048 15552 9076 15651
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 11146 15688 11152 15700
rect 11107 15660 11152 15688
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 10042 15580 10048 15632
rect 10100 15620 10106 15632
rect 10182 15623 10240 15629
rect 10182 15620 10194 15623
rect 10100 15592 10194 15620
rect 10100 15580 10106 15592
rect 10182 15589 10194 15592
rect 10228 15589 10240 15623
rect 11790 15620 11796 15632
rect 10182 15583 10240 15589
rect 10796 15592 11796 15620
rect 8251 15524 9076 15552
rect 8251 15521 8263 15524
rect 8205 15515 8263 15521
rect 9490 15512 9496 15564
rect 9548 15552 9554 15564
rect 9674 15552 9680 15564
rect 9548 15524 9680 15552
rect 9548 15512 9554 15524
rect 9674 15512 9680 15524
rect 9732 15552 9738 15564
rect 10796 15561 10824 15592
rect 11790 15580 11796 15592
rect 11848 15580 11854 15632
rect 11974 15580 11980 15632
rect 12032 15620 12038 15632
rect 13538 15620 13544 15632
rect 12032 15592 13544 15620
rect 12032 15580 12038 15592
rect 13538 15580 13544 15592
rect 13596 15580 13602 15632
rect 9861 15555 9919 15561
rect 9861 15552 9873 15555
rect 9732 15524 9873 15552
rect 9732 15512 9738 15524
rect 9861 15521 9873 15524
rect 9907 15521 9919 15555
rect 9861 15515 9919 15521
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15521 10839 15555
rect 10781 15515 10839 15521
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 4154 15484 4160 15496
rect 3007 15456 4160 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 4154 15444 4160 15456
rect 4212 15444 4218 15496
rect 6454 15484 6460 15496
rect 6415 15456 6460 15484
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 6914 15484 6920 15496
rect 6875 15456 6920 15484
rect 6914 15444 6920 15456
rect 6972 15444 6978 15496
rect 8110 15444 8116 15496
rect 8168 15484 8174 15496
rect 8389 15487 8447 15493
rect 8389 15484 8401 15487
rect 8168 15456 8401 15484
rect 8168 15444 8174 15456
rect 8389 15453 8401 15456
rect 8435 15453 8447 15487
rect 11698 15484 11704 15496
rect 11659 15456 11704 15484
rect 8389 15447 8447 15453
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 11974 15484 11980 15496
rect 11935 15456 11980 15484
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 5537 15419 5595 15425
rect 5537 15385 5549 15419
rect 5583 15416 5595 15419
rect 6822 15416 6828 15428
rect 5583 15388 6828 15416
rect 5583 15385 5595 15388
rect 5537 15379 5595 15385
rect 6822 15376 6828 15388
rect 6880 15376 6886 15428
rect 8021 15419 8079 15425
rect 8021 15385 8033 15419
rect 8067 15416 8079 15419
rect 8202 15416 8208 15428
rect 8067 15388 8208 15416
rect 8067 15385 8079 15388
rect 8021 15379 8079 15385
rect 8202 15376 8208 15388
rect 8260 15376 8266 15428
rect 5626 15308 5632 15360
rect 5684 15348 5690 15360
rect 6181 15351 6239 15357
rect 6181 15348 6193 15351
rect 5684 15320 6193 15348
rect 5684 15308 5690 15320
rect 6181 15317 6193 15320
rect 6227 15348 6239 15351
rect 6454 15348 6460 15360
rect 6227 15320 6460 15348
rect 6227 15317 6239 15320
rect 6181 15311 6239 15317
rect 6454 15308 6460 15320
rect 6512 15308 6518 15360
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 7374 15348 7380 15360
rect 7064 15320 7380 15348
rect 7064 15308 7070 15320
rect 7374 15308 7380 15320
rect 7432 15348 7438 15360
rect 7469 15351 7527 15357
rect 7469 15348 7481 15351
rect 7432 15320 7481 15348
rect 7432 15308 7438 15320
rect 7469 15317 7481 15320
rect 7515 15348 7527 15351
rect 8110 15348 8116 15360
rect 7515 15320 8116 15348
rect 7515 15317 7527 15320
rect 7469 15311 7527 15317
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 3881 15147 3939 15153
rect 3881 15113 3893 15147
rect 3927 15144 3939 15147
rect 4062 15144 4068 15156
rect 3927 15116 4068 15144
rect 3927 15113 3939 15116
rect 3881 15107 3939 15113
rect 4062 15104 4068 15116
rect 4120 15144 4126 15156
rect 5258 15144 5264 15156
rect 4120 15116 5264 15144
rect 4120 15104 4126 15116
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 5534 15144 5540 15156
rect 5495 15116 5540 15144
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 6546 15144 6552 15156
rect 6507 15116 6552 15144
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 7929 15147 7987 15153
rect 7929 15113 7941 15147
rect 7975 15144 7987 15147
rect 8202 15144 8208 15156
rect 7975 15116 8208 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 9398 15144 9404 15156
rect 8352 15116 8397 15144
rect 9359 15116 9404 15144
rect 8352 15104 8358 15116
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 10229 15147 10287 15153
rect 10229 15144 10241 15147
rect 9824 15116 10241 15144
rect 9824 15104 9830 15116
rect 10229 15113 10241 15116
rect 10275 15113 10287 15147
rect 11054 15144 11060 15156
rect 11015 15116 11060 15144
rect 10229 15107 10287 15113
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 3418 15076 3424 15088
rect 2700 15048 3424 15076
rect 2498 14900 2504 14952
rect 2556 14940 2562 14952
rect 2700 14949 2728 15048
rect 3418 15036 3424 15048
rect 3476 15036 3482 15088
rect 4706 15036 4712 15088
rect 4764 15076 4770 15088
rect 5905 15079 5963 15085
rect 5905 15076 5917 15079
rect 4764 15048 5917 15076
rect 4764 15036 4770 15048
rect 5905 15045 5917 15048
rect 5951 15045 5963 15079
rect 5905 15039 5963 15045
rect 6273 15079 6331 15085
rect 6273 15045 6285 15079
rect 6319 15076 6331 15079
rect 6638 15076 6644 15088
rect 6319 15048 6644 15076
rect 6319 15045 6331 15048
rect 6273 15039 6331 15045
rect 4338 15008 4344 15020
rect 2976 14980 4344 15008
rect 2976 14949 3004 14980
rect 4338 14968 4344 14980
rect 4396 15008 4402 15020
rect 4724 15008 4752 15036
rect 4396 14980 4752 15008
rect 4396 14968 4402 14980
rect 2685 14943 2743 14949
rect 2685 14940 2697 14943
rect 2556 14912 2697 14940
rect 2556 14900 2562 14912
rect 2685 14909 2697 14912
rect 2731 14909 2743 14943
rect 2685 14903 2743 14909
rect 2961 14943 3019 14949
rect 2961 14909 2973 14943
rect 3007 14909 3019 14943
rect 2961 14903 3019 14909
rect 3973 14943 4031 14949
rect 3973 14909 3985 14943
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14940 5779 14943
rect 6288 14940 6316 15039
rect 6638 15036 6644 15048
rect 6696 15036 6702 15088
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7193 15011 7251 15017
rect 7193 15008 7205 15011
rect 6972 14980 7205 15008
rect 6972 14968 6978 14980
rect 7193 14977 7205 14980
rect 7239 14977 7251 15011
rect 7193 14971 7251 14977
rect 8110 14968 8116 15020
rect 8168 15008 8174 15020
rect 8168 14980 8708 15008
rect 8168 14968 8174 14980
rect 8680 14952 8708 14980
rect 5767 14912 6316 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 2317 14875 2375 14881
rect 2317 14841 2329 14875
rect 2363 14872 2375 14875
rect 2976 14872 3004 14903
rect 2363 14844 3004 14872
rect 3145 14875 3203 14881
rect 2363 14841 2375 14844
rect 2317 14835 2375 14841
rect 3145 14841 3157 14875
rect 3191 14872 3203 14875
rect 3421 14875 3479 14881
rect 3421 14872 3433 14875
rect 3191 14844 3433 14872
rect 3191 14841 3203 14844
rect 3145 14835 3203 14841
rect 3421 14841 3433 14844
rect 3467 14872 3479 14875
rect 3988 14872 4016 14903
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 8389 14943 8447 14949
rect 8389 14940 8401 14943
rect 8352 14912 8401 14940
rect 8352 14900 8358 14912
rect 8389 14909 8401 14912
rect 8435 14909 8447 14943
rect 8389 14903 8447 14909
rect 8662 14900 8668 14952
rect 8720 14940 8726 14952
rect 8849 14943 8907 14949
rect 8849 14940 8861 14943
rect 8720 14912 8861 14940
rect 8720 14900 8726 14912
rect 8849 14909 8861 14912
rect 8895 14909 8907 14943
rect 8849 14903 8907 14909
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14940 10747 14943
rect 11425 14943 11483 14949
rect 11425 14940 11437 14943
rect 10735 14912 11437 14940
rect 10735 14909 10747 14912
rect 10689 14903 10747 14909
rect 11425 14909 11437 14912
rect 11471 14940 11483 14943
rect 11790 14940 11796 14952
rect 11471 14912 11796 14940
rect 11471 14909 11483 14912
rect 11425 14903 11483 14909
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 3467 14844 4016 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 4062 14832 4068 14884
rect 4120 14872 4126 14884
rect 4294 14875 4352 14881
rect 4294 14872 4306 14875
rect 4120 14844 4306 14872
rect 4120 14832 4126 14844
rect 4294 14841 4306 14844
rect 4340 14841 4352 14875
rect 4294 14835 4352 14841
rect 5810 14832 5816 14884
rect 5868 14872 5874 14884
rect 6917 14875 6975 14881
rect 6917 14872 6929 14875
rect 5868 14844 6929 14872
rect 5868 14832 5874 14844
rect 6917 14841 6929 14844
rect 6963 14841 6975 14875
rect 6917 14835 6975 14841
rect 7009 14875 7067 14881
rect 7009 14841 7021 14875
rect 7055 14841 7067 14875
rect 7009 14835 7067 14841
rect 4614 14764 4620 14816
rect 4672 14804 4678 14816
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 4672 14776 4905 14804
rect 4672 14764 4678 14776
rect 4893 14773 4905 14776
rect 4939 14773 4951 14807
rect 4893 14767 4951 14773
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 7024 14804 7052 14835
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 11330 14872 11336 14884
rect 10928 14844 11336 14872
rect 10928 14832 10934 14844
rect 11330 14832 11336 14844
rect 11388 14832 11394 14884
rect 11698 14832 11704 14884
rect 11756 14832 11762 14884
rect 8478 14804 8484 14816
rect 6880 14776 7052 14804
rect 8439 14776 8484 14804
rect 6880 14764 6886 14776
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9732 14776 9873 14804
rect 9732 14764 9738 14776
rect 9861 14773 9873 14776
rect 9907 14804 9919 14807
rect 10042 14804 10048 14816
rect 9907 14776 10048 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 11716 14804 11744 14832
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 10652 14776 12173 14804
rect 10652 14764 10658 14776
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 12161 14767 12219 14773
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 2498 14600 2504 14612
rect 2459 14572 2504 14600
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 3142 14560 3148 14612
rect 3200 14600 3206 14612
rect 5902 14600 5908 14612
rect 3200 14572 5908 14600
rect 3200 14560 3206 14572
rect 5902 14560 5908 14572
rect 5960 14560 5966 14612
rect 6822 14600 6828 14612
rect 6783 14572 6828 14600
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7193 14603 7251 14609
rect 7193 14569 7205 14603
rect 7239 14600 7251 14603
rect 8846 14600 8852 14612
rect 7239 14572 8852 14600
rect 7239 14569 7251 14572
rect 7193 14563 7251 14569
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 9490 14600 9496 14612
rect 9451 14572 9496 14600
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 9674 14560 9680 14612
rect 9732 14560 9738 14612
rect 4614 14492 4620 14544
rect 4672 14532 4678 14544
rect 4709 14535 4767 14541
rect 4709 14532 4721 14535
rect 4672 14504 4721 14532
rect 4672 14492 4678 14504
rect 4709 14501 4721 14504
rect 4755 14501 4767 14535
rect 4709 14495 4767 14501
rect 7558 14492 7564 14544
rect 7616 14541 7622 14544
rect 7616 14535 7664 14541
rect 7616 14501 7618 14535
rect 7652 14501 7664 14535
rect 9692 14532 9720 14560
rect 9998 14535 10056 14541
rect 9998 14532 10010 14535
rect 9692 14504 10010 14532
rect 7616 14495 7664 14501
rect 9998 14501 10010 14504
rect 10044 14501 10056 14535
rect 9998 14495 10056 14501
rect 7616 14492 7622 14495
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 6362 14464 6368 14476
rect 6319 14436 6368 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 6362 14424 6368 14436
rect 6420 14464 6426 14476
rect 6730 14464 6736 14476
rect 6420 14436 6736 14464
rect 6420 14424 6426 14436
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 7285 14467 7343 14473
rect 7285 14433 7297 14467
rect 7331 14464 7343 14467
rect 7742 14464 7748 14476
rect 7331 14436 7748 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 7742 14424 7748 14436
rect 7800 14464 7806 14476
rect 8478 14464 8484 14476
rect 7800 14436 8484 14464
rect 7800 14424 7806 14436
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9640 14436 9689 14464
rect 9640 14424 9646 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 11330 14424 11336 14476
rect 11388 14464 11394 14476
rect 11460 14467 11518 14473
rect 11460 14464 11472 14467
rect 11388 14436 11472 14464
rect 11388 14424 11394 14436
rect 11460 14433 11472 14436
rect 11506 14433 11518 14467
rect 11460 14427 11518 14433
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 4212 14368 4629 14396
rect 4212 14356 4218 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 4246 14288 4252 14340
rect 4304 14328 4310 14340
rect 4908 14328 4936 14359
rect 4304 14300 4936 14328
rect 4304 14288 4310 14300
rect 4982 14288 4988 14340
rect 5040 14328 5046 14340
rect 6457 14331 6515 14337
rect 6457 14328 6469 14331
rect 5040 14300 6469 14328
rect 5040 14288 5046 14300
rect 6457 14297 6469 14300
rect 6503 14328 6515 14331
rect 6822 14328 6828 14340
rect 6503 14300 6828 14328
rect 6503 14297 6515 14300
rect 6457 14291 6515 14297
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 5534 14260 5540 14272
rect 5495 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6089 14263 6147 14269
rect 6089 14260 6101 14263
rect 5868 14232 6101 14260
rect 5868 14220 5874 14232
rect 6089 14229 6101 14232
rect 6135 14229 6147 14263
rect 8202 14260 8208 14272
rect 8163 14232 8208 14260
rect 6089 14223 6147 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8573 14263 8631 14269
rect 8573 14229 8585 14263
rect 8619 14260 8631 14263
rect 8662 14260 8668 14272
rect 8619 14232 8668 14260
rect 8619 14229 8631 14232
rect 8573 14223 8631 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 10686 14260 10692 14272
rect 10643 14232 10692 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 11563 14263 11621 14269
rect 11563 14260 11575 14263
rect 11020 14232 11575 14260
rect 11020 14220 11026 14232
rect 11563 14229 11575 14232
rect 11609 14229 11621 14263
rect 11563 14223 11621 14229
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 4617 14059 4675 14065
rect 4617 14056 4629 14059
rect 4212 14028 4629 14056
rect 4212 14016 4218 14028
rect 4617 14025 4629 14028
rect 4663 14025 4675 14059
rect 4617 14019 4675 14025
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 5994 14056 6000 14068
rect 4764 14028 6000 14056
rect 4764 14016 4770 14028
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 6362 14056 6368 14068
rect 6323 14028 6368 14056
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 7193 14059 7251 14065
rect 7193 14025 7205 14059
rect 7239 14056 7251 14059
rect 7558 14056 7564 14068
rect 7239 14028 7564 14056
rect 7239 14025 7251 14028
rect 7193 14019 7251 14025
rect 7558 14016 7564 14028
rect 7616 14016 7622 14068
rect 9033 14059 9091 14065
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 9582 14056 9588 14068
rect 9079 14028 9588 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 10962 14056 10968 14068
rect 10923 14028 10968 14056
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 5810 13988 5816 14000
rect 5771 13960 5816 13988
rect 5810 13948 5816 13960
rect 5868 13948 5874 14000
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13920 3571 13923
rect 3559 13892 4108 13920
rect 3559 13889 3571 13892
rect 3513 13883 3571 13889
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 4080 13861 4108 13892
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 4212 13892 5273 13920
rect 4212 13880 4218 13892
rect 5261 13889 5273 13892
rect 5307 13920 5319 13923
rect 5534 13920 5540 13932
rect 5307 13892 5540 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 7098 13880 7104 13932
rect 7156 13920 7162 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 7156 13892 7297 13920
rect 7156 13880 7162 13892
rect 7285 13889 7297 13892
rect 7331 13920 7343 13923
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 7331 13892 8493 13920
rect 7331 13889 7343 13892
rect 7285 13883 7343 13889
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 9674 13920 9680 13932
rect 9635 13892 9680 13920
rect 8481 13883 8539 13889
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 10980 13920 11008 14016
rect 11330 13948 11336 14000
rect 11388 13988 11394 14000
rect 11425 13991 11483 13997
rect 11425 13988 11437 13991
rect 11388 13960 11437 13988
rect 11388 13948 11394 13960
rect 11425 13957 11437 13960
rect 11471 13957 11483 13991
rect 11425 13951 11483 13957
rect 9999 13892 11008 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 3605 13855 3663 13861
rect 3605 13852 3617 13855
rect 3476 13824 3617 13852
rect 3476 13812 3482 13824
rect 3605 13821 3617 13824
rect 3651 13821 3663 13855
rect 3605 13815 3663 13821
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4982 13852 4988 13864
rect 4111 13824 4988 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 8205 13855 8263 13861
rect 8205 13821 8217 13855
rect 8251 13852 8263 13855
rect 8294 13852 8300 13864
rect 8251 13824 8300 13852
rect 8251 13821 8263 13824
rect 8205 13815 8263 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 9401 13855 9459 13861
rect 9401 13821 9413 13855
rect 9447 13852 9459 13855
rect 9447 13824 9812 13852
rect 9447 13821 9459 13824
rect 9401 13815 9459 13821
rect 5353 13787 5411 13793
rect 5353 13753 5365 13787
rect 5399 13753 5411 13787
rect 5353 13747 5411 13753
rect 3878 13716 3884 13728
rect 3839 13688 3884 13716
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 5077 13719 5135 13725
rect 5077 13685 5089 13719
rect 5123 13716 5135 13719
rect 5368 13716 5396 13747
rect 7558 13744 7564 13796
rect 7616 13793 7622 13796
rect 7616 13787 7664 13793
rect 7616 13753 7618 13787
rect 7652 13753 7664 13787
rect 9784 13784 9812 13824
rect 10045 13787 10103 13793
rect 10045 13784 10057 13787
rect 9784 13756 10057 13784
rect 7616 13747 7664 13753
rect 10045 13753 10057 13756
rect 10091 13753 10103 13787
rect 10594 13784 10600 13796
rect 10555 13756 10600 13784
rect 10045 13747 10103 13753
rect 7616 13744 7622 13747
rect 5994 13716 6000 13728
rect 5123 13688 6000 13716
rect 5123 13685 5135 13688
rect 5077 13679 5135 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 10060 13716 10088 13747
rect 10594 13744 10600 13756
rect 10652 13744 10658 13796
rect 10686 13716 10692 13728
rect 10060 13688 10692 13716
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 3099 13515 3157 13521
rect 3099 13481 3111 13515
rect 3145 13512 3157 13515
rect 4062 13512 4068 13524
rect 3145 13484 4068 13512
rect 3145 13481 3157 13484
rect 3099 13475 3157 13481
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4614 13512 4620 13524
rect 4575 13484 4620 13512
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 7377 13515 7435 13521
rect 7377 13481 7389 13515
rect 7423 13512 7435 13515
rect 7558 13512 7564 13524
rect 7423 13484 7564 13512
rect 7423 13481 7435 13484
rect 7377 13475 7435 13481
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 7742 13512 7748 13524
rect 7703 13484 7748 13512
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 3418 13404 3424 13456
rect 3476 13444 3482 13456
rect 3605 13447 3663 13453
rect 3605 13444 3617 13447
rect 3476 13416 3617 13444
rect 3476 13404 3482 13416
rect 3605 13413 3617 13416
rect 3651 13413 3663 13447
rect 3605 13407 3663 13413
rect 5258 13404 5264 13456
rect 5316 13444 5322 13456
rect 5398 13447 5456 13453
rect 5398 13444 5410 13447
rect 5316 13416 5410 13444
rect 5316 13404 5322 13416
rect 5398 13413 5410 13416
rect 5444 13413 5456 13447
rect 8202 13444 8208 13456
rect 8163 13416 8208 13444
rect 5398 13407 5456 13413
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 10042 13444 10048 13456
rect 10003 13416 10048 13444
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 10594 13444 10600 13456
rect 10555 13416 10600 13444
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 2958 13336 2964 13388
rect 3016 13385 3022 13388
rect 3016 13379 3054 13385
rect 3042 13345 3054 13379
rect 3016 13339 3054 13345
rect 4132 13379 4190 13385
rect 4132 13345 4144 13379
rect 4178 13376 4190 13379
rect 4706 13376 4712 13388
rect 4178 13348 4712 13376
rect 4178 13345 4190 13348
rect 4132 13339 4190 13345
rect 3016 13336 3022 13339
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 11330 13336 11336 13388
rect 11388 13376 11394 13388
rect 11460 13379 11518 13385
rect 11460 13376 11472 13379
rect 11388 13348 11472 13376
rect 11388 13336 11394 13348
rect 11460 13345 11472 13348
rect 11506 13345 11518 13379
rect 11460 13339 11518 13345
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13277 5135 13311
rect 6822 13308 6828 13320
rect 6783 13280 6828 13308
rect 5077 13271 5135 13277
rect 4246 13249 4252 13252
rect 4203 13243 4252 13249
rect 4203 13240 4215 13243
rect 4159 13212 4215 13240
rect 4203 13209 4215 13212
rect 4249 13209 4252 13243
rect 4203 13203 4252 13209
rect 4246 13200 4252 13203
rect 4304 13240 4310 13252
rect 4982 13240 4988 13252
rect 4304 13212 4988 13240
rect 4304 13200 4310 13212
rect 4982 13200 4988 13212
rect 5040 13200 5046 13252
rect 4338 13132 4344 13184
rect 4396 13172 4402 13184
rect 4893 13175 4951 13181
rect 4893 13172 4905 13175
rect 4396 13144 4905 13172
rect 4396 13132 4402 13144
rect 4893 13141 4905 13144
rect 4939 13172 4951 13175
rect 5092 13172 5120 13271
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13308 8171 13311
rect 8570 13308 8576 13320
rect 8159 13280 8576 13308
rect 8159 13277 8171 13280
rect 8113 13271 8171 13277
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 8846 13308 8852 13320
rect 8803 13280 8852 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 9953 13311 10011 13317
rect 9953 13308 9965 13311
rect 9640 13280 9965 13308
rect 9640 13268 9646 13280
rect 9953 13277 9965 13280
rect 9999 13308 10011 13311
rect 11563 13311 11621 13317
rect 11563 13308 11575 13311
rect 9999 13280 11575 13308
rect 9999 13277 10011 13280
rect 9953 13271 10011 13277
rect 11563 13277 11575 13280
rect 11609 13277 11621 13311
rect 11563 13271 11621 13277
rect 5994 13172 6000 13184
rect 4939 13144 5120 13172
rect 5955 13144 6000 13172
rect 4939 13141 4951 13144
rect 4893 13135 4951 13141
rect 5994 13132 6000 13144
rect 6052 13132 6058 13184
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8812 13144 9045 13172
rect 8812 13132 8818 13144
rect 9033 13141 9045 13144
rect 9079 13141 9091 13175
rect 9033 13135 9091 13141
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 2958 12968 2964 12980
rect 2919 12940 2964 12968
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 3421 12971 3479 12977
rect 3421 12968 3433 12971
rect 3384 12940 3433 12968
rect 3384 12928 3390 12940
rect 3421 12937 3433 12940
rect 3467 12937 3479 12971
rect 6178 12968 6184 12980
rect 6139 12940 6184 12968
rect 3421 12931 3479 12937
rect 3436 12776 3464 12931
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 8110 12968 8116 12980
rect 8071 12940 8116 12968
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 8389 12971 8447 12977
rect 8389 12968 8401 12971
rect 8352 12940 8401 12968
rect 8352 12928 8358 12940
rect 8389 12937 8401 12940
rect 8435 12937 8447 12971
rect 8389 12931 8447 12937
rect 5077 12903 5135 12909
rect 5077 12869 5089 12903
rect 5123 12900 5135 12903
rect 5166 12900 5172 12912
rect 5123 12872 5172 12900
rect 5123 12869 5135 12872
rect 5077 12863 5135 12869
rect 5166 12860 5172 12872
rect 5224 12900 5230 12912
rect 5224 12872 6132 12900
rect 5224 12860 5230 12872
rect 4338 12832 4344 12844
rect 4299 12804 4344 12832
rect 4338 12792 4344 12804
rect 4396 12792 4402 12844
rect 4982 12792 4988 12844
rect 5040 12832 5046 12844
rect 5261 12835 5319 12841
rect 5261 12832 5273 12835
rect 5040 12804 5273 12832
rect 5040 12792 5046 12804
rect 5261 12801 5273 12804
rect 5307 12801 5319 12835
rect 5626 12832 5632 12844
rect 5587 12804 5632 12832
rect 5261 12795 5319 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 3418 12764 3424 12776
rect 3331 12736 3424 12764
rect 3418 12724 3424 12736
rect 3476 12764 3482 12776
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 3476 12736 3617 12764
rect 3476 12724 3482 12736
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 4154 12764 4160 12776
rect 4115 12736 4160 12764
rect 3605 12727 3663 12733
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 6104 12764 6132 12872
rect 6196 12832 6224 12928
rect 8478 12860 8484 12912
rect 8536 12900 8542 12912
rect 8536 12872 8892 12900
rect 8536 12860 8542 12872
rect 8864 12844 8892 12872
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 11425 12903 11483 12909
rect 11425 12900 11437 12903
rect 11388 12872 11437 12900
rect 11388 12860 11394 12872
rect 11425 12869 11437 12872
rect 11471 12869 11483 12903
rect 11425 12863 11483 12869
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6196 12804 6837 12832
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12832 8723 12835
rect 8754 12832 8760 12844
rect 8711 12804 8760 12832
rect 8711 12801 8723 12804
rect 8665 12795 8723 12801
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8904 12804 8953 12832
rect 8904 12792 8910 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10042 12832 10048 12844
rect 9999 12804 10048 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 10042 12792 10048 12804
rect 10100 12832 10106 12844
rect 10137 12835 10195 12841
rect 10137 12832 10149 12835
rect 10100 12804 10149 12832
rect 10100 12792 10106 12804
rect 10137 12801 10149 12804
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 6104 12736 6561 12764
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 10686 12764 10692 12776
rect 10647 12736 10692 12764
rect 6549 12727 6607 12733
rect 5353 12699 5411 12705
rect 5353 12665 5365 12699
rect 5399 12665 5411 12699
rect 6564 12696 6592 12727
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 7146 12699 7204 12705
rect 7146 12696 7158 12699
rect 6564 12668 7158 12696
rect 5353 12659 5411 12665
rect 7146 12665 7158 12668
rect 7192 12696 7204 12699
rect 7374 12696 7380 12708
rect 7192 12668 7380 12696
rect 7192 12665 7204 12668
rect 7146 12659 7204 12665
rect 4706 12628 4712 12640
rect 4667 12600 4712 12628
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 5368 12628 5396 12659
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 8757 12699 8815 12705
rect 8757 12696 8769 12699
rect 8352 12668 8769 12696
rect 8352 12656 8358 12668
rect 8757 12665 8769 12668
rect 8803 12665 8815 12699
rect 8757 12659 8815 12665
rect 10502 12656 10508 12708
rect 10560 12696 10566 12708
rect 11330 12696 11336 12708
rect 10560 12668 11336 12696
rect 10560 12656 10566 12668
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 5994 12628 6000 12640
rect 5368 12600 6000 12628
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 7742 12628 7748 12640
rect 7703 12600 7748 12628
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 3050 12384 3056 12436
rect 3108 12433 3114 12436
rect 3108 12427 3157 12433
rect 3108 12393 3111 12427
rect 3145 12393 3157 12427
rect 3108 12387 3157 12393
rect 3108 12384 3114 12387
rect 3326 12384 3332 12436
rect 3384 12424 3390 12436
rect 3510 12424 3516 12436
rect 3384 12396 3516 12424
rect 3384 12384 3390 12396
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 3697 12427 3755 12433
rect 3697 12393 3709 12427
rect 3743 12424 3755 12427
rect 4062 12424 4068 12436
rect 3743 12396 4068 12424
rect 3743 12393 3755 12396
rect 3697 12387 3755 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4246 12384 4252 12436
rect 4304 12424 4310 12436
rect 4709 12427 4767 12433
rect 4709 12424 4721 12427
rect 4304 12396 4721 12424
rect 4304 12384 4310 12396
rect 4709 12393 4721 12396
rect 4755 12393 4767 12427
rect 5994 12424 6000 12436
rect 5955 12396 6000 12424
rect 4709 12387 4767 12393
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 7745 12427 7803 12433
rect 7745 12424 7757 12427
rect 7708 12396 7757 12424
rect 7708 12384 7714 12396
rect 7745 12393 7757 12396
rect 7791 12424 7803 12427
rect 7791 12396 8524 12424
rect 7791 12393 7803 12396
rect 7745 12387 7803 12393
rect 4982 12316 4988 12368
rect 5040 12356 5046 12368
rect 5077 12359 5135 12365
rect 5077 12356 5089 12359
rect 5040 12328 5089 12356
rect 5040 12316 5046 12328
rect 5077 12325 5089 12328
rect 5123 12325 5135 12359
rect 5077 12319 5135 12325
rect 6641 12359 6699 12365
rect 6641 12325 6653 12359
rect 6687 12356 6699 12359
rect 7006 12356 7012 12368
rect 6687 12328 7012 12356
rect 6687 12325 6699 12328
rect 6641 12319 6699 12325
rect 7006 12316 7012 12328
rect 7064 12356 7070 12368
rect 8202 12356 8208 12368
rect 7064 12328 7788 12356
rect 8163 12328 8208 12356
rect 7064 12316 7070 12328
rect 7760 12300 7788 12328
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 8496 12356 8524 12396
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8628 12396 9045 12424
rect 8628 12384 8634 12396
rect 9033 12393 9045 12396
rect 9079 12424 9091 12427
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 9079 12396 9229 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9217 12393 9229 12396
rect 9263 12393 9275 12427
rect 9217 12387 9275 12393
rect 9493 12427 9551 12433
rect 9493 12393 9505 12427
rect 9539 12424 9551 12427
rect 9582 12424 9588 12436
rect 9539 12396 9588 12424
rect 9539 12393 9551 12396
rect 9493 12387 9551 12393
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 9769 12427 9827 12433
rect 9769 12393 9781 12427
rect 9815 12393 9827 12427
rect 10686 12424 10692 12436
rect 10647 12396 10692 12424
rect 9769 12387 9827 12393
rect 9784 12356 9812 12387
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 8496 12328 9812 12356
rect 11974 12316 11980 12368
rect 12032 12356 12038 12368
rect 12434 12356 12440 12368
rect 12032 12328 12440 12356
rect 12032 12316 12038 12328
rect 12434 12316 12440 12328
rect 12492 12316 12498 12368
rect 3050 12297 3056 12300
rect 3028 12291 3056 12297
rect 3028 12257 3040 12291
rect 3028 12251 3056 12257
rect 3050 12248 3056 12251
rect 3108 12248 3114 12300
rect 7742 12248 7748 12300
rect 7800 12248 7806 12300
rect 9950 12288 9956 12300
rect 9911 12260 9956 12288
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 11308 12291 11366 12297
rect 11308 12257 11320 12291
rect 11354 12288 11366 12291
rect 12250 12288 12256 12300
rect 11354 12260 12256 12288
rect 11354 12257 11366 12260
rect 11308 12251 11366 12257
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 4985 12223 5043 12229
rect 4985 12220 4997 12223
rect 4856 12192 4997 12220
rect 4856 12180 4862 12192
rect 4985 12189 4997 12192
rect 5031 12189 5043 12223
rect 5626 12220 5632 12232
rect 5587 12192 5632 12220
rect 4985 12183 5043 12189
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 6822 12220 6828 12232
rect 6595 12192 6828 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8570 12220 8576 12232
rect 8159 12192 8576 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 8570 12180 8576 12192
rect 8628 12220 8634 12232
rect 8628 12192 9352 12220
rect 8628 12180 8634 12192
rect 7098 12152 7104 12164
rect 7011 12124 7104 12152
rect 7098 12112 7104 12124
rect 7156 12152 7162 12164
rect 8478 12152 8484 12164
rect 7156 12124 8484 12152
rect 7156 12112 7162 12124
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 8665 12155 8723 12161
rect 8665 12121 8677 12155
rect 8711 12152 8723 12155
rect 8754 12152 8760 12164
rect 8711 12124 8760 12152
rect 8711 12121 8723 12124
rect 8665 12115 8723 12121
rect 8754 12112 8760 12124
rect 8812 12112 8818 12164
rect 9324 12152 9352 12192
rect 11379 12155 11437 12161
rect 11379 12152 11391 12155
rect 9324 12124 11391 12152
rect 11379 12121 11391 12124
rect 11425 12121 11437 12155
rect 11379 12115 11437 12121
rect 9217 12087 9275 12093
rect 9217 12053 9229 12087
rect 9263 12084 9275 12087
rect 10042 12084 10048 12096
rect 9263 12056 10048 12084
rect 9263 12053 9275 12056
rect 9217 12047 9275 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 3050 11880 3056 11892
rect 3011 11852 3056 11880
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 4982 11880 4988 11892
rect 4663 11852 4988 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 6549 11883 6607 11889
rect 6549 11849 6561 11883
rect 6595 11880 6607 11883
rect 6822 11880 6828 11892
rect 6595 11852 6828 11880
rect 6595 11849 6607 11852
rect 6549 11843 6607 11849
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7006 11880 7012 11892
rect 6967 11852 7012 11880
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 7469 11883 7527 11889
rect 7469 11880 7481 11883
rect 7432 11852 7481 11880
rect 7432 11840 7438 11852
rect 7469 11849 7481 11852
rect 7515 11849 7527 11883
rect 7469 11843 7527 11849
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 8260 11852 8585 11880
rect 8260 11840 8266 11852
rect 8573 11849 8585 11852
rect 8619 11880 8631 11883
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8619 11852 8861 11880
rect 8619 11849 8631 11852
rect 8573 11843 8631 11849
rect 8849 11849 8861 11852
rect 8895 11880 8907 11883
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 8895 11852 9137 11880
rect 8895 11849 8907 11852
rect 8849 11843 8907 11849
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9125 11843 9183 11849
rect 9309 11883 9367 11889
rect 9309 11849 9321 11883
rect 9355 11880 9367 11883
rect 10134 11880 10140 11892
rect 9355 11852 10140 11880
rect 9355 11849 9367 11852
rect 9309 11843 9367 11849
rect 4614 11744 4620 11756
rect 3804 11716 4620 11744
rect 3804 11685 3832 11716
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3467 11648 3801 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 4062 11676 4068 11688
rect 4023 11648 4068 11676
rect 3789 11639 3847 11645
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4246 11608 4252 11620
rect 4207 11580 4252 11608
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 5000 11540 5028 11840
rect 8662 11772 8668 11824
rect 8720 11812 8726 11824
rect 9324 11812 9352 11843
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 10962 11840 10968 11892
rect 11020 11880 11026 11892
rect 11422 11880 11428 11892
rect 11020 11852 11428 11880
rect 11020 11840 11026 11852
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 10042 11812 10048 11824
rect 8720 11784 9352 11812
rect 10003 11784 10048 11812
rect 8720 11772 8726 11784
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 5258 11744 5264 11756
rect 5215 11716 5264 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 5258 11704 5264 11716
rect 5316 11744 5322 11756
rect 6089 11747 6147 11753
rect 6089 11744 6101 11747
rect 5316 11716 6101 11744
rect 5316 11704 5322 11716
rect 6089 11713 6101 11716
rect 6135 11713 6147 11747
rect 7650 11744 7656 11756
rect 7611 11716 7656 11744
rect 6089 11707 6147 11713
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11744 9551 11747
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 9539 11716 10793 11744
rect 9539 11713 9551 11716
rect 9493 11707 9551 11713
rect 10781 11713 10793 11716
rect 10827 11744 10839 11747
rect 11103 11747 11161 11753
rect 11103 11744 11115 11747
rect 10827 11716 11115 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11103 11713 11115 11716
rect 11149 11713 11161 11747
rect 11103 11707 11161 11713
rect 10962 11636 10968 11688
rect 11020 11685 11026 11688
rect 11020 11679 11058 11685
rect 11046 11645 11058 11679
rect 11020 11639 11058 11645
rect 11020 11636 11026 11639
rect 5261 11611 5319 11617
rect 5261 11577 5273 11611
rect 5307 11577 5319 11611
rect 5810 11608 5816 11620
rect 5771 11580 5816 11608
rect 5261 11571 5319 11577
rect 5074 11540 5080 11552
rect 4987 11512 5080 11540
rect 5074 11500 5080 11512
rect 5132 11540 5138 11552
rect 5276 11540 5304 11571
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 7374 11568 7380 11620
rect 7432 11608 7438 11620
rect 7974 11611 8032 11617
rect 7974 11608 7986 11611
rect 7432 11580 7986 11608
rect 7432 11568 7438 11580
rect 7974 11577 7986 11580
rect 8020 11577 8032 11611
rect 7974 11571 8032 11577
rect 9125 11611 9183 11617
rect 9125 11577 9137 11611
rect 9171 11608 9183 11611
rect 9490 11608 9496 11620
rect 9171 11580 9496 11608
rect 9171 11577 9183 11580
rect 9125 11571 9183 11577
rect 9490 11568 9496 11580
rect 9548 11608 9554 11620
rect 9585 11611 9643 11617
rect 9585 11608 9597 11611
rect 9548 11580 9597 11608
rect 9548 11568 9554 11580
rect 9585 11577 9597 11580
rect 9631 11577 9643 11611
rect 9585 11571 9643 11577
rect 5132 11512 5304 11540
rect 5132 11500 5138 11512
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10413 11543 10471 11549
rect 10413 11540 10425 11543
rect 10008 11512 10425 11540
rect 10008 11500 10014 11512
rect 10413 11509 10425 11512
rect 10459 11509 10471 11543
rect 10413 11503 10471 11509
rect 11885 11543 11943 11549
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 12066 11540 12072 11552
rect 11931 11512 12072 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 12066 11500 12072 11512
rect 12124 11540 12130 11552
rect 12250 11540 12256 11552
rect 12124 11512 12256 11540
rect 12124 11500 12130 11512
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 3605 11339 3663 11345
rect 3605 11305 3617 11339
rect 3651 11336 3663 11339
rect 4062 11336 4068 11348
rect 3651 11308 4068 11336
rect 3651 11305 3663 11308
rect 3605 11299 3663 11305
rect 3620 11268 3648 11299
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 5132 11308 5181 11336
rect 5132 11296 5138 11308
rect 5169 11305 5181 11308
rect 5215 11305 5227 11339
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 5169 11299 5227 11305
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 9490 11336 9496 11348
rect 9451 11308 9496 11336
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 2976 11240 3648 11268
rect 2976 11212 3004 11240
rect 4338 11228 4344 11280
rect 4396 11268 4402 11280
rect 4611 11271 4669 11277
rect 4611 11268 4623 11271
rect 4396 11240 4623 11268
rect 4396 11228 4402 11240
rect 4611 11237 4623 11240
rect 4657 11268 4669 11271
rect 4657 11240 5212 11268
rect 4657 11237 4669 11240
rect 4611 11231 4669 11237
rect 5184 11212 5212 11240
rect 7374 11228 7380 11280
rect 7432 11268 7438 11280
rect 7606 11271 7664 11277
rect 7606 11268 7618 11271
rect 7432 11240 7618 11268
rect 7432 11228 7438 11240
rect 7606 11237 7618 11240
rect 7652 11237 7664 11271
rect 9858 11268 9864 11280
rect 9819 11240 9864 11268
rect 7606 11231 7664 11237
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 10042 11228 10048 11280
rect 10100 11268 10106 11280
rect 10413 11271 10471 11277
rect 10413 11268 10425 11271
rect 10100 11240 10425 11268
rect 10100 11228 10106 11240
rect 10413 11237 10425 11240
rect 10459 11237 10471 11271
rect 11422 11268 11428 11280
rect 11383 11240 11428 11268
rect 10413 11231 10471 11237
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2958 11200 2964 11212
rect 2871 11172 2964 11200
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 3145 11203 3203 11209
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 4154 11200 4160 11212
rect 3191 11172 4160 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 5166 11160 5172 11212
rect 5224 11160 5230 11212
rect 6178 11160 6184 11212
rect 6236 11200 6242 11212
rect 6308 11203 6366 11209
rect 6308 11200 6320 11203
rect 6236 11172 6320 11200
rect 6236 11160 6242 11172
rect 6308 11169 6320 11172
rect 6354 11169 6366 11203
rect 6308 11163 6366 11169
rect 4246 11132 4252 11144
rect 4159 11104 4252 11132
rect 4246 11092 4252 11104
rect 4304 11132 4310 11144
rect 5442 11132 5448 11144
rect 4304 11104 5448 11132
rect 4304 11092 4310 11104
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 7282 11132 7288 11144
rect 7243 11104 7288 11132
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 10594 11132 10600 11144
rect 9815 11104 10600 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11101 11391 11135
rect 11606 11132 11612 11144
rect 11567 11104 11612 11132
rect 11333 11095 11391 11101
rect 3050 11024 3056 11076
rect 3108 11064 3114 11076
rect 3878 11064 3884 11076
rect 3108 11036 3884 11064
rect 3108 11024 3114 11036
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4798 11064 4804 11076
rect 4080 11036 4804 11064
rect 4080 11008 4108 11036
rect 4798 11024 4804 11036
rect 4856 11064 4862 11076
rect 5537 11067 5595 11073
rect 5537 11064 5549 11067
rect 4856 11036 5549 11064
rect 4856 11024 4862 11036
rect 5537 11033 5549 11036
rect 5583 11033 5595 11067
rect 5537 11027 5595 11033
rect 6411 11067 6469 11073
rect 6411 11033 6423 11067
rect 6457 11064 6469 11067
rect 6822 11064 6828 11076
rect 6457 11036 6828 11064
rect 6457 11033 6469 11036
rect 6411 11027 6469 11033
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 7300 11064 7328 11092
rect 11348 11064 11376 11095
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 11514 11064 11520 11076
rect 7300 11036 8340 11064
rect 11348 11036 11520 11064
rect 4062 10956 4068 11008
rect 4120 10956 4126 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 8205 10999 8263 11005
rect 8205 10996 8217 10999
rect 8168 10968 8217 10996
rect 8168 10956 8174 10968
rect 8205 10965 8217 10968
rect 8251 10965 8263 10999
rect 8312 10996 8340 11036
rect 11514 11024 11520 11036
rect 11572 11024 11578 11076
rect 8386 10996 8392 11008
rect 8312 10968 8392 10996
rect 8205 10959 8263 10965
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 2958 10792 2964 10804
rect 2915 10764 2964 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 3559 10795 3617 10801
rect 3559 10761 3571 10795
rect 3605 10792 3617 10795
rect 4062 10792 4068 10804
rect 3605 10764 4068 10792
rect 3605 10761 3617 10764
rect 3559 10755 3617 10761
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4338 10792 4344 10804
rect 4299 10764 4344 10792
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5592 10764 5641 10792
rect 5592 10752 5598 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 7374 10792 7380 10804
rect 7335 10764 7380 10792
rect 5629 10755 5687 10761
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 8386 10752 8392 10804
rect 8444 10792 8450 10804
rect 8665 10795 8723 10801
rect 8665 10792 8677 10795
rect 8444 10764 8677 10792
rect 8444 10752 8450 10764
rect 8665 10761 8677 10764
rect 8711 10761 8723 10795
rect 8665 10755 8723 10761
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 9916 10764 10241 10792
rect 9916 10752 9922 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10594 10792 10600 10804
rect 10555 10764 10600 10792
rect 10229 10755 10287 10761
rect 10594 10752 10600 10764
rect 10652 10792 10658 10804
rect 10919 10795 10977 10801
rect 10919 10792 10931 10795
rect 10652 10764 10931 10792
rect 10652 10752 10658 10764
rect 10919 10761 10931 10764
rect 10965 10761 10977 10795
rect 10919 10755 10977 10761
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11609 10795 11667 10801
rect 11609 10792 11621 10795
rect 11480 10764 11621 10792
rect 11480 10752 11486 10764
rect 11609 10761 11621 10764
rect 11655 10761 11667 10795
rect 11609 10755 11667 10761
rect 4706 10684 4712 10736
rect 4764 10724 4770 10736
rect 9398 10724 9404 10736
rect 4764 10696 9404 10724
rect 4764 10684 4770 10696
rect 9398 10684 9404 10696
rect 9456 10684 9462 10736
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4212 10628 4445 10656
rect 4212 10616 4218 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10656 10011 10659
rect 10042 10656 10048 10668
rect 9999 10628 10048 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 3488 10591 3546 10597
rect 3488 10557 3500 10591
rect 3534 10588 3546 10591
rect 7469 10591 7527 10597
rect 3534 10560 3924 10588
rect 3534 10557 3546 10560
rect 3488 10551 3546 10557
rect 3896 10464 3924 10560
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7558 10588 7564 10600
rect 7515 10560 7564 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8435 10560 9168 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 4338 10480 4344 10532
rect 4396 10520 4402 10532
rect 4706 10520 4712 10532
rect 4396 10492 4712 10520
rect 4396 10480 4402 10492
rect 4706 10480 4712 10492
rect 4764 10529 4770 10532
rect 4764 10523 4812 10529
rect 4764 10489 4766 10523
rect 4800 10489 4812 10523
rect 4764 10483 4812 10489
rect 4764 10480 4770 10483
rect 7374 10480 7380 10532
rect 7432 10520 7438 10532
rect 7790 10523 7848 10529
rect 7790 10520 7802 10523
rect 7432 10492 7802 10520
rect 7432 10480 7438 10492
rect 7790 10489 7802 10492
rect 7836 10489 7848 10523
rect 7790 10483 7848 10489
rect 2406 10452 2412 10464
rect 2367 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 3878 10452 3884 10464
rect 3839 10424 3884 10452
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 5350 10452 5356 10464
rect 5311 10424 5356 10452
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 6178 10452 6184 10464
rect 5776 10424 6184 10452
rect 5776 10412 5782 10424
rect 6178 10412 6184 10424
rect 6236 10452 6242 10464
rect 9140 10461 9168 10560
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 10816 10591 10874 10597
rect 10816 10588 10828 10591
rect 10376 10560 10828 10588
rect 10376 10548 10382 10560
rect 10816 10557 10828 10560
rect 10862 10588 10874 10591
rect 11241 10591 11299 10597
rect 11241 10588 11253 10591
rect 10862 10560 11253 10588
rect 10862 10557 10874 10560
rect 10816 10551 10874 10557
rect 11241 10557 11253 10560
rect 11287 10557 11299 10591
rect 11241 10551 11299 10557
rect 9306 10520 9312 10532
rect 9267 10492 9312 10520
rect 9306 10480 9312 10492
rect 9364 10480 9370 10532
rect 9401 10523 9459 10529
rect 9401 10489 9413 10523
rect 9447 10520 9459 10523
rect 9490 10520 9496 10532
rect 9447 10492 9496 10520
rect 9447 10489 9459 10492
rect 9401 10483 9459 10489
rect 6273 10455 6331 10461
rect 6273 10452 6285 10455
rect 6236 10424 6285 10452
rect 6236 10412 6242 10424
rect 6273 10421 6285 10424
rect 6319 10421 6331 10455
rect 6273 10415 6331 10421
rect 9125 10455 9183 10461
rect 9125 10421 9137 10455
rect 9171 10452 9183 10455
rect 9416 10452 9444 10483
rect 9490 10480 9496 10492
rect 9548 10480 9554 10532
rect 9171 10424 9444 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 11977 10455 12035 10461
rect 11977 10452 11989 10455
rect 11572 10424 11989 10452
rect 11572 10412 11578 10424
rect 11977 10421 11989 10424
rect 12023 10421 12035 10455
rect 11977 10415 12035 10421
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 3099 10251 3157 10257
rect 3099 10217 3111 10251
rect 3145 10248 3157 10251
rect 3970 10248 3976 10260
rect 3145 10220 3976 10248
rect 3145 10217 3157 10220
rect 3099 10211 3157 10217
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 4212 10220 5089 10248
rect 4212 10208 4218 10220
rect 5077 10217 5089 10220
rect 5123 10217 5135 10251
rect 5077 10211 5135 10217
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 7432 10220 7481 10248
rect 7432 10208 7438 10220
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 9306 10248 9312 10260
rect 9267 10220 9312 10248
rect 7469 10211 7527 10217
rect 9306 10208 9312 10220
rect 9364 10248 9370 10260
rect 9815 10251 9873 10257
rect 9815 10248 9827 10251
rect 9364 10220 9827 10248
rect 9364 10208 9370 10220
rect 9815 10217 9827 10220
rect 9861 10217 9873 10251
rect 9815 10211 9873 10217
rect 4706 10180 4712 10192
rect 4667 10152 4712 10180
rect 4706 10140 4712 10152
rect 4764 10140 4770 10192
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 5445 10183 5503 10189
rect 5445 10180 5457 10183
rect 5408 10152 5457 10180
rect 5408 10140 5414 10152
rect 5445 10149 5457 10152
rect 5491 10149 5503 10183
rect 5445 10143 5503 10149
rect 8110 10140 8116 10192
rect 8168 10180 8174 10192
rect 8205 10183 8263 10189
rect 8205 10180 8217 10183
rect 8168 10152 8217 10180
rect 8168 10140 8174 10152
rect 8205 10149 8217 10152
rect 8251 10149 8263 10183
rect 8754 10180 8760 10192
rect 8715 10152 8760 10180
rect 8205 10143 8263 10149
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 3050 10121 3056 10124
rect 3028 10115 3056 10121
rect 3028 10081 3040 10115
rect 3028 10075 3056 10081
rect 3050 10072 3056 10075
rect 3108 10072 3114 10124
rect 4300 10115 4358 10121
rect 4300 10081 4312 10115
rect 4346 10112 4358 10115
rect 4522 10112 4528 10124
rect 4346 10084 4528 10112
rect 4346 10081 4358 10084
rect 4300 10075 4358 10081
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 9766 10121 9772 10124
rect 9744 10115 9772 10121
rect 9744 10081 9756 10115
rect 9824 10112 9830 10124
rect 10778 10112 10784 10124
rect 9824 10084 10784 10112
rect 9744 10075 9772 10081
rect 9766 10072 9772 10075
rect 9824 10072 9830 10084
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4387 10047 4445 10053
rect 4387 10044 4399 10047
rect 4120 10016 4399 10044
rect 4120 10004 4126 10016
rect 4387 10013 4399 10016
rect 4433 10044 4445 10047
rect 5353 10047 5411 10053
rect 5353 10044 5365 10047
rect 4433 10016 5365 10044
rect 4433 10013 4445 10016
rect 4387 10007 4445 10013
rect 5353 10013 5365 10016
rect 5399 10013 5411 10047
rect 5626 10044 5632 10056
rect 5587 10016 5632 10044
rect 5353 10007 5411 10013
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 6972 10016 8125 10044
rect 6972 10004 6978 10016
rect 8113 10013 8125 10016
rect 8159 10044 8171 10047
rect 8386 10044 8392 10056
rect 8159 10016 8392 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 4522 9936 4528 9988
rect 4580 9976 4586 9988
rect 7466 9976 7472 9988
rect 4580 9948 7472 9976
rect 4580 9936 4586 9948
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7616 9880 7849 9908
rect 7616 9868 7622 9880
rect 7837 9877 7849 9880
rect 7883 9877 7895 9911
rect 7837 9871 7895 9877
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4617 9707 4675 9713
rect 4617 9704 4629 9707
rect 4580 9676 4629 9704
rect 4580 9664 4586 9676
rect 4617 9673 4629 9676
rect 4663 9673 4675 9707
rect 8110 9704 8116 9716
rect 8071 9676 8116 9704
rect 4617 9667 4675 9673
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8202 9664 8208 9716
rect 8260 9704 8266 9716
rect 8294 9704 8300 9716
rect 8260 9676 8300 9704
rect 8260 9664 8266 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 10410 9704 10416 9716
rect 10284 9676 10416 9704
rect 10284 9664 10290 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 4062 9636 4068 9648
rect 4023 9608 4068 9636
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 5810 9636 5816 9648
rect 5771 9608 5816 9636
rect 5810 9596 5816 9608
rect 5868 9596 5874 9648
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 9217 9639 9275 9645
rect 9217 9636 9229 9639
rect 8444 9608 9229 9636
rect 8444 9596 8450 9608
rect 9217 9605 9229 9608
rect 9263 9605 9275 9639
rect 9217 9599 9275 9605
rect 11974 9596 11980 9648
rect 12032 9636 12038 9648
rect 13814 9636 13820 9648
rect 12032 9608 13820 9636
rect 12032 9596 12038 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 6546 9568 6552 9580
rect 6507 9540 6552 9568
rect 6546 9528 6552 9540
rect 6604 9568 6610 9580
rect 7558 9568 7564 9580
rect 6604 9540 6868 9568
rect 7519 9540 7564 9568
rect 6604 9528 6610 9540
rect 4208 9503 4266 9509
rect 4208 9469 4220 9503
rect 4254 9500 4266 9503
rect 5074 9500 5080 9512
rect 4254 9472 5080 9500
rect 4254 9469 4266 9472
rect 4208 9463 4266 9469
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 6840 9509 6868 9540
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8527 9571 8585 9577
rect 8527 9537 8539 9571
rect 8573 9568 8585 9571
rect 9582 9568 9588 9580
rect 8573 9540 9588 9568
rect 8573 9537 8585 9540
rect 8527 9531 8585 9537
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 7190 9500 7196 9512
rect 6871 9472 7196 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9469 7435 9503
rect 8386 9500 8392 9512
rect 8350 9472 8392 9500
rect 7377 9463 7435 9469
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 4295 9435 4353 9441
rect 4295 9432 4307 9435
rect 3743 9404 4307 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 4295 9401 4307 9404
rect 4341 9432 4353 9435
rect 5261 9435 5319 9441
rect 5261 9432 5273 9435
rect 4341 9404 5273 9432
rect 4341 9401 4353 9404
rect 4295 9395 4353 9401
rect 5261 9401 5273 9404
rect 5307 9401 5319 9435
rect 5261 9395 5319 9401
rect 5350 9392 5356 9444
rect 5408 9432 5414 9444
rect 6273 9435 6331 9441
rect 5408 9404 5453 9432
rect 5408 9392 5414 9404
rect 6273 9401 6285 9435
rect 6319 9432 6331 9435
rect 7098 9432 7104 9444
rect 6319 9404 7104 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 7098 9392 7104 9404
rect 7156 9432 7162 9444
rect 7392 9432 7420 9463
rect 8386 9460 8392 9472
rect 8444 9509 8450 9512
rect 8444 9503 8498 9509
rect 8444 9469 8452 9503
rect 8486 9500 8498 9503
rect 8846 9500 8852 9512
rect 8486 9472 8852 9500
rect 8486 9469 8498 9472
rect 8444 9463 8498 9469
rect 8444 9460 8450 9463
rect 8846 9460 8852 9472
rect 8904 9500 8910 9512
rect 8904 9472 8984 9500
rect 8904 9460 8910 9472
rect 8662 9432 8668 9444
rect 7156 9404 8668 9432
rect 7156 9392 7162 9404
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 8956 9441 8984 9472
rect 8941 9435 8999 9441
rect 8941 9401 8953 9435
rect 8987 9432 8999 9435
rect 10134 9432 10140 9444
rect 8987 9404 10140 9432
rect 8987 9401 8999 9404
rect 8941 9395 8999 9401
rect 10134 9392 10140 9404
rect 10192 9392 10198 9444
rect 3050 9364 3056 9376
rect 3011 9336 3056 9364
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 8570 9364 8576 9376
rect 3384 9336 8576 9364
rect 3384 9324 3390 9336
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 9766 9364 9772 9376
rect 9727 9336 9772 9364
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 5408 9132 5641 9160
rect 5408 9120 5414 9132
rect 5629 9129 5641 9132
rect 5675 9160 5687 9163
rect 5997 9163 6055 9169
rect 5997 9160 6009 9163
rect 5675 9132 6009 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 5997 9129 6009 9132
rect 6043 9129 6055 9163
rect 5997 9123 6055 9129
rect 4614 9092 4620 9104
rect 4540 9064 4620 9092
rect 4540 9033 4568 9064
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 6457 9095 6515 9101
rect 6457 9061 6469 9095
rect 6503 9092 6515 9095
rect 7282 9092 7288 9104
rect 6503 9064 7144 9092
rect 7243 9064 7288 9092
rect 6503 9061 6515 9064
rect 6457 9055 6515 9061
rect 7116 9036 7144 9064
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 4525 9027 4583 9033
rect 4525 8993 4537 9027
rect 4571 8993 4583 9027
rect 4706 9024 4712 9036
rect 4667 8996 4712 9024
rect 4525 8987 4583 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 6549 9027 6607 9033
rect 6549 9024 6561 9027
rect 6236 8996 6561 9024
rect 6236 8984 6242 8996
rect 6549 8993 6561 8996
rect 6595 8993 6607 9027
rect 7098 9024 7104 9036
rect 7059 8996 7104 9024
rect 6549 8987 6607 8993
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 8113 9027 8171 9033
rect 8113 8993 8125 9027
rect 8159 9024 8171 9027
rect 8294 9024 8300 9036
rect 8159 8996 8300 9024
rect 8159 8993 8171 8996
rect 8113 8987 8171 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 4798 8956 4804 8968
rect 4759 8928 4804 8956
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 8297 8891 8355 8897
rect 8297 8888 8309 8891
rect 5368 8860 8309 8888
rect 5368 8832 5396 8860
rect 8297 8857 8309 8860
rect 8343 8888 8355 8891
rect 8573 8891 8631 8897
rect 8573 8888 8585 8891
rect 8343 8860 8585 8888
rect 8343 8857 8355 8860
rect 8297 8851 8355 8857
rect 8573 8857 8585 8860
rect 8619 8888 8631 8891
rect 8754 8888 8760 8900
rect 8619 8860 8760 8888
rect 8619 8857 8631 8860
rect 8573 8851 8631 8857
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 5350 8820 5356 8832
rect 5311 8792 5356 8820
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 7650 8820 7656 8832
rect 7611 8792 7656 8820
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8720 8792 8953 8820
rect 8720 8780 8726 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 4430 8576 4436 8628
rect 4488 8616 4494 8628
rect 4985 8619 5043 8625
rect 4985 8616 4997 8619
rect 4488 8588 4997 8616
rect 4488 8576 4494 8588
rect 4985 8585 4997 8588
rect 5031 8585 5043 8619
rect 4985 8579 5043 8585
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8294 8616 8300 8628
rect 8251 8588 8300 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8480 3571 8483
rect 4448 8480 4476 8576
rect 4614 8548 4620 8560
rect 4575 8520 4620 8548
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 3559 8452 4476 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 3896 8421 3924 8452
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 4246 8412 4252 8424
rect 4203 8384 4252 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 4246 8372 4252 8384
rect 4304 8412 4310 8424
rect 4706 8412 4712 8424
rect 4304 8384 4712 8412
rect 4304 8372 4310 8384
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 5000 8412 5028 8579
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7650 8480 7656 8492
rect 6871 8452 7656 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 7650 8440 7656 8452
rect 7708 8480 7714 8492
rect 9125 8483 9183 8489
rect 9125 8480 9137 8483
rect 7708 8452 9137 8480
rect 7708 8440 7714 8452
rect 9125 8449 9137 8452
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 5000 8384 5181 8412
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5350 8372 5356 8424
rect 5408 8412 5414 8424
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 5408 8384 5641 8412
rect 5408 8372 5414 8384
rect 5629 8381 5641 8384
rect 5675 8381 5687 8415
rect 6178 8412 6184 8424
rect 6139 8384 6184 8412
rect 5629 8375 5687 8381
rect 6178 8372 6184 8384
rect 6236 8372 6242 8424
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 8662 8412 8668 8424
rect 6687 8384 6868 8412
rect 8623 8384 8668 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 4338 8344 4344 8356
rect 4299 8316 4344 8344
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 5905 8347 5963 8353
rect 5905 8313 5917 8347
rect 5951 8344 5963 8347
rect 6730 8344 6736 8356
rect 5951 8316 6736 8344
rect 5951 8313 5963 8316
rect 5905 8307 5963 8313
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 6840 8344 6868 8384
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8812 8384 9045 8412
rect 8812 8372 8818 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 7187 8347 7245 8353
rect 7187 8344 7199 8347
rect 6840 8316 7199 8344
rect 7187 8313 7199 8316
rect 7233 8344 7245 8347
rect 7374 8344 7380 8356
rect 7233 8316 7380 8344
rect 7233 8313 7245 8316
rect 7187 8307 7245 8313
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 7745 8279 7803 8285
rect 7745 8276 7757 8279
rect 6696 8248 7757 8276
rect 6696 8236 6702 8248
rect 7745 8245 7757 8248
rect 7791 8245 7803 8279
rect 7745 8239 7803 8245
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 3237 8075 3295 8081
rect 3237 8041 3249 8075
rect 3283 8072 3295 8075
rect 3510 8072 3516 8084
rect 3283 8044 3516 8072
rect 3283 8041 3295 8044
rect 3237 8035 3295 8041
rect 3510 8032 3516 8044
rect 3568 8072 3574 8084
rect 3697 8075 3755 8081
rect 3697 8072 3709 8075
rect 3568 8044 3709 8072
rect 3568 8032 3574 8044
rect 3697 8041 3709 8044
rect 3743 8072 3755 8075
rect 4246 8072 4252 8084
rect 3743 8044 4252 8072
rect 3743 8041 3755 8044
rect 3697 8035 3755 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4798 8072 4804 8084
rect 4759 8044 4804 8072
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7708 8044 7757 8072
rect 7708 8032 7714 8044
rect 7745 8041 7757 8044
rect 7791 8072 7803 8075
rect 9769 8075 9827 8081
rect 9769 8072 9781 8075
rect 7791 8044 9781 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 9769 8041 9781 8044
rect 9815 8041 9827 8075
rect 9769 8035 9827 8041
rect 6638 8004 6644 8016
rect 6599 7976 6644 8004
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 8202 8004 8208 8016
rect 8163 7976 8208 8004
rect 8202 7964 8208 7976
rect 8260 7964 8266 8016
rect 8754 7964 8760 8016
rect 8812 8004 8818 8016
rect 8812 7976 10180 8004
rect 8812 7964 8818 7976
rect 4890 7936 4896 7948
rect 4851 7908 4896 7936
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 5350 7936 5356 7948
rect 5263 7908 5356 7936
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 5276 7868 5304 7908
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 9950 7936 9956 7948
rect 9911 7908 9956 7936
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10152 7945 10180 7976
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7905 10195 7939
rect 10137 7899 10195 7905
rect 5442 7868 5448 7880
rect 4304 7840 5304 7868
rect 5403 7840 5448 7868
rect 4304 7828 4310 7840
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 6822 7868 6828 7880
rect 6595 7840 6828 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7006 7868 7012 7880
rect 6967 7840 7012 7868
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 8110 7868 8116 7880
rect 8071 7840 8116 7868
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 9306 7868 9312 7880
rect 8803 7840 9312 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 9490 7732 9496 7744
rect 9451 7704 9496 7732
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 6638 7488 6644 7540
rect 6696 7528 6702 7540
rect 7009 7531 7067 7537
rect 7009 7528 7021 7531
rect 6696 7500 7021 7528
rect 6696 7488 6702 7500
rect 7009 7497 7021 7500
rect 7055 7497 7067 7531
rect 7009 7491 7067 7497
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 7432 7500 7481 7528
rect 7432 7488 7438 7500
rect 7469 7497 7481 7500
rect 7515 7497 7527 7531
rect 7469 7491 7527 7497
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8573 7531 8631 7537
rect 8573 7528 8585 7531
rect 8260 7500 8585 7528
rect 8260 7488 8266 7500
rect 8573 7497 8585 7500
rect 8619 7528 8631 7531
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 8619 7500 8861 7528
rect 8619 7497 8631 7500
rect 8573 7491 8631 7497
rect 8849 7497 8861 7500
rect 8895 7497 8907 7531
rect 8849 7491 8907 7497
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 4614 7460 4620 7472
rect 4028 7432 4620 7460
rect 4028 7420 4034 7432
rect 4614 7420 4620 7432
rect 4672 7420 4678 7472
rect 6549 7463 6607 7469
rect 6549 7429 6561 7463
rect 6595 7460 6607 7463
rect 6822 7460 6828 7472
rect 6595 7432 6828 7460
rect 6595 7429 6607 7432
rect 6549 7423 6607 7429
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 4430 7392 4436 7404
rect 3436 7364 4436 7392
rect 3436 7336 3464 7364
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 4798 7392 4804 7404
rect 4755 7364 4804 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7324 3111 7327
rect 3418 7324 3424 7336
rect 3099 7296 3424 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 3605 7327 3663 7333
rect 3605 7324 3617 7327
rect 3568 7296 3617 7324
rect 3568 7284 3574 7296
rect 3605 7293 3617 7296
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 3881 7259 3939 7265
rect 3881 7225 3893 7259
rect 3927 7256 3939 7259
rect 4062 7256 4068 7268
rect 3927 7228 4068 7256
rect 3927 7225 3939 7228
rect 3881 7219 3939 7225
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 5074 7265 5080 7268
rect 4617 7259 4675 7265
rect 4617 7225 4629 7259
rect 4663 7256 4675 7259
rect 5071 7256 5080 7265
rect 4663 7228 5080 7256
rect 4663 7225 4675 7228
rect 4617 7219 4675 7225
rect 5071 7219 5080 7228
rect 5074 7216 5080 7219
rect 5132 7216 5138 7268
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 7834 7256 7840 7268
rect 7432 7228 7840 7256
rect 7432 7216 7438 7228
rect 7834 7216 7840 7228
rect 7892 7256 7898 7268
rect 7974 7259 8032 7265
rect 7974 7256 7986 7259
rect 7892 7228 7986 7256
rect 7892 7216 7898 7228
rect 7974 7225 7986 7228
rect 8020 7225 8032 7259
rect 8864 7256 8892 7491
rect 9950 7488 9956 7540
rect 10008 7528 10014 7540
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 10008 7500 10425 7528
rect 10008 7488 10014 7500
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 10413 7491 10471 7497
rect 9490 7392 9496 7404
rect 9403 7364 9496 7392
rect 9490 7352 9496 7364
rect 9548 7392 9554 7404
rect 11103 7395 11161 7401
rect 11103 7392 11115 7395
rect 9548 7364 11115 7392
rect 9548 7352 9554 7364
rect 11103 7361 11115 7364
rect 11149 7361 11161 7395
rect 11103 7355 11161 7361
rect 11016 7327 11074 7333
rect 11016 7293 11028 7327
rect 11062 7324 11074 7327
rect 11422 7324 11428 7336
rect 11062 7296 11428 7324
rect 11062 7293 11074 7296
rect 11016 7287 11074 7293
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 9490 7256 9496 7268
rect 8864 7228 9496 7256
rect 7974 7219 8032 7225
rect 9490 7216 9496 7228
rect 9548 7256 9554 7268
rect 9585 7259 9643 7265
rect 9585 7256 9597 7259
rect 9548 7228 9597 7256
rect 9548 7216 9554 7228
rect 9585 7225 9597 7228
rect 9631 7225 9643 7259
rect 9585 7219 9643 7225
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 9732 7228 10149 7256
rect 9732 7216 9738 7228
rect 10137 7225 10149 7228
rect 10183 7225 10195 7259
rect 10137 7219 10195 7225
rect 4246 7188 4252 7200
rect 4207 7160 4252 7188
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 5629 7191 5687 7197
rect 5629 7188 5641 7191
rect 5592 7160 5641 7188
rect 5592 7148 5598 7160
rect 5629 7157 5641 7160
rect 5675 7157 5687 7191
rect 5629 7151 5687 7157
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 8812 7160 9229 7188
rect 8812 7148 8818 7160
rect 9217 7157 9229 7160
rect 9263 7157 9275 7191
rect 9217 7151 9275 7157
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 3510 6944 3516 6996
rect 3568 6984 3574 6996
rect 3970 6984 3976 6996
rect 3568 6956 3976 6984
rect 3568 6944 3574 6956
rect 3970 6944 3976 6956
rect 4028 6984 4034 6996
rect 4433 6987 4491 6993
rect 4433 6984 4445 6987
rect 4028 6956 4445 6984
rect 4028 6944 4034 6956
rect 4433 6953 4445 6956
rect 4479 6953 4491 6987
rect 4890 6984 4896 6996
rect 4851 6956 4896 6984
rect 4433 6947 4491 6953
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 5902 6984 5908 6996
rect 5224 6956 5908 6984
rect 5224 6944 5230 6956
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 9490 6984 9496 6996
rect 9451 6956 9496 6984
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 2961 6851 3019 6857
rect 2731 6820 2912 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 2884 6712 2912 6820
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 3528 6848 3556 6944
rect 5074 6876 5080 6928
rect 5132 6916 5138 6928
rect 7834 6925 7840 6928
rect 5582 6919 5640 6925
rect 5582 6916 5594 6919
rect 5132 6888 5594 6916
rect 5132 6876 5138 6888
rect 5582 6885 5594 6888
rect 5628 6885 5640 6919
rect 7831 6916 7840 6925
rect 7795 6888 7840 6916
rect 5582 6879 5640 6885
rect 7831 6879 7840 6888
rect 7834 6876 7840 6879
rect 7892 6876 7898 6928
rect 9858 6916 9864 6928
rect 9819 6888 9864 6916
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 3007 6820 3556 6848
rect 4249 6851 4307 6857
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 4249 6817 4261 6851
rect 4295 6817 4307 6851
rect 4249 6811 4307 6817
rect 3142 6780 3148 6792
rect 3103 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 4264 6780 4292 6811
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 4396 6820 6469 6848
rect 4396 6808 4402 6820
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 6972 6820 7481 6848
rect 6972 6808 6978 6820
rect 7469 6817 7481 6820
rect 7515 6848 7527 6851
rect 8202 6848 8208 6860
rect 7515 6820 8208 6848
rect 7515 6817 7527 6820
rect 7469 6811 7527 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 4522 6780 4528 6792
rect 4264 6752 4528 6780
rect 4522 6740 4528 6752
rect 4580 6780 4586 6792
rect 4982 6780 4988 6792
rect 4580 6752 4988 6780
rect 4580 6740 4586 6752
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 5261 6743 5319 6749
rect 9692 6752 9781 6780
rect 2958 6712 2964 6724
rect 2871 6684 2964 6712
rect 2958 6672 2964 6684
rect 3016 6712 3022 6724
rect 3326 6712 3332 6724
rect 3016 6684 3332 6712
rect 3016 6672 3022 6684
rect 3326 6672 3332 6684
rect 3384 6672 3390 6724
rect 5276 6656 5304 6743
rect 9692 6724 9720 6752
rect 9769 6749 9781 6752
rect 9815 6749 9827 6783
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 9769 6743 9827 6749
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 8168 6684 8800 6712
rect 8168 6672 8174 6684
rect 8772 6656 8800 6684
rect 9674 6672 9680 6724
rect 9732 6672 9738 6724
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 5258 6644 5264 6656
rect 4212 6616 5264 6644
rect 4212 6604 4218 6616
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 6052 6616 6193 6644
rect 6052 6604 6058 6616
rect 6181 6613 6193 6616
rect 6227 6613 6239 6647
rect 6181 6607 6239 6613
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8570 6644 8576 6656
rect 8435 6616 8576 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 2547 6443 2605 6449
rect 2547 6409 2559 6443
rect 2593 6440 2605 6443
rect 2682 6440 2688 6452
rect 2593 6412 2688 6440
rect 2593 6409 2605 6412
rect 2547 6403 2605 6409
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 2958 6440 2964 6452
rect 2919 6412 2964 6440
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3234 6440 3240 6452
rect 3195 6412 3240 6440
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 4522 6440 4528 6452
rect 4483 6412 4528 6440
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 5258 6400 5264 6452
rect 5316 6440 5322 6452
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 5316 6412 6193 6440
rect 5316 6400 5322 6412
rect 6181 6409 6193 6412
rect 6227 6409 6239 6443
rect 6181 6403 6239 6409
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 7374 6440 7380 6452
rect 6687 6412 7380 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 4893 6375 4951 6381
rect 4893 6341 4905 6375
rect 4939 6372 4951 6375
rect 5074 6372 5080 6384
rect 4939 6344 5080 6372
rect 4939 6341 4951 6344
rect 4893 6335 4951 6341
rect 5074 6332 5080 6344
rect 5132 6372 5138 6384
rect 6656 6372 6684 6403
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 8628 6412 8953 6440
rect 8628 6400 8634 6412
rect 8941 6409 8953 6412
rect 8987 6440 8999 6443
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 8987 6412 9045 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 9033 6409 9045 6412
rect 9079 6409 9091 6443
rect 9033 6403 9091 6409
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 9732 6412 10609 6440
rect 9732 6400 9738 6412
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 5132 6344 6684 6372
rect 8389 6375 8447 6381
rect 5132 6332 5138 6344
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 3510 6304 3516 6316
rect 2363 6276 3516 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 3510 6264 3516 6276
rect 3568 6304 3574 6316
rect 3568 6276 4016 6304
rect 3568 6264 3574 6276
rect 3988 6248 4016 6276
rect 4338 6264 4344 6316
rect 4396 6304 4402 6316
rect 4985 6307 5043 6313
rect 4985 6304 4997 6307
rect 4396 6276 4997 6304
rect 4396 6264 4402 6276
rect 4985 6273 4997 6276
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 2498 6245 2504 6248
rect 2476 6239 2504 6245
rect 2476 6205 2488 6239
rect 2476 6199 2504 6205
rect 2498 6196 2504 6199
rect 2556 6196 2562 6248
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3292 6208 3433 6236
rect 3292 6196 3298 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3970 6236 3976 6248
rect 3931 6208 3976 6236
rect 3421 6199 3479 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5368 6180 5396 6344
rect 8389 6341 8401 6375
rect 8435 6372 8447 6375
rect 9858 6372 9864 6384
rect 8435 6344 9864 6372
rect 8435 6341 8447 6344
rect 8389 6335 8447 6341
rect 9858 6332 9864 6344
rect 9916 6372 9922 6384
rect 10229 6375 10287 6381
rect 10229 6372 10241 6375
rect 9916 6344 10241 6372
rect 9916 6332 9922 6344
rect 10229 6341 10241 6344
rect 10275 6341 10287 6375
rect 10229 6335 10287 6341
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6304 7530 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 7524 6276 8677 6304
rect 7524 6264 7530 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 9674 6304 9680 6316
rect 9635 6276 9680 6304
rect 8665 6267 8723 6273
rect 9674 6264 9680 6276
rect 9732 6304 9738 6316
rect 10042 6304 10048 6316
rect 9732 6276 10048 6304
rect 9732 6264 9738 6276
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 4154 6168 4160 6180
rect 4115 6140 4160 6168
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 5350 6177 5356 6180
rect 5347 6168 5356 6177
rect 5263 6140 5356 6168
rect 5347 6131 5356 6140
rect 5350 6128 5356 6131
rect 5408 6128 5414 6180
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 7790 6171 7848 6177
rect 7790 6168 7802 6171
rect 7432 6140 7802 6168
rect 7432 6128 7438 6140
rect 7790 6137 7802 6140
rect 7836 6137 7848 6171
rect 9306 6168 9312 6180
rect 9267 6140 9312 6168
rect 7790 6131 7848 6137
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 9401 6171 9459 6177
rect 9401 6137 9413 6171
rect 9447 6137 9459 6171
rect 9401 6131 9459 6137
rect 5902 6100 5908 6112
rect 5863 6072 5908 6100
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 8941 6103 8999 6109
rect 8941 6069 8953 6103
rect 8987 6100 8999 6103
rect 9416 6100 9444 6131
rect 8987 6072 9444 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 2498 5896 2504 5908
rect 2459 5868 2504 5896
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 3510 5896 3516 5908
rect 3471 5868 3516 5896
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 5350 5896 5356 5908
rect 5311 5868 5356 5896
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 7282 5896 7288 5908
rect 7243 5868 7288 5896
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 8202 5896 8208 5908
rect 8163 5868 8208 5896
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 9815 5899 9873 5905
rect 9815 5896 9827 5899
rect 8812 5868 9827 5896
rect 8812 5856 8818 5868
rect 9815 5865 9827 5868
rect 9861 5865 9873 5899
rect 9815 5859 9873 5865
rect 4430 5828 4436 5840
rect 4264 5800 4436 5828
rect 4264 5769 4292 5800
rect 4430 5788 4436 5800
rect 4488 5788 4494 5840
rect 5813 5831 5871 5837
rect 5813 5797 5825 5831
rect 5859 5828 5871 5831
rect 5902 5828 5908 5840
rect 5859 5800 5908 5828
rect 5859 5797 5871 5800
rect 5813 5791 5871 5797
rect 5902 5788 5908 5800
rect 5960 5828 5966 5840
rect 6178 5828 6184 5840
rect 5960 5800 6184 5828
rect 5960 5788 5966 5800
rect 6178 5788 6184 5800
rect 6236 5788 6242 5840
rect 4249 5763 4307 5769
rect 4249 5729 4261 5763
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 4396 5732 4537 5760
rect 4396 5720 4402 5732
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 7190 5760 7196 5772
rect 7151 5732 7196 5760
rect 4525 5723 4583 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7653 5763 7711 5769
rect 7653 5729 7665 5763
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 4798 5692 4804 5704
rect 4759 5664 4804 5692
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5692 5779 5695
rect 6086 5692 6092 5704
rect 5767 5664 6092 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7668 5692 7696 5723
rect 9674 5720 9680 5772
rect 9732 5769 9738 5772
rect 9732 5763 9770 5769
rect 9758 5729 9770 5763
rect 9732 5723 9770 5729
rect 9732 5720 9738 5723
rect 6972 5664 7696 5692
rect 6972 5652 6978 5664
rect 5626 5584 5632 5636
rect 5684 5624 5690 5636
rect 6273 5627 6331 5633
rect 6273 5624 6285 5627
rect 5684 5596 6285 5624
rect 5684 5584 5690 5596
rect 6273 5593 6285 5596
rect 6319 5593 6331 5627
rect 6273 5587 6331 5593
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4890 5556 4896 5568
rect 4120 5528 4896 5556
rect 4120 5516 4126 5528
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 9217 5559 9275 5565
rect 9217 5556 9229 5559
rect 8812 5528 9229 5556
rect 8812 5516 8818 5528
rect 9217 5525 9229 5528
rect 9263 5556 9275 5559
rect 9306 5556 9312 5568
rect 9263 5528 9312 5556
rect 9263 5525 9275 5528
rect 9217 5519 9275 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4488 5324 4629 5352
rect 4488 5312 4494 5324
rect 4617 5321 4629 5324
rect 4663 5321 4675 5355
rect 6178 5352 6184 5364
rect 6139 5324 6184 5352
rect 4617 5315 4675 5321
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7745 5355 7803 5361
rect 7745 5352 7757 5355
rect 7248 5324 7757 5352
rect 7248 5312 7254 5324
rect 7745 5321 7757 5324
rect 7791 5321 7803 5355
rect 9674 5352 9680 5364
rect 9635 5324 9680 5352
rect 7745 5315 7803 5321
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 4062 5244 4068 5296
rect 4120 5244 4126 5296
rect 4338 5244 4344 5296
rect 4396 5284 4402 5296
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 4396 5256 6561 5284
rect 4396 5244 4402 5256
rect 6549 5253 6561 5256
rect 6595 5284 6607 5287
rect 6822 5284 6828 5296
rect 6595 5256 6828 5284
rect 6595 5253 6607 5256
rect 6549 5247 6607 5253
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5216 3571 5219
rect 4080 5216 4108 5244
rect 8754 5216 8760 5228
rect 3559 5188 4108 5216
rect 8715 5188 8760 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3896 5157 3924 5188
rect 8754 5176 8760 5188
rect 8812 5176 8818 5228
rect 3881 5151 3939 5157
rect 3881 5117 3893 5151
rect 3927 5117 3939 5151
rect 3881 5111 3939 5117
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 4065 5151 4123 5157
rect 4065 5148 4077 5151
rect 4028 5120 4077 5148
rect 4028 5108 4034 5120
rect 4065 5117 4077 5120
rect 4111 5117 4123 5151
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 4065 5111 4123 5117
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 6880 5120 7389 5148
rect 6880 5108 6886 5120
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 9858 5108 9864 5160
rect 9916 5157 9922 5160
rect 9916 5151 9954 5157
rect 9942 5148 9954 5151
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 9942 5120 10333 5148
rect 9942 5117 9954 5120
rect 9916 5111 9954 5117
rect 10321 5117 10333 5120
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 9916 5108 9922 5111
rect 4341 5083 4399 5089
rect 4341 5049 4353 5083
rect 4387 5080 4399 5083
rect 4706 5080 4712 5092
rect 4387 5052 4712 5080
rect 4387 5049 4399 5052
rect 4341 5043 4399 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 5258 5080 5264 5092
rect 5219 5052 5264 5080
rect 5258 5040 5264 5052
rect 5316 5040 5322 5092
rect 5353 5083 5411 5089
rect 5353 5049 5365 5083
rect 5399 5080 5411 5083
rect 5442 5080 5448 5092
rect 5399 5052 5448 5080
rect 5399 5049 5411 5052
rect 5353 5043 5411 5049
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5368 5012 5396 5043
rect 5442 5040 5448 5052
rect 5500 5040 5506 5092
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6086 5080 6092 5092
rect 5951 5052 6092 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 6086 5040 6092 5052
rect 6144 5040 6150 5092
rect 8386 5080 8392 5092
rect 8347 5052 8392 5080
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5049 8539 5083
rect 8481 5043 8539 5049
rect 7006 5012 7012 5024
rect 5123 4984 5396 5012
rect 6967 4984 7012 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 8202 5012 8208 5024
rect 8163 4984 8208 5012
rect 8202 4972 8208 4984
rect 8260 5012 8266 5024
rect 8496 5012 8524 5043
rect 8260 4984 8524 5012
rect 8260 4972 8266 4984
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 9999 5015 10057 5021
rect 9999 5012 10011 5015
rect 9824 4984 10011 5012
rect 9824 4972 9830 4984
rect 9999 4981 10011 4984
rect 10045 4981 10057 5015
rect 9999 4975 10057 4981
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 3697 4811 3755 4817
rect 3697 4777 3709 4811
rect 3743 4808 3755 4811
rect 3970 4808 3976 4820
rect 3743 4780 3976 4808
rect 3743 4777 3755 4780
rect 3697 4771 3755 4777
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 4338 4808 4344 4820
rect 4299 4780 4344 4808
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 5905 4811 5963 4817
rect 5905 4808 5917 4811
rect 5316 4780 5917 4808
rect 5316 4768 5322 4780
rect 5905 4777 5917 4780
rect 5951 4777 5963 4811
rect 7098 4808 7104 4820
rect 7059 4780 7104 4808
rect 5905 4771 5963 4777
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 8202 4808 8208 4820
rect 8163 4780 8208 4808
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 5071 4743 5129 4749
rect 5071 4709 5083 4743
rect 5117 4740 5129 4743
rect 5350 4740 5356 4752
rect 5117 4712 5356 4740
rect 5117 4709 5129 4712
rect 5071 4703 5129 4709
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 7374 4700 7380 4752
rect 7432 4740 7438 4752
rect 7606 4743 7664 4749
rect 7606 4740 7618 4743
rect 7432 4712 7618 4740
rect 7432 4700 7438 4712
rect 7606 4709 7618 4712
rect 7652 4709 7664 4743
rect 7606 4703 7664 4709
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 2996 4675 3054 4681
rect 2996 4672 3008 4675
rect 2832 4644 3008 4672
rect 2832 4632 2838 4644
rect 2996 4641 3008 4644
rect 3042 4641 3054 4675
rect 7282 4672 7288 4684
rect 7243 4644 7288 4672
rect 2996 4635 3054 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 9728 4675 9786 4681
rect 9728 4641 9740 4675
rect 9774 4672 9786 4675
rect 10318 4672 10324 4684
rect 9774 4644 10324 4672
rect 9774 4641 9786 4644
rect 9728 4635 9786 4641
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 10686 4632 10692 4684
rect 10744 4681 10750 4684
rect 10744 4675 10782 4681
rect 10770 4641 10782 4675
rect 10744 4635 10782 4641
rect 10744 4632 10750 4635
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8444 4576 8585 4604
rect 8444 4564 8450 4576
rect 8573 4573 8585 4576
rect 8619 4604 8631 4607
rect 9815 4607 9873 4613
rect 9815 4604 9827 4607
rect 8619 4576 9827 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9815 4573 9827 4576
rect 9861 4573 9873 4607
rect 9815 4567 9873 4573
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 8904 4508 8953 4536
rect 8904 4496 8910 4508
rect 8941 4505 8953 4508
rect 8987 4536 8999 4539
rect 10827 4539 10885 4545
rect 10827 4536 10839 4539
rect 8987 4508 10839 4536
rect 8987 4505 8999 4508
rect 8941 4499 8999 4505
rect 10827 4505 10839 4508
rect 10873 4505 10885 4539
rect 10827 4499 10885 4505
rect 2590 4428 2596 4480
rect 2648 4468 2654 4480
rect 3099 4471 3157 4477
rect 3099 4468 3111 4471
rect 2648 4440 3111 4468
rect 2648 4428 2654 4440
rect 3099 4437 3111 4440
rect 3145 4437 3157 4471
rect 5626 4468 5632 4480
rect 5587 4440 5632 4468
rect 3099 4431 3157 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 6086 4428 6092 4480
rect 6144 4468 6150 4480
rect 6273 4471 6331 4477
rect 6273 4468 6285 4471
rect 6144 4440 6285 4468
rect 6144 4428 6150 4440
rect 6273 4437 6285 4440
rect 6319 4437 6331 4471
rect 6273 4431 6331 4437
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 3418 4264 3424 4276
rect 2832 4236 3424 4264
rect 2832 4224 2838 4236
rect 3418 4224 3424 4236
rect 3476 4224 3482 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 4801 4267 4859 4273
rect 4801 4264 4813 4267
rect 4488 4236 4813 4264
rect 4488 4224 4494 4236
rect 4801 4233 4813 4236
rect 4847 4264 4859 4267
rect 5350 4264 5356 4276
rect 4847 4236 5356 4264
rect 4847 4233 4859 4236
rect 4801 4227 4859 4233
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 8202 4224 8208 4276
rect 8260 4264 8266 4276
rect 8665 4267 8723 4273
rect 8665 4264 8677 4267
rect 8260 4236 8677 4264
rect 8260 4224 8266 4236
rect 8665 4233 8677 4236
rect 8711 4233 8723 4267
rect 8665 4227 8723 4233
rect 9953 4267 10011 4273
rect 9953 4233 9965 4267
rect 9999 4264 10011 4267
rect 10318 4264 10324 4276
rect 9999 4236 10324 4264
rect 9999 4233 10011 4236
rect 9953 4227 10011 4233
rect 3145 4199 3203 4205
rect 3145 4196 3157 4199
rect 2659 4168 3157 4196
rect 1648 4063 1706 4069
rect 1648 4029 1660 4063
rect 1694 4060 1706 4063
rect 1694 4032 2176 4060
rect 1694 4029 1706 4032
rect 1648 4023 1706 4029
rect 2148 3936 2176 4032
rect 2222 4020 2228 4072
rect 2280 4060 2286 4072
rect 2659 4069 2687 4168
rect 3145 4165 3157 4168
rect 3191 4196 3203 4199
rect 3234 4196 3240 4208
rect 3191 4168 3240 4196
rect 3191 4165 3203 4168
rect 3145 4159 3203 4165
rect 3234 4156 3240 4168
rect 3292 4156 3298 4208
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 7282 4196 7288 4208
rect 4764 4168 5488 4196
rect 4764 4156 4770 4168
rect 2731 4131 2789 4137
rect 2731 4097 2743 4131
rect 2777 4128 2789 4131
rect 5258 4128 5264 4140
rect 2777 4100 5264 4128
rect 2777 4097 2789 4100
rect 2731 4091 2789 4097
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5460 4128 5488 4168
rect 6932 4168 7288 4196
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 5460 4100 6193 4128
rect 6181 4097 6193 4100
rect 6227 4097 6239 4131
rect 6181 4091 6239 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6932 4128 6960 4168
rect 7282 4156 7288 4168
rect 7340 4156 7346 4208
rect 7098 4128 7104 4140
rect 6687 4100 6960 4128
rect 7059 4100 7104 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 2644 4063 2702 4069
rect 2644 4060 2656 4063
rect 2280 4032 2656 4060
rect 2280 4020 2286 4032
rect 2644 4029 2656 4032
rect 2690 4029 2702 4063
rect 2644 4023 2702 4029
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3992 2559 3995
rect 3694 3992 3700 4004
rect 2547 3964 3700 3992
rect 2547 3961 2559 3964
rect 2501 3955 2559 3961
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 3786 3952 3792 4004
rect 3844 3992 3850 4004
rect 4338 3992 4344 4004
rect 3844 3964 3889 3992
rect 4251 3964 4344 3992
rect 3844 3952 3850 3964
rect 4338 3952 4344 3964
rect 4396 3992 4402 4004
rect 5353 3995 5411 4001
rect 4396 3964 4844 3992
rect 4396 3952 4402 3964
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1719 3927 1777 3933
rect 1719 3924 1731 3927
rect 1452 3896 1731 3924
rect 1452 3884 1458 3896
rect 1719 3893 1731 3896
rect 1765 3893 1777 3927
rect 2130 3924 2136 3936
rect 2091 3896 2136 3924
rect 1719 3887 1777 3893
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 4816 3924 4844 3964
rect 5353 3961 5365 3995
rect 5399 3992 5411 3995
rect 5442 3992 5448 4004
rect 5399 3964 5448 3992
rect 5399 3961 5411 3964
rect 5353 3955 5411 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 5902 3992 5908 4004
rect 5863 3964 5908 3992
rect 5902 3952 5908 3964
rect 5960 3992 5966 4004
rect 6178 3992 6184 4004
rect 5960 3964 6184 3992
rect 5960 3952 5966 3964
rect 6178 3952 6184 3964
rect 6236 3952 6242 4004
rect 7374 3952 7380 4004
rect 7432 4001 7438 4004
rect 7432 3995 7480 4001
rect 7432 3961 7434 3995
rect 7468 3961 7480 3995
rect 8680 3992 8708 4227
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 10686 4224 10692 4276
rect 10744 4264 10750 4276
rect 10965 4267 11023 4273
rect 10965 4264 10977 4267
rect 10744 4236 10977 4264
rect 10744 4224 10750 4236
rect 10965 4233 10977 4236
rect 11011 4233 11023 4267
rect 10965 4227 11023 4233
rect 8846 4156 8852 4208
rect 8904 4156 8910 4208
rect 8864 4128 8892 4156
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8864 4100 8953 4128
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 9214 4128 9220 4140
rect 9175 4100 9220 4128
rect 8941 4091 8999 4097
rect 9214 4088 9220 4100
rect 9272 4128 9278 4140
rect 9582 4128 9588 4140
rect 9272 4100 9588 4128
rect 9272 4088 9278 4100
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 10318 4020 10324 4072
rect 10376 4060 10382 4072
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10376 4032 10425 4060
rect 10376 4020 10382 4032
rect 10413 4029 10425 4032
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 9033 3995 9091 4001
rect 9033 3992 9045 3995
rect 8680 3964 9045 3992
rect 7432 3955 7480 3961
rect 9033 3961 9045 3964
rect 9079 3961 9091 3995
rect 11054 3992 11060 4004
rect 9033 3955 9091 3961
rect 10612 3964 11060 3992
rect 7432 3952 7438 3955
rect 5534 3924 5540 3936
rect 4816 3896 5540 3924
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8202 3924 8208 3936
rect 8067 3896 8208 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 10612 3933 10640 3964
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 10597 3927 10655 3933
rect 10597 3893 10609 3927
rect 10643 3893 10655 3927
rect 10597 3887 10655 3893
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 3697 3723 3755 3729
rect 3697 3689 3709 3723
rect 3743 3720 3755 3723
rect 3786 3720 3792 3732
rect 3743 3692 3792 3720
rect 3743 3689 3755 3692
rect 3697 3683 3755 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 5258 3680 5264 3732
rect 5316 3720 5322 3732
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 5316 3692 5641 3720
rect 5316 3680 5322 3692
rect 5629 3689 5641 3692
rect 5675 3689 5687 3723
rect 5629 3683 5687 3689
rect 7193 3723 7251 3729
rect 7193 3689 7205 3723
rect 7239 3720 7251 3723
rect 7374 3720 7380 3732
rect 7239 3692 7380 3720
rect 7239 3689 7251 3692
rect 7193 3683 7251 3689
rect 7374 3680 7380 3692
rect 7432 3720 7438 3732
rect 7469 3723 7527 3729
rect 7469 3720 7481 3723
rect 7432 3692 7481 3720
rect 7432 3680 7438 3692
rect 7469 3689 7481 3692
rect 7515 3689 7527 3723
rect 7469 3683 7527 3689
rect 7929 3723 7987 3729
rect 7929 3689 7941 3723
rect 7975 3720 7987 3723
rect 8018 3720 8024 3732
rect 7975 3692 8024 3720
rect 7975 3689 7987 3692
rect 7929 3683 7987 3689
rect 8018 3680 8024 3692
rect 8076 3720 8082 3732
rect 10919 3723 10977 3729
rect 10919 3720 10931 3723
rect 8076 3692 10931 3720
rect 8076 3680 8082 3692
rect 10919 3689 10931 3692
rect 10965 3689 10977 3723
rect 10919 3683 10977 3689
rect 1857 3655 1915 3661
rect 1857 3621 1869 3655
rect 1903 3652 1915 3655
rect 2590 3652 2596 3664
rect 1903 3624 2596 3652
rect 1903 3621 1915 3624
rect 1857 3615 1915 3621
rect 2590 3612 2596 3624
rect 2648 3612 2654 3664
rect 4430 3661 4436 3664
rect 4427 3652 4436 3661
rect 4391 3624 4436 3652
rect 4427 3615 4436 3624
rect 4430 3612 4436 3615
rect 4488 3612 4494 3664
rect 5353 3655 5411 3661
rect 5353 3621 5365 3655
rect 5399 3652 5411 3655
rect 5442 3652 5448 3664
rect 5399 3624 5448 3652
rect 5399 3621 5411 3624
rect 5353 3615 5411 3621
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 5994 3652 6000 3664
rect 5955 3624 6000 3652
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 8202 3652 8208 3664
rect 8163 3624 8208 3652
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 8757 3655 8815 3661
rect 8757 3621 8769 3655
rect 8803 3652 8815 3655
rect 9214 3652 9220 3664
rect 8803 3624 9220 3652
rect 8803 3621 8815 3624
rect 8757 3615 8815 3621
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 2000 3587 2058 3593
rect 2000 3553 2012 3587
rect 2046 3584 2058 3587
rect 2314 3584 2320 3596
rect 2046 3556 2320 3584
rect 2046 3553 2058 3556
rect 2000 3547 2058 3553
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3200 3556 4077 3584
rect 3200 3544 3206 3556
rect 4065 3553 4077 3556
rect 4111 3584 4123 3587
rect 5258 3584 5264 3596
rect 4111 3556 5264 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3584 9738 3596
rect 10134 3584 10140 3596
rect 9732 3556 10140 3584
rect 9732 3544 9738 3556
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10848 3587 10906 3593
rect 10848 3553 10860 3587
rect 10894 3584 10906 3587
rect 11330 3584 11336 3596
rect 10894 3556 11336 3584
rect 10894 3553 10906 3556
rect 10848 3547 10906 3553
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 2087 3519 2145 3525
rect 2087 3485 2099 3519
rect 2133 3516 2145 3519
rect 2498 3516 2504 3528
rect 2133 3488 2504 3516
rect 2133 3485 2145 3488
rect 2087 3479 2145 3485
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 2682 3476 2688 3528
rect 2740 3516 2746 3528
rect 2961 3519 3019 3525
rect 2961 3516 2973 3519
rect 2740 3488 2973 3516
rect 2740 3476 2746 3488
rect 2961 3485 2973 3488
rect 3007 3485 3019 3519
rect 5902 3516 5908 3528
rect 5863 3488 5908 3516
rect 2961 3479 3019 3485
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 6178 3516 6184 3528
rect 6139 3488 6184 3516
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 9582 3516 9588 3528
rect 8159 3488 9588 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 2685 3383 2743 3389
rect 2685 3349 2697 3383
rect 2731 3380 2743 3383
rect 2774 3380 2780 3392
rect 2731 3352 2780 3380
rect 2731 3349 2743 3352
rect 2685 3343 2743 3349
rect 2774 3340 2780 3352
rect 2832 3340 2838 3392
rect 4246 3340 4252 3392
rect 4304 3380 4310 3392
rect 4985 3383 5043 3389
rect 4985 3380 4997 3383
rect 4304 3352 4997 3380
rect 4304 3340 4310 3352
rect 4985 3349 4997 3352
rect 5031 3349 5043 3383
rect 4985 3343 5043 3349
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 9364 3352 9873 3380
rect 9364 3340 9370 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 9861 3343 9919 3349
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 2409 3179 2467 3185
rect 2409 3176 2421 3179
rect 2372 3148 2421 3176
rect 2372 3136 2378 3148
rect 2409 3145 2421 3148
rect 2455 3145 2467 3179
rect 2409 3139 2467 3145
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 5353 3179 5411 3185
rect 5353 3176 5365 3179
rect 5316 3148 5365 3176
rect 5316 3136 5322 3148
rect 5353 3145 5365 3148
rect 5399 3145 5411 3179
rect 5353 3139 5411 3145
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 5994 3176 6000 3188
rect 5951 3148 6000 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 8021 3179 8079 3185
rect 8021 3145 8033 3179
rect 8067 3176 8079 3179
rect 8202 3176 8208 3188
rect 8067 3148 8208 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9217 3179 9275 3185
rect 9217 3145 9229 3179
rect 9263 3176 9275 3179
rect 9582 3176 9588 3188
rect 9263 3148 9588 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 10229 3179 10287 3185
rect 10229 3176 10241 3179
rect 10192 3148 10241 3176
rect 10192 3136 10198 3148
rect 10229 3145 10241 3148
rect 10275 3145 10287 3179
rect 10229 3139 10287 3145
rect 11330 3136 11336 3188
rect 11388 3176 11394 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 11388 3148 11621 3176
rect 11388 3136 11394 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 11609 3139 11667 3145
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 8754 3108 8760 3120
rect 2648 3080 2728 3108
rect 8715 3080 8760 3108
rect 2648 3068 2654 3080
rect 2700 3049 2728 3080
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3009 2743 3043
rect 3326 3040 3332 3052
rect 3287 3012 3332 3040
rect 2685 3003 2743 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 4154 3040 4160 3052
rect 4115 3012 4160 3040
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 5960 3012 6193 3040
rect 5960 3000 5966 3012
rect 6181 3009 6193 3012
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 8076 3012 8217 3040
rect 8076 3000 8082 3012
rect 8205 3009 8217 3012
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3040 9643 3043
rect 9858 3040 9864 3052
rect 9631 3012 9864 3040
rect 9631 3009 9643 3012
rect 9585 3003 9643 3009
rect 1210 2932 1216 2984
rect 1268 2972 1274 2984
rect 1670 2981 1676 2984
rect 1648 2975 1676 2981
rect 1648 2972 1660 2975
rect 1268 2944 1660 2972
rect 1268 2932 1274 2944
rect 1648 2941 1660 2944
rect 1728 2972 1734 2984
rect 2041 2975 2099 2981
rect 2041 2972 2053 2975
rect 1728 2944 2053 2972
rect 1648 2935 1676 2941
rect 1670 2932 1676 2935
rect 1728 2932 1734 2944
rect 2041 2941 2053 2944
rect 2087 2941 2099 2975
rect 3510 2972 3516 2984
rect 2041 2935 2099 2941
rect 3344 2944 3516 2972
rect 2774 2864 2780 2916
rect 2832 2904 2838 2916
rect 2832 2876 2925 2904
rect 2832 2864 2838 2876
rect 3050 2864 3056 2916
rect 3108 2904 3114 2916
rect 3344 2904 3372 2944
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3697 2975 3755 2981
rect 3697 2941 3709 2975
rect 3743 2972 3755 2975
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 3743 2944 4077 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 4065 2941 4077 2944
rect 4111 2972 4123 2975
rect 6822 2972 6828 2984
rect 4111 2944 4476 2972
rect 6735 2944 6828 2972
rect 4111 2941 4123 2944
rect 4065 2935 4123 2941
rect 4448 2916 4476 2944
rect 6822 2932 6828 2944
rect 6880 2972 6886 2984
rect 9692 2981 9720 3012
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 6880 2944 7389 2972
rect 6880 2932 6886 2944
rect 7377 2941 7389 2944
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 9723 2944 9757 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 10778 2932 10784 2984
rect 10836 2981 10842 2984
rect 10836 2975 10874 2981
rect 10862 2972 10874 2975
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 10862 2944 11253 2972
rect 10862 2941 10874 2944
rect 10836 2935 10874 2941
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 10836 2932 10842 2935
rect 3108 2876 3372 2904
rect 3436 2876 4384 2904
rect 3108 2864 3114 2876
rect 1719 2839 1777 2845
rect 1719 2805 1731 2839
rect 1765 2836 1777 2839
rect 2314 2836 2320 2848
rect 1765 2808 2320 2836
rect 1765 2805 1777 2808
rect 1719 2799 1777 2805
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 2792 2836 2820 2864
rect 3436 2836 3464 2876
rect 4356 2848 4384 2876
rect 4430 2864 4436 2916
rect 4488 2913 4494 2916
rect 4488 2907 4536 2913
rect 4488 2873 4490 2907
rect 4524 2873 4536 2907
rect 4488 2867 4536 2873
rect 4488 2864 4494 2867
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 8352 2876 8397 2904
rect 8352 2864 8358 2876
rect 2792 2808 3464 2836
rect 4338 2796 4344 2848
rect 4396 2836 4402 2848
rect 5077 2839 5135 2845
rect 5077 2836 5089 2839
rect 4396 2808 5089 2836
rect 4396 2796 4402 2808
rect 5077 2805 5089 2808
rect 5123 2805 5135 2839
rect 7006 2836 7012 2848
rect 6967 2808 7012 2836
rect 5077 2799 5135 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 9861 2839 9919 2845
rect 9861 2805 9873 2839
rect 9907 2836 9919 2839
rect 10134 2836 10140 2848
rect 9907 2808 10140 2836
rect 9907 2805 9919 2808
rect 9861 2799 9919 2805
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 10318 2796 10324 2848
rect 10376 2836 10382 2848
rect 10919 2839 10977 2845
rect 10919 2836 10931 2839
rect 10376 2808 10931 2836
rect 10376 2796 10382 2808
rect 10919 2805 10931 2808
rect 10965 2805 10977 2839
rect 10919 2799 10977 2805
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 1535 2635 1593 2641
rect 1535 2601 1547 2635
rect 1581 2632 1593 2635
rect 2406 2632 2412 2644
rect 1581 2604 2412 2632
rect 1581 2601 1593 2604
rect 1535 2595 1593 2601
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 2866 2632 2872 2644
rect 2516 2604 2872 2632
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 2516 2564 2544 2604
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4249 2635 4307 2641
rect 4249 2632 4261 2635
rect 4212 2604 4261 2632
rect 4212 2592 4218 2604
rect 4249 2601 4261 2604
rect 4295 2601 4307 2635
rect 4249 2595 4307 2601
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 4709 2635 4767 2641
rect 4709 2632 4721 2635
rect 4396 2604 4721 2632
rect 4396 2592 4402 2604
rect 4709 2601 4721 2604
rect 4755 2632 4767 2635
rect 4755 2604 5120 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 1995 2536 2544 2564
rect 2593 2567 2651 2573
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 2593 2533 2605 2567
rect 2639 2564 2651 2567
rect 3513 2567 3571 2573
rect 3513 2564 3525 2567
rect 2639 2536 3525 2564
rect 2639 2533 2651 2536
rect 2593 2527 2651 2533
rect 3513 2533 3525 2536
rect 3559 2564 3571 2567
rect 4062 2564 4068 2576
rect 3559 2536 4068 2564
rect 3559 2533 3571 2536
rect 3513 2527 3571 2533
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 1964 2496 1992 2527
rect 4062 2524 4068 2536
rect 4120 2524 4126 2576
rect 4982 2564 4988 2576
rect 4943 2536 4988 2564
rect 4982 2524 4988 2536
rect 5040 2524 5046 2576
rect 5092 2573 5120 2604
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 6052 2604 6653 2632
rect 6052 2592 6058 2604
rect 6641 2601 6653 2604
rect 6687 2632 6699 2635
rect 8113 2635 8171 2641
rect 6687 2604 7144 2632
rect 6687 2601 6699 2604
rect 6641 2595 6699 2601
rect 5077 2567 5135 2573
rect 5077 2533 5089 2567
rect 5123 2533 5135 2567
rect 5077 2527 5135 2533
rect 5629 2567 5687 2573
rect 5629 2533 5641 2567
rect 5675 2564 5687 2567
rect 6178 2564 6184 2576
rect 5675 2536 6184 2564
rect 5675 2533 5687 2536
rect 5629 2527 5687 2533
rect 6178 2524 6184 2536
rect 6236 2524 6242 2576
rect 6365 2567 6423 2573
rect 6365 2533 6377 2567
rect 6411 2564 6423 2567
rect 7006 2564 7012 2576
rect 6411 2536 7012 2564
rect 6411 2533 6423 2536
rect 6365 2527 6423 2533
rect 7006 2524 7012 2536
rect 7064 2524 7070 2576
rect 7116 2573 7144 2604
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 8202 2632 8208 2644
rect 8159 2604 8208 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9490 2632 9496 2644
rect 9171 2604 9496 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2533 7159 2567
rect 7101 2527 7159 2533
rect 1510 2468 1992 2496
rect 8481 2499 8539 2505
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 9140 2496 9168 2595
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 12066 2632 12072 2644
rect 12027 2604 12072 2632
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 8527 2468 9168 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 10226 2456 10232 2508
rect 10284 2496 10290 2508
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 10284 2468 10333 2496
rect 10284 2456 10290 2468
rect 10321 2465 10333 2468
rect 10367 2496 10379 2499
rect 10873 2499 10931 2505
rect 10873 2496 10885 2499
rect 10367 2468 10885 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 10873 2465 10885 2468
rect 10919 2465 10931 2499
rect 10873 2459 10931 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 12084 2496 12112 2592
rect 13170 2496 13176 2508
rect 11471 2468 12112 2496
rect 13131 2468 13176 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 13170 2456 13176 2468
rect 13228 2496 13234 2508
rect 13725 2499 13783 2505
rect 13725 2496 13737 2499
rect 13228 2468 13737 2496
rect 13228 2456 13234 2468
rect 13725 2465 13737 2468
rect 13771 2465 13783 2499
rect 13725 2459 13783 2465
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2363 2400 2513 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2501 2397 2513 2400
rect 2547 2428 2559 2431
rect 2682 2428 2688 2440
rect 2547 2400 2688 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 2958 2428 2964 2440
rect 2919 2400 2964 2428
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5040 2400 5917 2428
rect 5040 2388 5046 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 7282 2428 7288 2440
rect 7243 2400 7288 2428
rect 5905 2391 5963 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 10505 2363 10563 2369
rect 10505 2329 10517 2363
rect 10551 2360 10563 2363
rect 11882 2360 11888 2372
rect 10551 2332 11888 2360
rect 10551 2329 10563 2332
rect 10505 2323 10563 2329
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 13357 2363 13415 2369
rect 13357 2329 13369 2363
rect 13403 2360 13415 2363
rect 14182 2360 14188 2372
rect 13403 2332 14188 2360
rect 13403 2329 13415 2332
rect 13357 2323 13415 2329
rect 14182 2320 14188 2332
rect 14240 2320 14246 2372
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8444 2264 8677 2292
rect 8444 2252 8450 2264
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 8665 2255 8723 2261
rect 11609 2295 11667 2301
rect 11609 2261 11621 2295
rect 11655 2292 11667 2295
rect 12342 2292 12348 2304
rect 11655 2264 12348 2292
rect 11655 2261 11667 2264
rect 11609 2255 11667 2261
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 3878 1980 3884 2032
rect 3936 2020 3942 2032
rect 4614 2020 4620 2032
rect 3936 1992 4620 2020
rect 3936 1980 3942 1992
rect 4614 1980 4620 1992
rect 4672 1980 4678 2032
rect 5166 552 5172 604
rect 5224 592 5230 604
rect 5718 592 5724 604
rect 5224 564 5724 592
rect 5224 552 5230 564
rect 5718 552 5724 564
rect 5776 552 5782 604
<< via1 >>
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 4068 37272 4120 37324
rect 6000 37272 6052 37324
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 9956 36524 10008 36576
rect 10692 36524 10744 36576
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 9312 36320 9364 36372
rect 8576 36252 8628 36304
rect 7472 36227 7524 36236
rect 7472 36193 7516 36227
rect 7516 36193 7524 36227
rect 7472 36184 7524 36193
rect 9588 36184 9640 36236
rect 9772 36227 9824 36236
rect 9772 36193 9790 36227
rect 9790 36193 9824 36227
rect 9772 36184 9824 36193
rect 8300 36048 8352 36100
rect 10324 35980 10376 36032
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 7472 35776 7524 35828
rect 9588 35776 9640 35828
rect 7012 35751 7064 35760
rect 7012 35717 7021 35751
rect 7021 35717 7055 35751
rect 7055 35717 7064 35751
rect 7012 35708 7064 35717
rect 8760 35683 8812 35692
rect 8760 35649 8769 35683
rect 8769 35649 8803 35683
rect 8803 35649 8812 35683
rect 8760 35640 8812 35649
rect 10324 35683 10376 35692
rect 10324 35649 10333 35683
rect 10333 35649 10367 35683
rect 10367 35649 10376 35683
rect 10324 35640 10376 35649
rect 10784 35683 10836 35692
rect 10784 35649 10793 35683
rect 10793 35649 10827 35683
rect 10827 35649 10836 35683
rect 10784 35640 10836 35649
rect 5632 35572 5684 35624
rect 8300 35547 8352 35556
rect 8300 35513 8309 35547
rect 8309 35513 8343 35547
rect 8343 35513 8352 35547
rect 8300 35504 8352 35513
rect 8576 35504 8628 35556
rect 10416 35547 10468 35556
rect 10416 35513 10425 35547
rect 10425 35513 10459 35547
rect 10459 35513 10468 35547
rect 10416 35504 10468 35513
rect 9772 35479 9824 35488
rect 9772 35445 9781 35479
rect 9781 35445 9815 35479
rect 9815 35445 9824 35479
rect 9772 35436 9824 35445
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 6000 35232 6052 35284
rect 8300 35232 8352 35284
rect 9956 35232 10008 35284
rect 13176 35275 13228 35284
rect 13176 35241 13185 35275
rect 13185 35241 13219 35275
rect 13219 35241 13228 35275
rect 13176 35232 13228 35241
rect 8576 35164 8628 35216
rect 10600 35207 10652 35216
rect 10600 35173 10609 35207
rect 10609 35173 10643 35207
rect 10643 35173 10652 35207
rect 10600 35164 10652 35173
rect 6736 35096 6788 35148
rect 7288 35096 7340 35148
rect 12072 35139 12124 35148
rect 12072 35105 12090 35139
rect 12090 35105 12124 35139
rect 12072 35096 12124 35105
rect 13084 35096 13136 35148
rect 8116 35071 8168 35080
rect 8116 35037 8125 35071
rect 8125 35037 8159 35071
rect 8159 35037 8168 35071
rect 8116 35028 8168 35037
rect 8208 34960 8260 35012
rect 7564 34935 7616 34944
rect 7564 34901 7573 34935
rect 7573 34901 7607 34935
rect 7607 34901 7616 34935
rect 7564 34892 7616 34901
rect 8024 34892 8076 34944
rect 10968 35028 11020 35080
rect 11520 35028 11572 35080
rect 12532 34892 12584 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 8116 34688 8168 34740
rect 10140 34688 10192 34740
rect 11060 34688 11112 34740
rect 5816 34663 5868 34672
rect 5816 34629 5825 34663
rect 5825 34629 5859 34663
rect 5859 34629 5868 34663
rect 5816 34620 5868 34629
rect 7564 34620 7616 34672
rect 8024 34595 8076 34604
rect 8024 34561 8033 34595
rect 8033 34561 8067 34595
rect 8067 34561 8076 34595
rect 8024 34552 8076 34561
rect 9956 34552 10008 34604
rect 10784 34595 10836 34604
rect 10784 34561 10793 34595
rect 10793 34561 10827 34595
rect 10827 34561 10836 34595
rect 10784 34552 10836 34561
rect 5540 34484 5592 34536
rect 6736 34484 6788 34536
rect 8668 34527 8720 34536
rect 8668 34493 8677 34527
rect 8677 34493 8711 34527
rect 8711 34493 8720 34527
rect 8668 34484 8720 34493
rect 8852 34484 8904 34536
rect 12072 34527 12124 34536
rect 12072 34493 12081 34527
rect 12081 34493 12115 34527
rect 12115 34493 12124 34527
rect 12072 34484 12124 34493
rect 12440 34527 12492 34536
rect 12440 34493 12449 34527
rect 12449 34493 12483 34527
rect 12483 34493 12492 34527
rect 12440 34484 12492 34493
rect 13084 34484 13136 34536
rect 7932 34416 7984 34468
rect 7288 34348 7340 34400
rect 10232 34348 10284 34400
rect 10600 34348 10652 34400
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 5356 34144 5408 34196
rect 13176 34187 13228 34196
rect 13176 34153 13185 34187
rect 13185 34153 13219 34187
rect 13219 34153 13228 34187
rect 13176 34144 13228 34153
rect 6368 34119 6420 34128
rect 6368 34085 6377 34119
rect 6377 34085 6411 34119
rect 6411 34085 6420 34119
rect 6368 34076 6420 34085
rect 7932 34119 7984 34128
rect 7932 34085 7941 34119
rect 7941 34085 7975 34119
rect 7975 34085 7984 34119
rect 7932 34076 7984 34085
rect 10048 34119 10100 34128
rect 10048 34085 10051 34119
rect 10051 34085 10085 34119
rect 10085 34085 10100 34119
rect 10048 34076 10100 34085
rect 5264 34051 5316 34060
rect 5264 34017 5282 34051
rect 5282 34017 5316 34051
rect 5264 34008 5316 34017
rect 11060 34076 11112 34128
rect 12164 34008 12216 34060
rect 13452 34008 13504 34060
rect 6184 33872 6236 33924
rect 8300 33940 8352 33992
rect 8760 33940 8812 33992
rect 9496 33940 9548 33992
rect 9680 33983 9732 33992
rect 9680 33949 9689 33983
rect 9689 33949 9723 33983
rect 9723 33949 9732 33983
rect 9680 33940 9732 33949
rect 11336 33940 11388 33992
rect 10784 33872 10836 33924
rect 7564 33847 7616 33856
rect 7564 33813 7573 33847
rect 7573 33813 7607 33847
rect 7607 33813 7616 33847
rect 7564 33804 7616 33813
rect 10968 33847 11020 33856
rect 10968 33813 10977 33847
rect 10977 33813 11011 33847
rect 11011 33813 11020 33847
rect 10968 33804 11020 33813
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 4896 33600 4948 33652
rect 6368 33600 6420 33652
rect 10232 33643 10284 33652
rect 10232 33609 10241 33643
rect 10241 33609 10275 33643
rect 10275 33609 10284 33643
rect 10232 33600 10284 33609
rect 11980 33600 12032 33652
rect 13452 33643 13504 33652
rect 13452 33609 13461 33643
rect 13461 33609 13495 33643
rect 13495 33609 13504 33643
rect 13452 33600 13504 33609
rect 7564 33507 7616 33516
rect 7564 33473 7573 33507
rect 7573 33473 7607 33507
rect 7607 33473 7616 33507
rect 7564 33464 7616 33473
rect 8024 33507 8076 33516
rect 8024 33473 8033 33507
rect 8033 33473 8067 33507
rect 8067 33473 8076 33507
rect 8024 33464 8076 33473
rect 9680 33464 9732 33516
rect 12532 33507 12584 33516
rect 12532 33473 12541 33507
rect 12541 33473 12575 33507
rect 12575 33473 12584 33507
rect 12532 33464 12584 33473
rect 12808 33507 12860 33516
rect 12808 33473 12817 33507
rect 12817 33473 12851 33507
rect 12851 33473 12860 33507
rect 12808 33464 12860 33473
rect 4712 33439 4764 33448
rect 4712 33405 4756 33439
rect 4756 33405 4764 33439
rect 5264 33439 5316 33448
rect 4712 33396 4764 33405
rect 5264 33405 5273 33439
rect 5273 33405 5307 33439
rect 5307 33405 5316 33439
rect 5264 33396 5316 33405
rect 9312 33439 9364 33448
rect 6092 33328 6144 33380
rect 9312 33405 9321 33439
rect 9321 33405 9355 33439
rect 9355 33405 9364 33439
rect 9312 33396 9364 33405
rect 11152 33396 11204 33448
rect 12256 33396 12308 33448
rect 7656 33371 7708 33380
rect 7656 33337 7665 33371
rect 7665 33337 7699 33371
rect 7699 33337 7708 33371
rect 7656 33328 7708 33337
rect 7288 33260 7340 33312
rect 9404 33260 9456 33312
rect 10876 33328 10928 33380
rect 10048 33260 10100 33312
rect 11060 33260 11112 33312
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 6184 33099 6236 33108
rect 6184 33065 6193 33099
rect 6193 33065 6227 33099
rect 6227 33065 6236 33099
rect 6184 33056 6236 33065
rect 7656 33099 7708 33108
rect 7656 33065 7665 33099
rect 7665 33065 7699 33099
rect 7699 33065 7708 33099
rect 7656 33056 7708 33065
rect 7932 33099 7984 33108
rect 7932 33065 7941 33099
rect 7941 33065 7975 33099
rect 7975 33065 7984 33099
rect 7932 33056 7984 33065
rect 8300 33099 8352 33108
rect 8300 33065 8309 33099
rect 8309 33065 8343 33099
rect 8343 33065 8352 33099
rect 8300 33056 8352 33065
rect 10416 33056 10468 33108
rect 10876 33056 10928 33108
rect 12532 33099 12584 33108
rect 12532 33065 12541 33099
rect 12541 33065 12575 33099
rect 12575 33065 12584 33099
rect 12532 33056 12584 33065
rect 7196 32988 7248 33040
rect 9404 32988 9456 33040
rect 11060 32988 11112 33040
rect 11704 32988 11756 33040
rect 6000 32920 6052 32972
rect 8576 32963 8628 32972
rect 8576 32929 8594 32963
rect 8594 32929 8628 32963
rect 8576 32920 8628 32929
rect 13084 32963 13136 32972
rect 13084 32929 13102 32963
rect 13102 32929 13136 32963
rect 13084 32920 13136 32929
rect 7472 32852 7524 32904
rect 10416 32852 10468 32904
rect 11520 32895 11572 32904
rect 11520 32861 11529 32895
rect 11529 32861 11563 32895
rect 11563 32861 11572 32895
rect 11520 32852 11572 32861
rect 11612 32852 11664 32904
rect 8760 32716 8812 32768
rect 9312 32759 9364 32768
rect 9312 32725 9321 32759
rect 9321 32725 9355 32759
rect 9355 32725 9364 32759
rect 9312 32716 9364 32725
rect 11336 32759 11388 32768
rect 11336 32725 11345 32759
rect 11345 32725 11379 32759
rect 11379 32725 11388 32759
rect 11336 32716 11388 32725
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 7932 32512 7984 32564
rect 8576 32512 8628 32564
rect 8668 32512 8720 32564
rect 11704 32555 11756 32564
rect 11704 32521 11713 32555
rect 11713 32521 11747 32555
rect 11747 32521 11756 32555
rect 11704 32512 11756 32521
rect 12440 32512 12492 32564
rect 8944 32444 8996 32496
rect 8760 32376 8812 32428
rect 6828 32351 6880 32360
rect 6828 32317 6837 32351
rect 6837 32317 6871 32351
rect 6871 32317 6880 32351
rect 6828 32308 6880 32317
rect 10692 32308 10744 32360
rect 7196 32283 7248 32292
rect 6000 32172 6052 32224
rect 7196 32249 7199 32283
rect 7199 32249 7233 32283
rect 7233 32249 7248 32283
rect 7196 32240 7248 32249
rect 9404 32240 9456 32292
rect 10232 32283 10284 32292
rect 10232 32249 10241 32283
rect 10241 32249 10275 32283
rect 10275 32249 10284 32283
rect 10232 32240 10284 32249
rect 10416 32215 10468 32224
rect 10416 32181 10425 32215
rect 10425 32181 10459 32215
rect 10459 32181 10468 32215
rect 10416 32172 10468 32181
rect 12164 32215 12216 32224
rect 12164 32181 12173 32215
rect 12173 32181 12207 32215
rect 12207 32181 12216 32215
rect 12164 32172 12216 32181
rect 13084 32215 13136 32224
rect 13084 32181 13093 32215
rect 13093 32181 13127 32215
rect 13127 32181 13136 32215
rect 13084 32172 13136 32181
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 9680 31968 9732 32020
rect 11520 31968 11572 32020
rect 6828 31943 6880 31952
rect 6828 31909 6837 31943
rect 6837 31909 6871 31943
rect 6871 31909 6880 31943
rect 6828 31900 6880 31909
rect 8760 31900 8812 31952
rect 10692 31943 10744 31952
rect 10692 31909 10701 31943
rect 10701 31909 10735 31943
rect 10735 31909 10744 31943
rect 10692 31900 10744 31909
rect 5816 31832 5868 31884
rect 6644 31875 6696 31884
rect 6644 31841 6653 31875
rect 6653 31841 6687 31875
rect 6687 31841 6696 31875
rect 6644 31832 6696 31841
rect 8116 31875 8168 31884
rect 7748 31764 7800 31816
rect 8116 31841 8125 31875
rect 8125 31841 8159 31875
rect 8159 31841 8168 31875
rect 8116 31832 8168 31841
rect 10232 31875 10284 31884
rect 10232 31841 10241 31875
rect 10241 31841 10275 31875
rect 10275 31841 10284 31875
rect 10232 31832 10284 31841
rect 11244 31875 11296 31884
rect 11244 31841 11288 31875
rect 11288 31841 11296 31875
rect 11244 31832 11296 31841
rect 10140 31764 10192 31816
rect 7380 31628 7432 31680
rect 8668 31671 8720 31680
rect 8668 31637 8677 31671
rect 8677 31637 8711 31671
rect 8711 31637 8720 31671
rect 8668 31628 8720 31637
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 5816 31467 5868 31476
rect 5816 31433 5825 31467
rect 5825 31433 5859 31467
rect 5859 31433 5868 31467
rect 5816 31424 5868 31433
rect 7380 31331 7432 31340
rect 7380 31297 7389 31331
rect 7389 31297 7423 31331
rect 7423 31297 7432 31331
rect 7380 31288 7432 31297
rect 9312 31331 9364 31340
rect 9312 31297 9321 31331
rect 9321 31297 9355 31331
rect 9355 31297 9364 31331
rect 9312 31288 9364 31297
rect 6920 31263 6972 31272
rect 6920 31229 6929 31263
rect 6929 31229 6963 31263
rect 6963 31229 6972 31263
rect 6920 31220 6972 31229
rect 6644 31127 6696 31136
rect 6644 31093 6653 31127
rect 6653 31093 6687 31127
rect 6687 31093 6696 31127
rect 8300 31220 8352 31272
rect 8668 31263 8720 31272
rect 8668 31229 8677 31263
rect 8677 31229 8711 31263
rect 8711 31229 8720 31263
rect 8668 31220 8720 31229
rect 10232 31424 10284 31476
rect 10784 31288 10836 31340
rect 10140 31263 10192 31272
rect 10140 31229 10149 31263
rect 10149 31229 10183 31263
rect 10183 31229 10192 31263
rect 10140 31220 10192 31229
rect 10968 31152 11020 31204
rect 12164 31152 12216 31204
rect 6644 31084 6696 31093
rect 8116 31084 8168 31136
rect 8668 31084 8720 31136
rect 11244 31084 11296 31136
rect 11520 31084 11572 31136
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 7748 30923 7800 30932
rect 7748 30889 7757 30923
rect 7757 30889 7791 30923
rect 7791 30889 7800 30923
rect 7748 30880 7800 30889
rect 9496 30923 9548 30932
rect 9496 30889 9505 30923
rect 9505 30889 9539 30923
rect 9539 30889 9548 30923
rect 10784 30923 10836 30932
rect 9496 30880 9548 30889
rect 8208 30855 8260 30864
rect 8208 30821 8217 30855
rect 8217 30821 8251 30855
rect 8251 30821 8260 30855
rect 8208 30812 8260 30821
rect 10784 30889 10793 30923
rect 10793 30889 10827 30923
rect 10827 30889 10836 30923
rect 10784 30880 10836 30889
rect 9864 30855 9916 30864
rect 9864 30821 9873 30855
rect 9873 30821 9907 30855
rect 9907 30821 9916 30855
rect 11428 30855 11480 30864
rect 9864 30812 9916 30821
rect 11428 30821 11437 30855
rect 11437 30821 11471 30855
rect 11471 30821 11480 30855
rect 11428 30812 11480 30821
rect 7012 30719 7064 30728
rect 7012 30685 7021 30719
rect 7021 30685 7055 30719
rect 7055 30685 7064 30719
rect 7012 30676 7064 30685
rect 7932 30676 7984 30728
rect 8392 30719 8444 30728
rect 8392 30685 8401 30719
rect 8401 30685 8435 30719
rect 8435 30685 8444 30719
rect 8392 30676 8444 30685
rect 11336 30719 11388 30728
rect 11336 30685 11345 30719
rect 11345 30685 11379 30719
rect 11379 30685 11388 30719
rect 11336 30676 11388 30685
rect 12164 30676 12216 30728
rect 6920 30583 6972 30592
rect 6920 30549 6929 30583
rect 6929 30549 6963 30583
rect 6963 30549 6972 30583
rect 6920 30540 6972 30549
rect 8392 30540 8444 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 8484 30268 8536 30320
rect 11428 30336 11480 30388
rect 11336 30200 11388 30252
rect 7472 30175 7524 30184
rect 7472 30141 7481 30175
rect 7481 30141 7515 30175
rect 7515 30141 7524 30175
rect 7472 30132 7524 30141
rect 8760 30175 8812 30184
rect 8760 30141 8769 30175
rect 8769 30141 8803 30175
rect 8803 30141 8812 30175
rect 8760 30132 8812 30141
rect 9956 30132 10008 30184
rect 6644 29996 6696 30048
rect 9772 30064 9824 30116
rect 7564 30039 7616 30048
rect 7564 30005 7573 30039
rect 7573 30005 7607 30039
rect 7607 30005 7616 30039
rect 7564 29996 7616 30005
rect 8300 30039 8352 30048
rect 8300 30005 8309 30039
rect 8309 30005 8343 30039
rect 8343 30005 8352 30039
rect 8300 29996 8352 30005
rect 9312 30039 9364 30048
rect 9312 30005 9321 30039
rect 9321 30005 9355 30039
rect 9355 30005 9364 30039
rect 9312 29996 9364 30005
rect 9404 29996 9456 30048
rect 10416 30064 10468 30116
rect 11060 30064 11112 30116
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 7472 29835 7524 29844
rect 7472 29801 7481 29835
rect 7481 29801 7515 29835
rect 7515 29801 7524 29835
rect 7472 29792 7524 29801
rect 7932 29835 7984 29844
rect 7932 29801 7941 29835
rect 7941 29801 7975 29835
rect 7975 29801 7984 29835
rect 7932 29792 7984 29801
rect 10968 29835 11020 29844
rect 10968 29801 10977 29835
rect 10977 29801 11011 29835
rect 11011 29801 11020 29835
rect 10968 29792 11020 29801
rect 8392 29724 8444 29776
rect 10416 29767 10468 29776
rect 10416 29733 10419 29767
rect 10419 29733 10453 29767
rect 10453 29733 10468 29767
rect 10416 29724 10468 29733
rect 11980 29767 12032 29776
rect 11980 29733 11989 29767
rect 11989 29733 12023 29767
rect 12023 29733 12032 29767
rect 11980 29724 12032 29733
rect 6644 29656 6696 29708
rect 8208 29699 8260 29708
rect 8208 29665 8217 29699
rect 8217 29665 8251 29699
rect 8251 29665 8260 29699
rect 8208 29656 8260 29665
rect 8668 29656 8720 29708
rect 6736 29588 6788 29640
rect 7196 29631 7248 29640
rect 7196 29597 7205 29631
rect 7205 29597 7239 29631
rect 7239 29597 7248 29631
rect 7196 29588 7248 29597
rect 8852 29588 8904 29640
rect 10692 29588 10744 29640
rect 11888 29631 11940 29640
rect 11888 29597 11897 29631
rect 11897 29597 11931 29631
rect 11931 29597 11940 29631
rect 11888 29588 11940 29597
rect 12164 29631 12216 29640
rect 12164 29597 12173 29631
rect 12173 29597 12207 29631
rect 12207 29597 12216 29631
rect 12164 29588 12216 29597
rect 5356 29452 5408 29504
rect 9956 29495 10008 29504
rect 9956 29461 9965 29495
rect 9965 29461 9999 29495
rect 9999 29461 10008 29495
rect 9956 29452 10008 29461
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 8300 29291 8352 29300
rect 8300 29257 8309 29291
rect 8309 29257 8343 29291
rect 8343 29257 8352 29291
rect 8300 29248 8352 29257
rect 8668 29291 8720 29300
rect 8668 29257 8677 29291
rect 8677 29257 8711 29291
rect 8711 29257 8720 29291
rect 8668 29248 8720 29257
rect 10416 29291 10468 29300
rect 8576 29180 8628 29232
rect 5264 29155 5316 29164
rect 5264 29121 5273 29155
rect 5273 29121 5307 29155
rect 5307 29121 5316 29155
rect 5264 29112 5316 29121
rect 5908 29155 5960 29164
rect 5908 29121 5917 29155
rect 5917 29121 5951 29155
rect 5951 29121 5960 29155
rect 5908 29112 5960 29121
rect 7196 29112 7248 29164
rect 8852 29112 8904 29164
rect 6644 29044 6696 29096
rect 7932 29044 7984 29096
rect 8576 29044 8628 29096
rect 4896 28976 4948 29028
rect 4988 28976 5040 29028
rect 5356 29019 5408 29028
rect 5356 28985 5365 29019
rect 5365 28985 5399 29019
rect 5399 28985 5408 29019
rect 5356 28976 5408 28985
rect 8116 28976 8168 29028
rect 10416 29257 10425 29291
rect 10425 29257 10459 29291
rect 10459 29257 10468 29291
rect 10416 29248 10468 29257
rect 11888 29291 11940 29300
rect 11888 29257 11897 29291
rect 11897 29257 11931 29291
rect 11931 29257 11940 29291
rect 11888 29248 11940 29257
rect 11980 29044 12032 29096
rect 9680 28976 9732 29028
rect 10324 28976 10376 29028
rect 10692 28951 10744 28960
rect 10692 28917 10701 28951
rect 10701 28917 10735 28951
rect 10735 28917 10744 28951
rect 10692 28908 10744 28917
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 7196 28704 7248 28756
rect 9312 28704 9364 28756
rect 9956 28747 10008 28756
rect 9956 28713 9965 28747
rect 9965 28713 9999 28747
rect 9999 28713 10008 28747
rect 9956 28704 10008 28713
rect 8116 28636 8168 28688
rect 8668 28636 8720 28688
rect 4896 28611 4948 28620
rect 4896 28577 4914 28611
rect 4914 28577 4948 28611
rect 4896 28568 4948 28577
rect 6368 28611 6420 28620
rect 6368 28577 6377 28611
rect 6377 28577 6411 28611
rect 6411 28577 6420 28611
rect 6368 28568 6420 28577
rect 6644 28611 6696 28620
rect 6644 28577 6653 28611
rect 6653 28577 6687 28611
rect 6687 28577 6696 28611
rect 6644 28568 6696 28577
rect 7564 28568 7616 28620
rect 8300 28568 8352 28620
rect 11244 28611 11296 28620
rect 6828 28543 6880 28552
rect 6828 28509 6837 28543
rect 6837 28509 6871 28543
rect 6871 28509 6880 28543
rect 6828 28500 6880 28509
rect 8392 28500 8444 28552
rect 11244 28577 11253 28611
rect 11253 28577 11287 28611
rect 11287 28577 11296 28611
rect 11244 28568 11296 28577
rect 10416 28500 10468 28552
rect 4804 28364 4856 28416
rect 5264 28407 5316 28416
rect 5264 28373 5273 28407
rect 5273 28373 5307 28407
rect 5307 28373 5316 28407
rect 5264 28364 5316 28373
rect 5356 28364 5408 28416
rect 6736 28364 6788 28416
rect 9404 28364 9456 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 6644 28160 6696 28212
rect 7564 28160 7616 28212
rect 8668 28160 8720 28212
rect 3240 27956 3292 28008
rect 5632 28092 5684 28144
rect 7748 28135 7800 28144
rect 7748 28101 7757 28135
rect 7757 28101 7791 28135
rect 7791 28101 7800 28135
rect 7748 28092 7800 28101
rect 8116 28135 8168 28144
rect 8116 28101 8125 28135
rect 8125 28101 8159 28135
rect 8159 28101 8168 28135
rect 8116 28092 8168 28101
rect 5356 28024 5408 28076
rect 6828 28067 6880 28076
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 8392 28024 8444 28076
rect 9404 27999 9456 28008
rect 9404 27965 9413 27999
rect 9413 27965 9447 27999
rect 9447 27965 9456 27999
rect 9404 27956 9456 27965
rect 11060 28203 11112 28212
rect 11060 28169 11069 28203
rect 11069 28169 11103 28203
rect 11103 28169 11112 28203
rect 11060 28160 11112 28169
rect 10692 28024 10744 28076
rect 10140 27956 10192 28008
rect 5264 27888 5316 27940
rect 5724 27931 5776 27940
rect 5724 27897 5733 27931
rect 5733 27897 5767 27931
rect 5767 27897 5776 27931
rect 5724 27888 5776 27897
rect 7932 27888 7984 27940
rect 8116 27888 8168 27940
rect 4068 27820 4120 27872
rect 4896 27863 4948 27872
rect 4896 27829 4905 27863
rect 4905 27829 4939 27863
rect 4939 27829 4948 27863
rect 4896 27820 4948 27829
rect 10324 27820 10376 27872
rect 11244 27820 11296 27872
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 4804 27659 4856 27668
rect 4804 27625 4813 27659
rect 4813 27625 4847 27659
rect 4847 27625 4856 27659
rect 4804 27616 4856 27625
rect 5264 27616 5316 27668
rect 6184 27616 6236 27668
rect 6828 27616 6880 27668
rect 5356 27548 5408 27600
rect 5632 27548 5684 27600
rect 6276 27548 6328 27600
rect 7104 27548 7156 27600
rect 7380 27548 7432 27600
rect 9864 27591 9916 27600
rect 9864 27557 9873 27591
rect 9873 27557 9907 27591
rect 9907 27557 9916 27591
rect 9864 27548 9916 27557
rect 11980 27548 12032 27600
rect 4528 27480 4580 27532
rect 8392 27523 8444 27532
rect 8392 27489 8436 27523
rect 8436 27489 8444 27523
rect 8392 27480 8444 27489
rect 12808 27523 12860 27532
rect 12808 27489 12852 27523
rect 12852 27489 12860 27523
rect 12808 27480 12860 27489
rect 5356 27455 5408 27464
rect 5356 27421 5365 27455
rect 5365 27421 5399 27455
rect 5399 27421 5408 27455
rect 5356 27412 5408 27421
rect 5724 27455 5776 27464
rect 5724 27421 5733 27455
rect 5733 27421 5767 27455
rect 5767 27421 5776 27455
rect 5724 27412 5776 27421
rect 7840 27412 7892 27464
rect 9772 27455 9824 27464
rect 9772 27421 9781 27455
rect 9781 27421 9815 27455
rect 9815 27421 9824 27455
rect 9772 27412 9824 27421
rect 10232 27412 10284 27464
rect 11520 27412 11572 27464
rect 12072 27412 12124 27464
rect 7012 27344 7064 27396
rect 6000 27276 6052 27328
rect 6644 27276 6696 27328
rect 8852 27276 8904 27328
rect 9404 27319 9456 27328
rect 9404 27285 9413 27319
rect 9413 27285 9447 27319
rect 9447 27285 9456 27319
rect 9404 27276 9456 27285
rect 12532 27276 12584 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 5356 27072 5408 27124
rect 6276 27115 6328 27124
rect 6276 27081 6285 27115
rect 6285 27081 6319 27115
rect 6319 27081 6328 27115
rect 6276 27072 6328 27081
rect 7840 27115 7892 27124
rect 7840 27081 7849 27115
rect 7849 27081 7883 27115
rect 7883 27081 7892 27115
rect 7840 27072 7892 27081
rect 11980 27115 12032 27124
rect 11980 27081 11989 27115
rect 11989 27081 12023 27115
rect 12023 27081 12032 27115
rect 11980 27072 12032 27081
rect 12808 27072 12860 27124
rect 13636 27072 13688 27124
rect 4528 27047 4580 27056
rect 4528 27013 4537 27047
rect 4537 27013 4571 27047
rect 4571 27013 4580 27047
rect 4528 27004 4580 27013
rect 5540 27004 5592 27056
rect 8392 27004 8444 27056
rect 10232 27047 10284 27056
rect 10232 27013 10241 27047
rect 10241 27013 10275 27047
rect 10275 27013 10284 27047
rect 10232 27004 10284 27013
rect 2872 26868 2924 26920
rect 4804 26936 4856 26988
rect 6920 26979 6972 26988
rect 6920 26945 6929 26979
rect 6929 26945 6963 26979
rect 6963 26945 6972 26979
rect 6920 26936 6972 26945
rect 7012 26936 7064 26988
rect 9864 26936 9916 26988
rect 11336 26936 11388 26988
rect 4160 26911 4212 26920
rect 4160 26877 4178 26911
rect 4178 26877 4212 26911
rect 4160 26868 4212 26877
rect 4436 26732 4488 26784
rect 6184 26868 6236 26920
rect 5264 26843 5316 26852
rect 5264 26809 5273 26843
rect 5273 26809 5307 26843
rect 5307 26809 5316 26843
rect 5264 26800 5316 26809
rect 5172 26732 5224 26784
rect 8300 26868 8352 26920
rect 11060 26868 11112 26920
rect 12256 26868 12308 26920
rect 9680 26843 9732 26852
rect 9680 26809 9689 26843
rect 9689 26809 9723 26843
rect 9723 26809 9732 26843
rect 9680 26800 9732 26809
rect 9772 26843 9824 26852
rect 9772 26809 9781 26843
rect 9781 26809 9815 26843
rect 9815 26809 9824 26843
rect 9772 26800 9824 26809
rect 12072 26800 12124 26852
rect 11060 26732 11112 26784
rect 11980 26732 12032 26784
rect 12716 26732 12768 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 5632 26571 5684 26580
rect 5632 26537 5641 26571
rect 5641 26537 5675 26571
rect 5675 26537 5684 26571
rect 5632 26528 5684 26537
rect 6920 26528 6972 26580
rect 9680 26528 9732 26580
rect 11520 26528 11572 26580
rect 12624 26528 12676 26580
rect 12900 26571 12952 26580
rect 12900 26537 12909 26571
rect 12909 26537 12943 26571
rect 12943 26537 12952 26571
rect 12900 26528 12952 26537
rect 4620 26460 4672 26512
rect 5356 26460 5408 26512
rect 6184 26460 6236 26512
rect 9588 26460 9640 26512
rect 9864 26503 9916 26512
rect 9864 26469 9873 26503
rect 9873 26469 9907 26503
rect 9907 26469 9916 26503
rect 9864 26460 9916 26469
rect 11336 26503 11388 26512
rect 11336 26469 11345 26503
rect 11345 26469 11379 26503
rect 11379 26469 11388 26503
rect 11336 26460 11388 26469
rect 12440 26503 12492 26512
rect 12440 26469 12449 26503
rect 12449 26469 12483 26503
rect 12483 26469 12492 26503
rect 12440 26460 12492 26469
rect 4436 26392 4488 26444
rect 5448 26324 5500 26376
rect 7564 26392 7616 26444
rect 8300 26435 8352 26444
rect 8300 26401 8309 26435
rect 8309 26401 8343 26435
rect 8343 26401 8352 26435
rect 8300 26392 8352 26401
rect 13360 26460 13412 26512
rect 6460 26324 6512 26376
rect 8392 26367 8444 26376
rect 8392 26333 8401 26367
rect 8401 26333 8435 26367
rect 8435 26333 8444 26367
rect 8392 26324 8444 26333
rect 9956 26324 10008 26376
rect 11060 26324 11112 26376
rect 11152 26324 11204 26376
rect 11980 26324 12032 26376
rect 12808 26324 12860 26376
rect 5632 26256 5684 26308
rect 7656 26188 7708 26240
rect 10048 26188 10100 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 5264 25984 5316 26036
rect 6460 26027 6512 26036
rect 6460 25993 6469 26027
rect 6469 25993 6503 26027
rect 6503 25993 6512 26027
rect 6460 25984 6512 25993
rect 8300 25984 8352 26036
rect 9312 25984 9364 26036
rect 9496 25984 9548 26036
rect 9864 25984 9916 26036
rect 11336 25984 11388 26036
rect 6920 25916 6972 25968
rect 7932 25916 7984 25968
rect 8392 25848 8444 25900
rect 7656 25780 7708 25832
rect 4620 25755 4672 25764
rect 4620 25721 4623 25755
rect 4623 25721 4657 25755
rect 4657 25721 4672 25755
rect 4620 25712 4672 25721
rect 12532 25891 12584 25900
rect 10048 25823 10100 25832
rect 10048 25789 10057 25823
rect 10057 25789 10091 25823
rect 10091 25789 10100 25823
rect 10048 25780 10100 25789
rect 12532 25857 12541 25891
rect 12541 25857 12575 25891
rect 12575 25857 12584 25891
rect 12532 25848 12584 25857
rect 12624 25848 12676 25900
rect 10968 25780 11020 25832
rect 10508 25712 10560 25764
rect 3976 25644 4028 25696
rect 5540 25687 5592 25696
rect 5540 25653 5549 25687
rect 5549 25653 5583 25687
rect 5583 25653 5592 25687
rect 5540 25644 5592 25653
rect 6092 25687 6144 25696
rect 6092 25653 6101 25687
rect 6101 25653 6135 25687
rect 6135 25653 6144 25687
rect 6092 25644 6144 25653
rect 7564 25644 7616 25696
rect 11980 25644 12032 25696
rect 12440 25644 12492 25696
rect 13360 25644 13412 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 6092 25440 6144 25492
rect 8392 25483 8444 25492
rect 8392 25449 8401 25483
rect 8401 25449 8435 25483
rect 8435 25449 8444 25483
rect 8392 25440 8444 25449
rect 8852 25440 8904 25492
rect 9956 25483 10008 25492
rect 9956 25449 9965 25483
rect 9965 25449 9999 25483
rect 9999 25449 10008 25483
rect 9956 25440 10008 25449
rect 10968 25483 11020 25492
rect 10968 25449 10977 25483
rect 10977 25449 11011 25483
rect 11011 25449 11020 25483
rect 10968 25440 11020 25449
rect 11980 25440 12032 25492
rect 12440 25440 12492 25492
rect 12532 25440 12584 25492
rect 13268 25440 13320 25492
rect 3148 25415 3200 25424
rect 3148 25381 3157 25415
rect 3157 25381 3191 25415
rect 3191 25381 3200 25415
rect 3148 25372 3200 25381
rect 4620 25372 4672 25424
rect 5264 25415 5316 25424
rect 5264 25381 5267 25415
rect 5267 25381 5301 25415
rect 5301 25381 5316 25415
rect 5264 25372 5316 25381
rect 7104 25415 7156 25424
rect 7104 25381 7107 25415
rect 7107 25381 7141 25415
rect 7141 25381 7156 25415
rect 7104 25372 7156 25381
rect 7932 25372 7984 25424
rect 10508 25372 10560 25424
rect 11796 25372 11848 25424
rect 2688 25347 2740 25356
rect 2688 25313 2697 25347
rect 2697 25313 2731 25347
rect 2731 25313 2740 25347
rect 2688 25304 2740 25313
rect 2964 25347 3016 25356
rect 2964 25313 2973 25347
rect 2973 25313 3007 25347
rect 3007 25313 3016 25347
rect 2964 25304 3016 25313
rect 10140 25304 10192 25356
rect 12716 25347 12768 25356
rect 12716 25313 12725 25347
rect 12725 25313 12759 25347
rect 12759 25313 12768 25347
rect 12716 25304 12768 25313
rect 13452 25304 13504 25356
rect 4160 25168 4212 25220
rect 5908 25100 5960 25152
rect 8484 25279 8536 25288
rect 8484 25245 8493 25279
rect 8493 25245 8527 25279
rect 8527 25245 8536 25279
rect 8484 25236 8536 25245
rect 11980 25236 12032 25288
rect 7288 25100 7340 25152
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 2688 24896 2740 24948
rect 2964 24896 3016 24948
rect 5908 24803 5960 24812
rect 5908 24769 5917 24803
rect 5917 24769 5951 24803
rect 5951 24769 5960 24803
rect 5908 24760 5960 24769
rect 6000 24760 6052 24812
rect 7012 24760 7064 24812
rect 8484 24896 8536 24948
rect 10048 24939 10100 24948
rect 10048 24905 10057 24939
rect 10057 24905 10091 24939
rect 10091 24905 10100 24939
rect 10048 24896 10100 24905
rect 8852 24803 8904 24812
rect 8852 24769 8861 24803
rect 8861 24769 8895 24803
rect 8895 24769 8904 24803
rect 8852 24760 8904 24769
rect 9496 24803 9548 24812
rect 9496 24769 9505 24803
rect 9505 24769 9539 24803
rect 9539 24769 9548 24803
rect 9496 24760 9548 24769
rect 3056 24556 3108 24608
rect 4252 24692 4304 24744
rect 5540 24692 5592 24744
rect 7288 24667 7340 24676
rect 7288 24633 7297 24667
rect 7297 24633 7331 24667
rect 7331 24633 7340 24667
rect 7288 24624 7340 24633
rect 7656 24624 7708 24676
rect 9312 24624 9364 24676
rect 10508 24896 10560 24948
rect 11796 24939 11848 24948
rect 11796 24905 11805 24939
rect 11805 24905 11839 24939
rect 11839 24905 11848 24939
rect 11796 24896 11848 24905
rect 13452 24896 13504 24948
rect 10784 24760 10836 24812
rect 12532 24828 12584 24880
rect 13360 24828 13412 24880
rect 10968 24692 11020 24744
rect 12532 24735 12584 24744
rect 12532 24701 12541 24735
rect 12541 24701 12575 24735
rect 12575 24701 12584 24735
rect 12532 24692 12584 24701
rect 12900 24735 12952 24744
rect 12900 24701 12909 24735
rect 12909 24701 12943 24735
rect 12943 24701 12952 24735
rect 12900 24692 12952 24701
rect 3976 24556 4028 24608
rect 5264 24556 5316 24608
rect 6644 24599 6696 24608
rect 6644 24565 6653 24599
rect 6653 24565 6687 24599
rect 6687 24565 6696 24599
rect 6644 24556 6696 24565
rect 7104 24556 7156 24608
rect 11244 24556 11296 24608
rect 12532 24599 12584 24608
rect 12532 24565 12541 24599
rect 12541 24565 12575 24599
rect 12575 24565 12584 24599
rect 12532 24556 12584 24565
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 8760 24395 8812 24404
rect 8760 24361 8769 24395
rect 8769 24361 8803 24395
rect 8803 24361 8812 24395
rect 8760 24352 8812 24361
rect 10140 24352 10192 24404
rect 12900 24352 12952 24404
rect 5448 24284 5500 24336
rect 7288 24284 7340 24336
rect 10416 24284 10468 24336
rect 10968 24327 11020 24336
rect 10968 24293 10977 24327
rect 10977 24293 11011 24327
rect 11011 24293 11020 24327
rect 10968 24284 11020 24293
rect 11244 24327 11296 24336
rect 11244 24293 11253 24327
rect 11253 24293 11287 24327
rect 11287 24293 11296 24327
rect 11244 24284 11296 24293
rect 12992 24284 13044 24336
rect 3148 24216 3200 24268
rect 4252 24216 4304 24268
rect 6276 24216 6328 24268
rect 8392 24216 8444 24268
rect 9680 24259 9732 24268
rect 9680 24225 9689 24259
rect 9689 24225 9723 24259
rect 9723 24225 9732 24259
rect 9680 24216 9732 24225
rect 12624 24259 12676 24268
rect 12624 24225 12668 24259
rect 12668 24225 12676 24259
rect 12624 24216 12676 24225
rect 4712 24148 4764 24200
rect 7932 24148 7984 24200
rect 11152 24191 11204 24200
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 11520 24191 11572 24200
rect 11520 24157 11529 24191
rect 11529 24157 11563 24191
rect 11563 24157 11572 24191
rect 11520 24148 11572 24157
rect 12072 24148 12124 24200
rect 5448 24080 5500 24132
rect 7656 24123 7708 24132
rect 7656 24089 7665 24123
rect 7665 24089 7699 24123
rect 7699 24089 7708 24123
rect 7656 24080 7708 24089
rect 8668 24080 8720 24132
rect 9864 24123 9916 24132
rect 9864 24089 9873 24123
rect 9873 24089 9907 24123
rect 9907 24089 9916 24123
rect 9864 24080 9916 24089
rect 3056 24012 3108 24064
rect 4252 24012 4304 24064
rect 5540 24055 5592 24064
rect 5540 24021 5549 24055
rect 5549 24021 5583 24055
rect 5583 24021 5592 24055
rect 5540 24012 5592 24021
rect 6828 24055 6880 24064
rect 6828 24021 6837 24055
rect 6837 24021 6871 24055
rect 6871 24021 6880 24055
rect 6828 24012 6880 24021
rect 10876 24012 10928 24064
rect 11980 24012 12032 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 3148 23808 3200 23860
rect 6644 23851 6696 23860
rect 6644 23817 6653 23851
rect 6653 23817 6687 23851
rect 6687 23817 6696 23851
rect 6644 23808 6696 23817
rect 11244 23851 11296 23860
rect 11244 23817 11253 23851
rect 11253 23817 11287 23851
rect 11287 23817 11296 23851
rect 11244 23808 11296 23817
rect 4712 23740 4764 23792
rect 11152 23740 11204 23792
rect 7656 23672 7708 23724
rect 10416 23672 10468 23724
rect 10876 23715 10928 23724
rect 10876 23681 10885 23715
rect 10885 23681 10919 23715
rect 10919 23681 10928 23715
rect 10876 23672 10928 23681
rect 3148 23536 3200 23588
rect 3332 23468 3384 23520
rect 4252 23604 4304 23656
rect 5080 23647 5132 23656
rect 5080 23613 5089 23647
rect 5089 23613 5123 23647
rect 5123 23613 5132 23647
rect 5448 23647 5500 23656
rect 5080 23604 5132 23613
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 5540 23604 5592 23656
rect 6276 23647 6328 23656
rect 6276 23613 6285 23647
rect 6285 23613 6319 23647
rect 6319 23613 6328 23647
rect 6276 23604 6328 23613
rect 6828 23647 6880 23656
rect 6828 23613 6837 23647
rect 6837 23613 6871 23647
rect 6871 23613 6880 23647
rect 6828 23604 6880 23613
rect 10232 23604 10284 23656
rect 12624 23647 12676 23656
rect 12624 23613 12633 23647
rect 12633 23613 12667 23647
rect 12667 23613 12676 23647
rect 12624 23604 12676 23613
rect 5908 23579 5960 23588
rect 5908 23545 5917 23579
rect 5917 23545 5951 23579
rect 5951 23545 5960 23579
rect 5908 23536 5960 23545
rect 6644 23536 6696 23588
rect 8668 23579 8720 23588
rect 4068 23468 4120 23520
rect 4712 23511 4764 23520
rect 4712 23477 4721 23511
rect 4721 23477 4755 23511
rect 4755 23477 4764 23511
rect 4712 23468 4764 23477
rect 5264 23468 5316 23520
rect 8392 23511 8444 23520
rect 8392 23477 8401 23511
rect 8401 23477 8435 23511
rect 8435 23477 8444 23511
rect 8392 23468 8444 23477
rect 8668 23545 8677 23579
rect 8677 23545 8711 23579
rect 8711 23545 8720 23579
rect 8668 23536 8720 23545
rect 9680 23579 9732 23588
rect 9680 23545 9689 23579
rect 9689 23545 9723 23579
rect 9723 23545 9732 23579
rect 9680 23536 9732 23545
rect 10416 23536 10468 23588
rect 11612 23536 11664 23588
rect 9864 23511 9916 23520
rect 9864 23477 9873 23511
rect 9873 23477 9907 23511
rect 9907 23477 9916 23511
rect 9864 23468 9916 23477
rect 10508 23468 10560 23520
rect 10784 23468 10836 23520
rect 12164 23468 12216 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 5908 23264 5960 23316
rect 7288 23307 7340 23316
rect 4988 23239 5040 23248
rect 4988 23205 4997 23239
rect 4997 23205 5031 23239
rect 5031 23205 5040 23239
rect 4988 23196 5040 23205
rect 2964 23171 3016 23180
rect 2964 23137 2973 23171
rect 2973 23137 3007 23171
rect 3007 23137 3016 23171
rect 2964 23128 3016 23137
rect 7288 23273 7297 23307
rect 7297 23273 7331 23307
rect 7331 23273 7340 23307
rect 7288 23264 7340 23273
rect 7932 23307 7984 23316
rect 7932 23273 7941 23307
rect 7941 23273 7975 23307
rect 7975 23273 7984 23307
rect 7932 23264 7984 23273
rect 8944 23307 8996 23316
rect 8944 23273 8953 23307
rect 8953 23273 8987 23307
rect 8987 23273 8996 23307
rect 8944 23264 8996 23273
rect 10232 23264 10284 23316
rect 6644 23196 6696 23248
rect 11428 23264 11480 23316
rect 11244 23239 11296 23248
rect 11244 23205 11253 23239
rect 11253 23205 11287 23239
rect 11287 23205 11296 23239
rect 11244 23196 11296 23205
rect 7012 23128 7064 23180
rect 8116 23171 8168 23180
rect 8116 23137 8125 23171
rect 8125 23137 8159 23171
rect 8159 23137 8168 23171
rect 8116 23128 8168 23137
rect 9680 23171 9732 23180
rect 9680 23137 9689 23171
rect 9689 23137 9723 23171
rect 9723 23137 9732 23171
rect 9680 23128 9732 23137
rect 3516 23060 3568 23112
rect 5632 23060 5684 23112
rect 11520 23103 11572 23112
rect 11520 23069 11529 23103
rect 11529 23069 11563 23103
rect 11563 23069 11572 23103
rect 11520 23060 11572 23069
rect 5448 23035 5500 23044
rect 5448 23001 5457 23035
rect 5457 23001 5491 23035
rect 5491 23001 5500 23035
rect 5448 22992 5500 23001
rect 3332 22924 3384 22976
rect 4252 22967 4304 22976
rect 4252 22933 4261 22967
rect 4261 22933 4295 22967
rect 4295 22933 4304 22967
rect 4252 22924 4304 22933
rect 4620 22967 4672 22976
rect 4620 22933 4629 22967
rect 4629 22933 4663 22967
rect 4663 22933 4672 22967
rect 4620 22924 4672 22933
rect 7380 22924 7432 22976
rect 8484 22924 8536 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2964 22763 3016 22772
rect 2964 22729 2973 22763
rect 2973 22729 3007 22763
rect 3007 22729 3016 22763
rect 2964 22720 3016 22729
rect 3516 22763 3568 22772
rect 3516 22729 3525 22763
rect 3525 22729 3559 22763
rect 3559 22729 3568 22763
rect 3516 22720 3568 22729
rect 4988 22720 5040 22772
rect 5448 22720 5500 22772
rect 4436 22652 4488 22704
rect 4620 22627 4672 22636
rect 4620 22593 4629 22627
rect 4629 22593 4663 22627
rect 4663 22593 4672 22627
rect 4620 22584 4672 22593
rect 4988 22584 5040 22636
rect 6644 22720 6696 22772
rect 8116 22763 8168 22772
rect 8116 22729 8125 22763
rect 8125 22729 8159 22763
rect 8159 22729 8168 22763
rect 8116 22720 8168 22729
rect 11428 22763 11480 22772
rect 11428 22729 11437 22763
rect 11437 22729 11471 22763
rect 11471 22729 11480 22763
rect 11428 22720 11480 22729
rect 12532 22720 12584 22772
rect 10600 22652 10652 22704
rect 7196 22627 7248 22636
rect 7196 22593 7205 22627
rect 7205 22593 7239 22627
rect 7239 22593 7248 22627
rect 7196 22584 7248 22593
rect 9864 22627 9916 22636
rect 9864 22593 9873 22627
rect 9873 22593 9907 22627
rect 9907 22593 9916 22627
rect 9864 22584 9916 22593
rect 10416 22627 10468 22636
rect 10416 22593 10425 22627
rect 10425 22593 10459 22627
rect 10459 22593 10468 22627
rect 10416 22584 10468 22593
rect 4344 22516 4396 22568
rect 8484 22559 8536 22568
rect 4988 22491 5040 22500
rect 4988 22457 4991 22491
rect 4991 22457 5025 22491
rect 5025 22457 5040 22491
rect 4988 22448 5040 22457
rect 8484 22525 8493 22559
rect 8493 22525 8527 22559
rect 8527 22525 8536 22559
rect 8484 22516 8536 22525
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 9680 22516 9732 22568
rect 10232 22559 10284 22568
rect 10232 22525 10241 22559
rect 10241 22525 10275 22559
rect 10275 22525 10284 22559
rect 10232 22516 10284 22525
rect 12532 22516 12584 22568
rect 13452 22559 13504 22568
rect 13452 22525 13461 22559
rect 13461 22525 13495 22559
rect 13495 22525 13504 22559
rect 13452 22516 13504 22525
rect 6920 22491 6972 22500
rect 6920 22457 6929 22491
rect 6929 22457 6963 22491
rect 6963 22457 6972 22491
rect 6920 22448 6972 22457
rect 7380 22448 7432 22500
rect 9128 22491 9180 22500
rect 9128 22457 9137 22491
rect 9137 22457 9171 22491
rect 9171 22457 9180 22491
rect 9128 22448 9180 22457
rect 10968 22423 11020 22432
rect 10968 22389 10977 22423
rect 10977 22389 11011 22423
rect 11011 22389 11020 22423
rect 10968 22380 11020 22389
rect 11060 22380 11112 22432
rect 11244 22380 11296 22432
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 5448 22219 5500 22228
rect 5448 22185 5457 22219
rect 5457 22185 5491 22219
rect 5491 22185 5500 22219
rect 5448 22176 5500 22185
rect 6828 22176 6880 22228
rect 6920 22176 6972 22228
rect 9128 22176 9180 22228
rect 4988 22108 5040 22160
rect 6000 22040 6052 22092
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 10048 22176 10100 22228
rect 10232 22176 10284 22228
rect 10968 22176 11020 22228
rect 12072 22176 12124 22228
rect 12532 22151 12584 22160
rect 4528 22015 4580 22024
rect 4528 21981 4537 22015
rect 4537 21981 4571 22015
rect 4571 21981 4580 22015
rect 4528 21972 4580 21981
rect 5540 21972 5592 22024
rect 6920 21972 6972 22024
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 12532 22117 12541 22151
rect 12541 22117 12575 22151
rect 12575 22117 12584 22151
rect 12532 22108 12584 22117
rect 11428 22040 11480 22092
rect 12072 22083 12124 22092
rect 12072 22049 12081 22083
rect 12081 22049 12115 22083
rect 12115 22049 12124 22083
rect 12072 22040 12124 22049
rect 9496 21972 9548 22024
rect 11152 21972 11204 22024
rect 10968 21947 11020 21956
rect 10968 21913 10977 21947
rect 10977 21913 11011 21947
rect 11011 21913 11020 21947
rect 10968 21904 11020 21913
rect 11888 21947 11940 21956
rect 11888 21913 11897 21947
rect 11897 21913 11931 21947
rect 11931 21913 11940 21947
rect 11888 21904 11940 21913
rect 4252 21836 4304 21888
rect 4620 21836 4672 21888
rect 9680 21836 9732 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 4988 21632 5040 21684
rect 5448 21632 5500 21684
rect 9496 21675 9548 21684
rect 6920 21607 6972 21616
rect 6920 21573 6929 21607
rect 6929 21573 6963 21607
rect 6963 21573 6972 21607
rect 6920 21564 6972 21573
rect 9496 21641 9505 21675
rect 9505 21641 9539 21675
rect 9539 21641 9548 21675
rect 9496 21632 9548 21641
rect 11152 21632 11204 21684
rect 8760 21564 8812 21616
rect 12624 21607 12676 21616
rect 12624 21573 12633 21607
rect 12633 21573 12667 21607
rect 12667 21573 12676 21607
rect 12624 21564 12676 21573
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 7564 21539 7616 21548
rect 7564 21505 7573 21539
rect 7573 21505 7607 21539
rect 7607 21505 7616 21539
rect 7564 21496 7616 21505
rect 9588 21496 9640 21548
rect 4620 21428 4672 21480
rect 6736 21428 6788 21480
rect 5080 21360 5132 21412
rect 8300 21428 8352 21480
rect 9680 21428 9732 21480
rect 3792 21335 3844 21344
rect 3792 21301 3801 21335
rect 3801 21301 3835 21335
rect 3835 21301 3844 21335
rect 3792 21292 3844 21301
rect 4344 21292 4396 21344
rect 4436 21292 4488 21344
rect 6000 21292 6052 21344
rect 8300 21335 8352 21344
rect 8300 21301 8309 21335
rect 8309 21301 8343 21335
rect 8343 21301 8352 21335
rect 8300 21292 8352 21301
rect 9772 21335 9824 21344
rect 9772 21301 9781 21335
rect 9781 21301 9815 21335
rect 9815 21301 9824 21335
rect 11520 21360 11572 21412
rect 11888 21360 11940 21412
rect 9772 21292 9824 21301
rect 11428 21292 11480 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 3792 21088 3844 21140
rect 4528 21088 4580 21140
rect 5632 21088 5684 21140
rect 6828 21088 6880 21140
rect 9496 21088 9548 21140
rect 10232 21088 10284 21140
rect 11152 21088 11204 21140
rect 12072 21088 12124 21140
rect 6644 21020 6696 21072
rect 10416 21020 10468 21072
rect 11980 21020 12032 21072
rect 4436 20995 4488 21004
rect 4436 20961 4445 20995
rect 4445 20961 4479 20995
rect 4479 20961 4488 20995
rect 4436 20952 4488 20961
rect 4620 20995 4672 21004
rect 4620 20961 4629 20995
rect 4629 20961 4663 20995
rect 4663 20961 4672 20995
rect 4620 20952 4672 20961
rect 7748 20952 7800 21004
rect 8576 20952 8628 21004
rect 3976 20884 4028 20936
rect 6276 20884 6328 20936
rect 7196 20859 7248 20868
rect 7196 20825 7205 20859
rect 7205 20825 7239 20859
rect 7239 20825 7248 20859
rect 7196 20816 7248 20825
rect 7380 20816 7432 20868
rect 6920 20748 6972 20800
rect 9680 20748 9732 20800
rect 9772 20748 9824 20800
rect 11152 20952 11204 21004
rect 11612 20952 11664 21004
rect 11520 20816 11572 20868
rect 12072 20816 12124 20868
rect 11612 20748 11664 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 6276 20587 6328 20596
rect 6276 20553 6285 20587
rect 6285 20553 6319 20587
rect 6319 20553 6328 20587
rect 6276 20544 6328 20553
rect 9772 20587 9824 20596
rect 9772 20553 9781 20587
rect 9781 20553 9815 20587
rect 9815 20553 9824 20587
rect 9772 20544 9824 20553
rect 11980 20587 12032 20596
rect 11980 20553 11989 20587
rect 11989 20553 12023 20587
rect 12023 20553 12032 20587
rect 11980 20544 12032 20553
rect 5356 20519 5408 20528
rect 5356 20485 5365 20519
rect 5365 20485 5399 20519
rect 5399 20485 5408 20519
rect 5356 20476 5408 20485
rect 10876 20476 10928 20528
rect 7380 20451 7432 20460
rect 7380 20417 7389 20451
rect 7389 20417 7423 20451
rect 7423 20417 7432 20451
rect 7380 20408 7432 20417
rect 8300 20383 8352 20392
rect 3976 20272 4028 20324
rect 8300 20349 8309 20383
rect 8309 20349 8343 20383
rect 8343 20349 8352 20383
rect 8760 20383 8812 20392
rect 8300 20340 8352 20349
rect 8760 20349 8769 20383
rect 8769 20349 8803 20383
rect 8803 20349 8812 20383
rect 8760 20340 8812 20349
rect 9680 20340 9732 20392
rect 10416 20340 10468 20392
rect 4804 20315 4856 20324
rect 4804 20281 4813 20315
rect 4813 20281 4847 20315
rect 4847 20281 4856 20315
rect 4804 20272 4856 20281
rect 4896 20315 4948 20324
rect 4896 20281 4905 20315
rect 4905 20281 4939 20315
rect 4939 20281 4948 20315
rect 6920 20315 6972 20324
rect 4896 20272 4948 20281
rect 6920 20281 6929 20315
rect 6929 20281 6963 20315
rect 6963 20281 6972 20315
rect 6920 20272 6972 20281
rect 7012 20315 7064 20324
rect 7012 20281 7021 20315
rect 7021 20281 7055 20315
rect 7055 20281 7064 20315
rect 10692 20315 10744 20324
rect 7012 20272 7064 20281
rect 10692 20281 10701 20315
rect 10701 20281 10735 20315
rect 10735 20281 10744 20315
rect 10692 20272 10744 20281
rect 11612 20272 11664 20324
rect 11980 20272 12032 20324
rect 3884 20204 3936 20256
rect 4252 20247 4304 20256
rect 4252 20213 4261 20247
rect 4261 20213 4295 20247
rect 4295 20213 4304 20247
rect 4252 20204 4304 20213
rect 4436 20204 4488 20256
rect 4620 20247 4672 20256
rect 4620 20213 4629 20247
rect 4629 20213 4663 20247
rect 4663 20213 4672 20247
rect 4620 20204 4672 20213
rect 6644 20247 6696 20256
rect 6644 20213 6653 20247
rect 6653 20213 6687 20247
rect 6687 20213 6696 20247
rect 6644 20204 6696 20213
rect 7748 20204 7800 20256
rect 8484 20204 8536 20256
rect 9588 20204 9640 20256
rect 12072 20204 12124 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 4160 20000 4212 20052
rect 4896 20000 4948 20052
rect 4804 19932 4856 19984
rect 5540 19932 5592 19984
rect 5724 19932 5776 19984
rect 10876 20000 10928 20052
rect 6644 19932 6696 19984
rect 7840 19932 7892 19984
rect 4068 19864 4120 19916
rect 5356 19864 5408 19916
rect 9680 19864 9732 19916
rect 10048 19864 10100 19916
rect 10416 19864 10468 19916
rect 10692 19864 10744 19916
rect 11520 19864 11572 19916
rect 5540 19839 5592 19848
rect 5540 19805 5549 19839
rect 5549 19805 5583 19839
rect 5583 19805 5592 19839
rect 5540 19796 5592 19805
rect 7196 19796 7248 19848
rect 8300 19796 8352 19848
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 7932 19771 7984 19780
rect 7932 19737 7941 19771
rect 7941 19737 7975 19771
rect 7975 19737 7984 19771
rect 7932 19728 7984 19737
rect 9956 19771 10008 19780
rect 9956 19737 9965 19771
rect 9965 19737 9999 19771
rect 9999 19737 10008 19771
rect 9956 19728 10008 19737
rect 10508 19728 10560 19780
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8392 19660 8444 19669
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 4896 19456 4948 19508
rect 5724 19456 5776 19508
rect 7840 19499 7892 19508
rect 7840 19465 7849 19499
rect 7849 19465 7883 19499
rect 7883 19465 7892 19499
rect 7840 19456 7892 19465
rect 10416 19456 10468 19508
rect 10876 19499 10928 19508
rect 10876 19465 10885 19499
rect 10885 19465 10919 19499
rect 10919 19465 10928 19499
rect 10876 19456 10928 19465
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 7012 19320 7064 19372
rect 7932 19320 7984 19372
rect 3240 19295 3292 19304
rect 3240 19261 3249 19295
rect 3249 19261 3283 19295
rect 3283 19261 3292 19295
rect 3240 19252 3292 19261
rect 4068 19252 4120 19304
rect 4160 19252 4212 19304
rect 2412 19116 2464 19168
rect 3056 19184 3108 19236
rect 5540 19252 5592 19304
rect 5724 19184 5776 19236
rect 6644 19159 6696 19168
rect 6644 19125 6653 19159
rect 6653 19125 6687 19159
rect 6687 19125 6696 19159
rect 7104 19184 7156 19236
rect 8392 19320 8444 19372
rect 8944 19363 8996 19372
rect 8944 19329 8953 19363
rect 8953 19329 8987 19363
rect 8987 19329 8996 19363
rect 8944 19320 8996 19329
rect 9220 19295 9272 19304
rect 9220 19261 9229 19295
rect 9229 19261 9263 19295
rect 9263 19261 9272 19295
rect 9220 19252 9272 19261
rect 9864 19252 9916 19304
rect 10876 19252 10928 19304
rect 8392 19227 8444 19236
rect 8392 19193 8401 19227
rect 8401 19193 8435 19227
rect 8435 19193 8444 19227
rect 8392 19184 8444 19193
rect 9956 19184 10008 19236
rect 6644 19116 6696 19125
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 2780 18955 2832 18964
rect 2780 18921 2789 18955
rect 2789 18921 2823 18955
rect 2823 18921 2832 18955
rect 2780 18912 2832 18921
rect 3424 18912 3476 18964
rect 8300 18955 8352 18964
rect 5724 18844 5776 18896
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 9588 18912 9640 18964
rect 9956 18912 10008 18964
rect 10048 18912 10100 18964
rect 10600 18912 10652 18964
rect 6920 18844 6972 18896
rect 8024 18844 8076 18896
rect 2044 18819 2096 18828
rect 2044 18785 2062 18819
rect 2062 18785 2096 18819
rect 2044 18776 2096 18785
rect 3148 18776 3200 18828
rect 4436 18776 4488 18828
rect 3424 18708 3476 18760
rect 5724 18708 5776 18760
rect 5632 18640 5684 18692
rect 9772 18776 9824 18828
rect 10416 18844 10468 18896
rect 11244 18776 11296 18828
rect 13084 18776 13136 18828
rect 6184 18708 6236 18760
rect 8576 18708 8628 18760
rect 10416 18751 10468 18760
rect 10416 18717 10425 18751
rect 10425 18717 10459 18751
rect 10459 18717 10468 18751
rect 10416 18708 10468 18717
rect 7932 18683 7984 18692
rect 7932 18649 7941 18683
rect 7941 18649 7975 18683
rect 7975 18649 7984 18683
rect 7932 18640 7984 18649
rect 9864 18640 9916 18692
rect 11428 18640 11480 18692
rect 12256 18640 12308 18692
rect 3240 18572 3292 18624
rect 4160 18572 4212 18624
rect 4896 18572 4948 18624
rect 5264 18572 5316 18624
rect 5540 18572 5592 18624
rect 6828 18615 6880 18624
rect 6828 18581 6837 18615
rect 6837 18581 6871 18615
rect 6871 18581 6880 18615
rect 6828 18572 6880 18581
rect 11152 18572 11204 18624
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 2780 18368 2832 18420
rect 3148 18368 3200 18420
rect 5264 18368 5316 18420
rect 5816 18368 5868 18420
rect 8024 18411 8076 18420
rect 4160 18275 4212 18284
rect 4160 18241 4169 18275
rect 4169 18241 4203 18275
rect 4203 18241 4212 18275
rect 4160 18232 4212 18241
rect 8024 18377 8033 18411
rect 8033 18377 8067 18411
rect 8067 18377 8076 18411
rect 8024 18368 8076 18377
rect 8484 18411 8536 18420
rect 8484 18377 8493 18411
rect 8493 18377 8527 18411
rect 8527 18377 8536 18411
rect 8484 18368 8536 18377
rect 9588 18411 9640 18420
rect 9588 18377 9597 18411
rect 9597 18377 9631 18411
rect 9631 18377 9640 18411
rect 9588 18368 9640 18377
rect 10140 18368 10192 18420
rect 6644 18300 6696 18352
rect 9864 18300 9916 18352
rect 2504 18164 2556 18216
rect 3424 18207 3476 18216
rect 3424 18173 3433 18207
rect 3433 18173 3467 18207
rect 3467 18173 3476 18207
rect 3424 18164 3476 18173
rect 3884 18207 3936 18216
rect 3884 18173 3893 18207
rect 3893 18173 3927 18207
rect 3927 18173 3936 18207
rect 3884 18164 3936 18173
rect 4896 18164 4948 18216
rect 5540 18207 5592 18216
rect 5540 18173 5549 18207
rect 5549 18173 5583 18207
rect 5583 18173 5592 18207
rect 5540 18164 5592 18173
rect 5816 18164 5868 18216
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 2044 18139 2096 18148
rect 2044 18105 2053 18139
rect 2053 18105 2087 18139
rect 2087 18105 2096 18139
rect 2044 18096 2096 18105
rect 5356 18096 5408 18148
rect 5724 18139 5776 18148
rect 5724 18105 5733 18139
rect 5733 18105 5767 18139
rect 5767 18105 5776 18139
rect 5724 18096 5776 18105
rect 10508 18368 10560 18420
rect 11244 18368 11296 18420
rect 11520 18232 11572 18284
rect 9772 18164 9824 18216
rect 10416 18164 10468 18216
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 9588 18096 9640 18148
rect 4436 18028 4488 18080
rect 10692 18071 10744 18080
rect 10692 18037 10701 18071
rect 10701 18037 10735 18071
rect 10735 18037 10744 18071
rect 10692 18028 10744 18037
rect 11060 18071 11112 18080
rect 11060 18037 11069 18071
rect 11069 18037 11103 18071
rect 11103 18037 11112 18071
rect 11060 18028 11112 18037
rect 12624 18071 12676 18080
rect 12624 18037 12633 18071
rect 12633 18037 12667 18071
rect 12667 18037 12676 18071
rect 12624 18028 12676 18037
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 3884 17824 3936 17876
rect 4804 17824 4856 17876
rect 5724 17824 5776 17876
rect 6644 17824 6696 17876
rect 3240 17756 3292 17808
rect 5816 17799 5868 17808
rect 3056 17688 3108 17740
rect 4160 17731 4212 17740
rect 4160 17697 4178 17731
rect 4178 17697 4212 17731
rect 4160 17688 4212 17697
rect 5080 17731 5132 17740
rect 5080 17697 5089 17731
rect 5089 17697 5123 17731
rect 5123 17697 5132 17731
rect 5080 17688 5132 17697
rect 5540 17731 5592 17740
rect 5540 17697 5549 17731
rect 5549 17697 5583 17731
rect 5583 17697 5592 17731
rect 5540 17688 5592 17697
rect 5816 17765 5825 17799
rect 5825 17765 5859 17799
rect 5859 17765 5868 17799
rect 5816 17756 5868 17765
rect 7380 17799 7432 17808
rect 7380 17765 7389 17799
rect 7389 17765 7423 17799
rect 7423 17765 7432 17799
rect 7380 17756 7432 17765
rect 9588 17824 9640 17876
rect 10600 17824 10652 17876
rect 6184 17688 6236 17740
rect 9772 17756 9824 17808
rect 10692 17756 10744 17808
rect 11520 17731 11572 17740
rect 5632 17620 5684 17672
rect 8300 17620 8352 17672
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 12808 17731 12860 17740
rect 12808 17697 12817 17731
rect 12817 17697 12851 17731
rect 12851 17697 12860 17731
rect 12808 17688 12860 17697
rect 13084 17731 13136 17740
rect 13084 17697 13093 17731
rect 13093 17697 13127 17731
rect 13127 17697 13136 17731
rect 13084 17688 13136 17697
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 8852 17552 8904 17604
rect 9864 17552 9916 17604
rect 12900 17595 12952 17604
rect 12900 17561 12909 17595
rect 12909 17561 12943 17595
rect 12943 17561 12952 17595
rect 12900 17552 12952 17561
rect 2504 17527 2556 17536
rect 2504 17493 2513 17527
rect 2513 17493 2547 17527
rect 2547 17493 2556 17527
rect 2504 17484 2556 17493
rect 4712 17484 4764 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 9680 17484 9732 17536
rect 10968 17484 11020 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 5080 17280 5132 17332
rect 5540 17280 5592 17332
rect 8300 17323 8352 17332
rect 8300 17289 8309 17323
rect 8309 17289 8343 17323
rect 8343 17289 8352 17323
rect 8300 17280 8352 17289
rect 9864 17280 9916 17332
rect 3056 17255 3108 17264
rect 3056 17221 3065 17255
rect 3065 17221 3099 17255
rect 3099 17221 3108 17255
rect 3056 17212 3108 17221
rect 11520 17280 11572 17332
rect 12808 17280 12860 17332
rect 4620 17144 4672 17196
rect 5080 17144 5132 17196
rect 6920 17144 6972 17196
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 4988 17051 5040 17060
rect 4988 17017 4997 17051
rect 4997 17017 5031 17051
rect 5031 17017 5040 17051
rect 4988 17008 5040 17017
rect 7196 17119 7248 17128
rect 7196 17085 7205 17119
rect 7205 17085 7239 17119
rect 7239 17085 7248 17119
rect 7196 17076 7248 17085
rect 13084 17212 13136 17264
rect 8576 17144 8628 17196
rect 7748 17076 7800 17128
rect 9128 17144 9180 17196
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 10600 17119 10652 17128
rect 7564 17008 7616 17060
rect 8300 17008 8352 17060
rect 8852 17008 8904 17060
rect 10600 17085 10609 17119
rect 10609 17085 10643 17119
rect 10643 17085 10652 17119
rect 10600 17076 10652 17085
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 11244 17076 11296 17128
rect 9680 17008 9732 17060
rect 9588 16983 9640 16992
rect 9588 16949 9597 16983
rect 9597 16949 9631 16983
rect 9631 16949 9640 16983
rect 9588 16940 9640 16949
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 4988 16736 5040 16788
rect 5632 16736 5684 16788
rect 7196 16779 7248 16788
rect 7196 16745 7205 16779
rect 7205 16745 7239 16779
rect 7239 16745 7248 16779
rect 7196 16736 7248 16745
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 9128 16779 9180 16788
rect 9128 16745 9137 16779
rect 9137 16745 9171 16779
rect 9171 16745 9180 16779
rect 9128 16736 9180 16745
rect 9404 16736 9456 16788
rect 4712 16643 4764 16652
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 6092 16600 6144 16652
rect 10876 16736 10928 16788
rect 12440 16736 12492 16788
rect 12808 16668 12860 16720
rect 7564 16643 7616 16652
rect 7564 16609 7573 16643
rect 7573 16609 7607 16643
rect 7607 16609 7616 16643
rect 7564 16600 7616 16609
rect 7748 16600 7800 16652
rect 8024 16600 8076 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10600 16600 10652 16652
rect 12440 16600 12492 16652
rect 13544 16643 13596 16652
rect 13544 16609 13588 16643
rect 13588 16609 13596 16643
rect 13544 16600 13596 16609
rect 4436 16532 4488 16584
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 8208 16532 8260 16584
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 9772 16507 9824 16516
rect 9772 16473 9781 16507
rect 9781 16473 9815 16507
rect 9815 16473 9824 16507
rect 9772 16464 9824 16473
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 3240 16192 3292 16244
rect 5264 16192 5316 16244
rect 6092 16235 6144 16244
rect 6092 16201 6101 16235
rect 6101 16201 6135 16235
rect 6135 16201 6144 16235
rect 6092 16192 6144 16201
rect 8208 16192 8260 16244
rect 9772 16192 9824 16244
rect 10968 16192 11020 16244
rect 13544 16235 13596 16244
rect 13544 16201 13553 16235
rect 13553 16201 13587 16235
rect 13587 16201 13596 16235
rect 13544 16192 13596 16201
rect 4436 16056 4488 16108
rect 4988 16056 5040 16108
rect 4252 15988 4304 16040
rect 11244 16124 11296 16176
rect 11980 16124 12032 16176
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 11152 16056 11204 16108
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 8852 16031 8904 16040
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 5264 15920 5316 15972
rect 8760 15920 8812 15972
rect 9404 15920 9456 15972
rect 10968 15963 11020 15972
rect 10968 15929 10977 15963
rect 10977 15929 11011 15963
rect 11011 15929 11020 15963
rect 10968 15920 11020 15929
rect 11980 15920 12032 15972
rect 5908 15852 5960 15904
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 9588 15895 9640 15904
rect 9588 15861 9597 15895
rect 9597 15861 9631 15895
rect 9631 15861 9640 15895
rect 9588 15852 9640 15861
rect 12440 15852 12492 15904
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 4712 15648 4764 15700
rect 7564 15648 7616 15700
rect 9496 15691 9548 15700
rect 5264 15580 5316 15632
rect 5908 15580 5960 15632
rect 6552 15623 6604 15632
rect 6552 15589 6561 15623
rect 6561 15589 6595 15623
rect 6595 15589 6604 15623
rect 6552 15580 6604 15589
rect 4804 15512 4856 15564
rect 5540 15512 5592 15564
rect 8852 15580 8904 15632
rect 8024 15512 8076 15564
rect 9496 15657 9505 15691
rect 9505 15657 9539 15691
rect 9539 15657 9548 15691
rect 9496 15648 9548 15657
rect 11152 15691 11204 15700
rect 11152 15657 11161 15691
rect 11161 15657 11195 15691
rect 11195 15657 11204 15691
rect 11152 15648 11204 15657
rect 10048 15580 10100 15632
rect 11796 15623 11848 15632
rect 9496 15512 9548 15564
rect 9680 15512 9732 15564
rect 11796 15589 11805 15623
rect 11805 15589 11839 15623
rect 11839 15589 11848 15623
rect 11796 15580 11848 15589
rect 11980 15580 12032 15632
rect 13544 15580 13596 15632
rect 4160 15444 4212 15496
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 6920 15487 6972 15496
rect 6920 15453 6929 15487
rect 6929 15453 6963 15487
rect 6963 15453 6972 15487
rect 6920 15444 6972 15453
rect 8116 15444 8168 15496
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 6828 15376 6880 15428
rect 8208 15376 8260 15428
rect 5632 15308 5684 15360
rect 6460 15308 6512 15360
rect 7012 15308 7064 15360
rect 7380 15308 7432 15360
rect 8116 15308 8168 15360
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 4068 15104 4120 15156
rect 5264 15147 5316 15156
rect 5264 15113 5273 15147
rect 5273 15113 5307 15147
rect 5307 15113 5316 15147
rect 5264 15104 5316 15113
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 8208 15104 8260 15156
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 9404 15147 9456 15156
rect 8300 15104 8352 15113
rect 9404 15113 9413 15147
rect 9413 15113 9447 15147
rect 9447 15113 9456 15147
rect 9404 15104 9456 15113
rect 9772 15104 9824 15156
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 2504 14900 2556 14952
rect 3424 15036 3476 15088
rect 4712 15036 4764 15088
rect 4344 14968 4396 15020
rect 6644 15036 6696 15088
rect 6920 14968 6972 15020
rect 8116 14968 8168 15020
rect 8300 14900 8352 14952
rect 8668 14900 8720 14952
rect 11796 14900 11848 14952
rect 4068 14832 4120 14884
rect 5816 14832 5868 14884
rect 4620 14764 4672 14816
rect 6828 14764 6880 14816
rect 10876 14832 10928 14884
rect 11336 14832 11388 14884
rect 11704 14832 11756 14884
rect 8484 14807 8536 14816
rect 8484 14773 8493 14807
rect 8493 14773 8527 14807
rect 8527 14773 8536 14807
rect 8484 14764 8536 14773
rect 9680 14764 9732 14816
rect 10048 14764 10100 14816
rect 10600 14764 10652 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 2504 14603 2556 14612
rect 2504 14569 2513 14603
rect 2513 14569 2547 14603
rect 2547 14569 2556 14603
rect 2504 14560 2556 14569
rect 3148 14560 3200 14612
rect 5908 14560 5960 14612
rect 6828 14603 6880 14612
rect 6828 14569 6837 14603
rect 6837 14569 6871 14603
rect 6871 14569 6880 14603
rect 6828 14560 6880 14569
rect 8852 14603 8904 14612
rect 8852 14569 8861 14603
rect 8861 14569 8895 14603
rect 8895 14569 8904 14603
rect 8852 14560 8904 14569
rect 9496 14603 9548 14612
rect 9496 14569 9505 14603
rect 9505 14569 9539 14603
rect 9539 14569 9548 14603
rect 9496 14560 9548 14569
rect 9680 14560 9732 14612
rect 4620 14492 4672 14544
rect 7564 14492 7616 14544
rect 6368 14424 6420 14476
rect 6736 14424 6788 14476
rect 7748 14424 7800 14476
rect 8484 14424 8536 14476
rect 9588 14424 9640 14476
rect 11336 14424 11388 14476
rect 4160 14356 4212 14408
rect 4252 14288 4304 14340
rect 4988 14288 5040 14340
rect 6828 14288 6880 14340
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 5816 14220 5868 14272
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 8668 14220 8720 14272
rect 10692 14220 10744 14272
rect 10968 14220 11020 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 4160 14016 4212 14068
rect 4712 14016 4764 14068
rect 6000 14016 6052 14068
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 7564 14016 7616 14068
rect 9588 14016 9640 14068
rect 10968 14059 11020 14068
rect 10968 14025 10977 14059
rect 10977 14025 11011 14059
rect 11011 14025 11020 14059
rect 10968 14016 11020 14025
rect 5816 13991 5868 14000
rect 5816 13957 5825 13991
rect 5825 13957 5859 13991
rect 5859 13957 5868 13991
rect 5816 13948 5868 13957
rect 3424 13812 3476 13864
rect 4160 13880 4212 13932
rect 5540 13880 5592 13932
rect 7104 13880 7156 13932
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 9680 13880 9732 13889
rect 11336 13948 11388 14000
rect 4988 13812 5040 13864
rect 8300 13812 8352 13864
rect 3884 13719 3936 13728
rect 3884 13685 3893 13719
rect 3893 13685 3927 13719
rect 3927 13685 3936 13719
rect 3884 13676 3936 13685
rect 7564 13744 7616 13796
rect 10600 13787 10652 13796
rect 6000 13676 6052 13728
rect 10600 13753 10609 13787
rect 10609 13753 10643 13787
rect 10643 13753 10652 13787
rect 10600 13744 10652 13753
rect 10692 13676 10744 13728
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 4068 13472 4120 13524
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 7564 13472 7616 13524
rect 7748 13515 7800 13524
rect 7748 13481 7757 13515
rect 7757 13481 7791 13515
rect 7791 13481 7800 13515
rect 7748 13472 7800 13481
rect 3424 13404 3476 13456
rect 5264 13404 5316 13456
rect 8208 13447 8260 13456
rect 8208 13413 8217 13447
rect 8217 13413 8251 13447
rect 8251 13413 8260 13447
rect 8208 13404 8260 13413
rect 10048 13447 10100 13456
rect 10048 13413 10057 13447
rect 10057 13413 10091 13447
rect 10091 13413 10100 13447
rect 10048 13404 10100 13413
rect 10600 13447 10652 13456
rect 10600 13413 10609 13447
rect 10609 13413 10643 13447
rect 10643 13413 10652 13447
rect 10600 13404 10652 13413
rect 2964 13379 3016 13388
rect 2964 13345 3008 13379
rect 3008 13345 3016 13379
rect 2964 13336 3016 13345
rect 4712 13336 4764 13388
rect 11336 13336 11388 13388
rect 6828 13311 6880 13320
rect 4252 13200 4304 13252
rect 4988 13200 5040 13252
rect 4344 13132 4396 13184
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 8576 13268 8628 13320
rect 8852 13268 8904 13320
rect 9588 13268 9640 13320
rect 6000 13175 6052 13184
rect 6000 13141 6009 13175
rect 6009 13141 6043 13175
rect 6043 13141 6052 13175
rect 6000 13132 6052 13141
rect 8760 13132 8812 13184
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 2964 12971 3016 12980
rect 2964 12937 2973 12971
rect 2973 12937 3007 12971
rect 3007 12937 3016 12971
rect 2964 12928 3016 12937
rect 3332 12928 3384 12980
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 8300 12928 8352 12980
rect 5172 12860 5224 12912
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 4988 12792 5040 12844
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 3424 12724 3476 12776
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 8484 12860 8536 12912
rect 11336 12860 11388 12912
rect 8760 12792 8812 12844
rect 8852 12792 8904 12844
rect 10048 12792 10100 12844
rect 10692 12767 10744 12776
rect 10692 12733 10701 12767
rect 10701 12733 10735 12767
rect 10735 12733 10744 12767
rect 10692 12724 10744 12733
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 7380 12656 7432 12708
rect 8300 12656 8352 12708
rect 10508 12656 10560 12708
rect 11336 12656 11388 12708
rect 6000 12588 6052 12640
rect 7748 12631 7800 12640
rect 7748 12597 7757 12631
rect 7757 12597 7791 12631
rect 7791 12597 7800 12631
rect 7748 12588 7800 12597
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 3056 12384 3108 12436
rect 3332 12384 3384 12436
rect 3516 12384 3568 12436
rect 4068 12384 4120 12436
rect 4252 12384 4304 12436
rect 6000 12427 6052 12436
rect 6000 12393 6009 12427
rect 6009 12393 6043 12427
rect 6043 12393 6052 12427
rect 6000 12384 6052 12393
rect 7656 12384 7708 12436
rect 4988 12316 5040 12368
rect 7012 12316 7064 12368
rect 8208 12359 8260 12368
rect 8208 12325 8217 12359
rect 8217 12325 8251 12359
rect 8251 12325 8260 12359
rect 8208 12316 8260 12325
rect 8576 12384 8628 12436
rect 9588 12384 9640 12436
rect 10692 12427 10744 12436
rect 10692 12393 10701 12427
rect 10701 12393 10735 12427
rect 10735 12393 10744 12427
rect 10692 12384 10744 12393
rect 11980 12316 12032 12368
rect 12440 12316 12492 12368
rect 3056 12291 3108 12300
rect 3056 12257 3074 12291
rect 3074 12257 3108 12291
rect 3056 12248 3108 12257
rect 7748 12248 7800 12300
rect 9956 12291 10008 12300
rect 9956 12257 9965 12291
rect 9965 12257 9999 12291
rect 9999 12257 10008 12291
rect 9956 12248 10008 12257
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 12256 12248 12308 12300
rect 4804 12180 4856 12232
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 6828 12180 6880 12232
rect 8576 12180 8628 12232
rect 7104 12155 7156 12164
rect 7104 12121 7113 12155
rect 7113 12121 7147 12155
rect 7147 12121 7156 12155
rect 7104 12112 7156 12121
rect 8484 12112 8536 12164
rect 8760 12112 8812 12164
rect 10048 12044 10100 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 3056 11883 3108 11892
rect 3056 11849 3065 11883
rect 3065 11849 3099 11883
rect 3099 11849 3108 11883
rect 3056 11840 3108 11849
rect 4988 11883 5040 11892
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 6828 11840 6880 11892
rect 7012 11883 7064 11892
rect 7012 11849 7021 11883
rect 7021 11849 7055 11883
rect 7055 11849 7064 11883
rect 7012 11840 7064 11849
rect 7380 11840 7432 11892
rect 8208 11840 8260 11892
rect 4620 11704 4672 11756
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 4252 11611 4304 11620
rect 4252 11577 4261 11611
rect 4261 11577 4295 11611
rect 4295 11577 4304 11611
rect 4252 11568 4304 11577
rect 8668 11772 8720 11824
rect 10140 11840 10192 11892
rect 10968 11840 11020 11892
rect 11428 11883 11480 11892
rect 11428 11849 11437 11883
rect 11437 11849 11471 11883
rect 11471 11849 11480 11883
rect 11428 11840 11480 11849
rect 10048 11815 10100 11824
rect 10048 11781 10057 11815
rect 10057 11781 10091 11815
rect 10091 11781 10100 11815
rect 10048 11772 10100 11781
rect 5264 11704 5316 11756
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 10968 11679 11020 11688
rect 10968 11645 11012 11679
rect 11012 11645 11020 11679
rect 10968 11636 11020 11645
rect 5816 11611 5868 11620
rect 5080 11500 5132 11552
rect 5816 11577 5825 11611
rect 5825 11577 5859 11611
rect 5859 11577 5868 11611
rect 5816 11568 5868 11577
rect 7380 11568 7432 11620
rect 9496 11568 9548 11620
rect 9956 11500 10008 11552
rect 12072 11500 12124 11552
rect 12256 11500 12308 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 4068 11296 4120 11348
rect 5080 11296 5132 11348
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 9496 11339 9548 11348
rect 9496 11305 9505 11339
rect 9505 11305 9539 11339
rect 9539 11305 9548 11339
rect 9496 11296 9548 11305
rect 4344 11228 4396 11280
rect 7380 11228 7432 11280
rect 9864 11271 9916 11280
rect 9864 11237 9873 11271
rect 9873 11237 9907 11271
rect 9907 11237 9916 11271
rect 9864 11228 9916 11237
rect 10048 11228 10100 11280
rect 11428 11271 11480 11280
rect 11428 11237 11437 11271
rect 11437 11237 11471 11271
rect 11471 11237 11480 11271
rect 11428 11228 11480 11237
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 2964 11203 3016 11212
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 4160 11160 4212 11212
rect 5172 11160 5224 11212
rect 6184 11160 6236 11212
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 5448 11092 5500 11144
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 10600 11092 10652 11144
rect 11612 11135 11664 11144
rect 3056 11024 3108 11076
rect 3884 11024 3936 11076
rect 4804 11024 4856 11076
rect 6828 11024 6880 11076
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 4068 10956 4120 11008
rect 8116 10956 8168 11008
rect 11520 11024 11572 11076
rect 8392 10956 8444 11008
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 2964 10752 3016 10804
rect 4068 10752 4120 10804
rect 4344 10795 4396 10804
rect 4344 10761 4353 10795
rect 4353 10761 4387 10795
rect 4387 10761 4396 10795
rect 4344 10752 4396 10761
rect 5540 10752 5592 10804
rect 7380 10795 7432 10804
rect 7380 10761 7389 10795
rect 7389 10761 7423 10795
rect 7423 10761 7432 10795
rect 7380 10752 7432 10761
rect 8392 10752 8444 10804
rect 9864 10752 9916 10804
rect 10600 10795 10652 10804
rect 10600 10761 10609 10795
rect 10609 10761 10643 10795
rect 10643 10761 10652 10795
rect 10600 10752 10652 10761
rect 11428 10752 11480 10804
rect 4712 10684 4764 10736
rect 9404 10684 9456 10736
rect 4160 10616 4212 10668
rect 10048 10616 10100 10668
rect 7564 10548 7616 10600
rect 4344 10480 4396 10532
rect 4712 10480 4764 10532
rect 7380 10480 7432 10532
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 3884 10455 3936 10464
rect 3884 10421 3893 10455
rect 3893 10421 3927 10455
rect 3927 10421 3936 10455
rect 3884 10412 3936 10421
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 5724 10412 5776 10464
rect 6184 10412 6236 10464
rect 10324 10548 10376 10600
rect 9312 10523 9364 10532
rect 9312 10489 9321 10523
rect 9321 10489 9355 10523
rect 9355 10489 9364 10523
rect 9312 10480 9364 10489
rect 9496 10480 9548 10532
rect 11520 10412 11572 10464
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 3976 10208 4028 10260
rect 4160 10208 4212 10260
rect 7380 10208 7432 10260
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 4712 10183 4764 10192
rect 4712 10149 4721 10183
rect 4721 10149 4755 10183
rect 4755 10149 4764 10183
rect 4712 10140 4764 10149
rect 5356 10140 5408 10192
rect 8116 10140 8168 10192
rect 8760 10183 8812 10192
rect 8760 10149 8769 10183
rect 8769 10149 8803 10183
rect 8803 10149 8812 10183
rect 8760 10140 8812 10149
rect 3056 10115 3108 10124
rect 3056 10081 3074 10115
rect 3074 10081 3108 10115
rect 3056 10072 3108 10081
rect 4528 10072 4580 10124
rect 9772 10115 9824 10124
rect 9772 10081 9790 10115
rect 9790 10081 9824 10115
rect 9772 10072 9824 10081
rect 10784 10072 10836 10124
rect 4068 10004 4120 10056
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 6920 10004 6972 10056
rect 8392 10004 8444 10056
rect 4528 9936 4580 9988
rect 7472 9936 7524 9988
rect 7564 9868 7616 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 4528 9664 4580 9716
rect 8116 9707 8168 9716
rect 8116 9673 8125 9707
rect 8125 9673 8159 9707
rect 8159 9673 8168 9707
rect 8116 9664 8168 9673
rect 8208 9664 8260 9716
rect 8300 9664 8352 9716
rect 10232 9664 10284 9716
rect 10416 9664 10468 9716
rect 4068 9639 4120 9648
rect 4068 9605 4077 9639
rect 4077 9605 4111 9639
rect 4111 9605 4120 9639
rect 4068 9596 4120 9605
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 8392 9596 8444 9648
rect 11980 9596 12032 9648
rect 13820 9596 13872 9648
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 7564 9571 7616 9580
rect 6552 9528 6604 9537
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 9588 9528 9640 9580
rect 7196 9460 7248 9512
rect 5356 9435 5408 9444
rect 5356 9401 5365 9435
rect 5365 9401 5399 9435
rect 5399 9401 5408 9435
rect 5356 9392 5408 9401
rect 7104 9392 7156 9444
rect 8392 9460 8444 9512
rect 8852 9460 8904 9512
rect 8668 9392 8720 9444
rect 10140 9392 10192 9444
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 3332 9324 3384 9376
rect 8576 9324 8628 9376
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 5356 9120 5408 9172
rect 4620 9052 4672 9104
rect 7288 9095 7340 9104
rect 7288 9061 7297 9095
rect 7297 9061 7331 9095
rect 7331 9061 7340 9095
rect 7288 9052 7340 9061
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 6184 8984 6236 9036
rect 7104 9027 7156 9036
rect 7104 8993 7113 9027
rect 7113 8993 7147 9027
rect 7147 8993 7156 9027
rect 7104 8984 7156 8993
rect 8300 8984 8352 9036
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 8760 8848 8812 8900
rect 5356 8823 5408 8832
rect 5356 8789 5365 8823
rect 5365 8789 5399 8823
rect 5399 8789 5408 8823
rect 5356 8780 5408 8789
rect 7656 8823 7708 8832
rect 7656 8789 7665 8823
rect 7665 8789 7699 8823
rect 7699 8789 7708 8823
rect 7656 8780 7708 8789
rect 8668 8780 8720 8832
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 4436 8576 4488 8628
rect 4620 8551 4672 8560
rect 4620 8517 4629 8551
rect 4629 8517 4663 8551
rect 4663 8517 4672 8551
rect 4620 8508 4672 8517
rect 4252 8372 4304 8424
rect 4712 8372 4764 8424
rect 8300 8576 8352 8628
rect 7656 8440 7708 8492
rect 5356 8372 5408 8424
rect 6184 8415 6236 8424
rect 6184 8381 6193 8415
rect 6193 8381 6227 8415
rect 6227 8381 6236 8415
rect 6184 8372 6236 8381
rect 8668 8415 8720 8424
rect 4344 8347 4396 8356
rect 4344 8313 4353 8347
rect 4353 8313 4387 8347
rect 4387 8313 4396 8347
rect 4344 8304 4396 8313
rect 6736 8304 6788 8356
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 8760 8372 8812 8424
rect 7380 8304 7432 8356
rect 6644 8236 6696 8288
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 3516 8032 3568 8084
rect 4252 8075 4304 8084
rect 4252 8041 4261 8075
rect 4261 8041 4295 8075
rect 4295 8041 4304 8075
rect 4252 8032 4304 8041
rect 4804 8075 4856 8084
rect 4804 8041 4813 8075
rect 4813 8041 4847 8075
rect 4847 8041 4856 8075
rect 4804 8032 4856 8041
rect 7656 8032 7708 8084
rect 6644 8007 6696 8016
rect 6644 7973 6653 8007
rect 6653 7973 6687 8007
rect 6687 7973 6696 8007
rect 6644 7964 6696 7973
rect 8208 8007 8260 8016
rect 8208 7973 8217 8007
rect 8217 7973 8251 8007
rect 8251 7973 8260 8007
rect 8208 7964 8260 7973
rect 8760 7964 8812 8016
rect 4896 7939 4948 7948
rect 4896 7905 4905 7939
rect 4905 7905 4939 7939
rect 4939 7905 4948 7939
rect 4896 7896 4948 7905
rect 5356 7939 5408 7948
rect 4252 7828 4304 7880
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 6828 7828 6880 7880
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 9312 7828 9364 7880
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 6644 7488 6696 7540
rect 7380 7488 7432 7540
rect 8208 7488 8260 7540
rect 3976 7420 4028 7472
rect 4620 7420 4672 7472
rect 6828 7420 6880 7472
rect 4436 7352 4488 7404
rect 4804 7352 4856 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 3516 7284 3568 7336
rect 4068 7216 4120 7268
rect 5080 7259 5132 7268
rect 5080 7225 5083 7259
rect 5083 7225 5117 7259
rect 5117 7225 5132 7259
rect 5080 7216 5132 7225
rect 7380 7216 7432 7268
rect 7840 7216 7892 7268
rect 9956 7488 10008 7540
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 11428 7327 11480 7336
rect 11428 7293 11437 7327
rect 11437 7293 11471 7327
rect 11471 7293 11480 7327
rect 11428 7284 11480 7293
rect 9496 7216 9548 7268
rect 9680 7216 9732 7268
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 5540 7148 5592 7200
rect 8760 7148 8812 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 3516 6944 3568 6996
rect 3976 6944 4028 6996
rect 4896 6987 4948 6996
rect 4896 6953 4905 6987
rect 4905 6953 4939 6987
rect 4939 6953 4948 6987
rect 4896 6944 4948 6953
rect 5172 6944 5224 6996
rect 5908 6944 5960 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 5080 6876 5132 6928
rect 7840 6919 7892 6928
rect 7840 6885 7843 6919
rect 7843 6885 7877 6919
rect 7877 6885 7892 6919
rect 7840 6876 7892 6885
rect 9864 6919 9916 6928
rect 9864 6885 9873 6919
rect 9873 6885 9907 6919
rect 9907 6885 9916 6919
rect 9864 6876 9916 6885
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 4344 6808 4396 6860
rect 6920 6808 6972 6860
rect 8208 6808 8260 6860
rect 4528 6740 4580 6792
rect 4988 6740 5040 6792
rect 2964 6672 3016 6724
rect 3332 6672 3384 6724
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 8116 6672 8168 6724
rect 9680 6672 9732 6724
rect 4160 6604 4212 6656
rect 5264 6604 5316 6656
rect 6000 6604 6052 6656
rect 8576 6604 8628 6656
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 2688 6400 2740 6452
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 3240 6443 3292 6452
rect 3240 6409 3249 6443
rect 3249 6409 3283 6443
rect 3283 6409 3292 6443
rect 3240 6400 3292 6409
rect 4528 6443 4580 6452
rect 4528 6409 4537 6443
rect 4537 6409 4571 6443
rect 4571 6409 4580 6443
rect 4528 6400 4580 6409
rect 5264 6400 5316 6452
rect 7380 6443 7432 6452
rect 5080 6332 5132 6384
rect 7380 6409 7389 6443
rect 7389 6409 7423 6443
rect 7423 6409 7432 6443
rect 7380 6400 7432 6409
rect 8576 6400 8628 6452
rect 9680 6400 9732 6452
rect 3516 6264 3568 6316
rect 4344 6264 4396 6316
rect 2504 6239 2556 6248
rect 2504 6205 2522 6239
rect 2522 6205 2556 6239
rect 2504 6196 2556 6205
rect 3240 6196 3292 6248
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 9864 6332 9916 6384
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 10048 6264 10100 6316
rect 4160 6171 4212 6180
rect 4160 6137 4169 6171
rect 4169 6137 4203 6171
rect 4203 6137 4212 6171
rect 4160 6128 4212 6137
rect 5356 6171 5408 6180
rect 5356 6137 5359 6171
rect 5359 6137 5393 6171
rect 5393 6137 5408 6171
rect 5356 6128 5408 6137
rect 7380 6128 7432 6180
rect 9312 6171 9364 6180
rect 9312 6137 9321 6171
rect 9321 6137 9355 6171
rect 9355 6137 9364 6171
rect 9312 6128 9364 6137
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 2504 5899 2556 5908
rect 2504 5865 2513 5899
rect 2513 5865 2547 5899
rect 2547 5865 2556 5899
rect 2504 5856 2556 5865
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 7288 5899 7340 5908
rect 7288 5865 7297 5899
rect 7297 5865 7331 5899
rect 7331 5865 7340 5899
rect 7288 5856 7340 5865
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 8760 5856 8812 5908
rect 4436 5788 4488 5840
rect 5908 5788 5960 5840
rect 6184 5788 6236 5840
rect 4344 5720 4396 5772
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7196 5720 7248 5729
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 6092 5652 6144 5704
rect 6920 5652 6972 5704
rect 9680 5763 9732 5772
rect 9680 5729 9724 5763
rect 9724 5729 9732 5763
rect 9680 5720 9732 5729
rect 5632 5584 5684 5636
rect 4068 5516 4120 5568
rect 4896 5516 4948 5568
rect 8760 5516 8812 5568
rect 9312 5516 9364 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 4436 5312 4488 5364
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 7196 5312 7248 5364
rect 9680 5355 9732 5364
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 4068 5244 4120 5296
rect 4344 5244 4396 5296
rect 6828 5244 6880 5296
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 3976 5108 4028 5160
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 9864 5151 9916 5160
rect 9864 5117 9908 5151
rect 9908 5117 9916 5151
rect 9864 5108 9916 5117
rect 4712 5040 4764 5092
rect 5264 5083 5316 5092
rect 5264 5049 5273 5083
rect 5273 5049 5307 5083
rect 5307 5049 5316 5083
rect 5264 5040 5316 5049
rect 5448 5040 5500 5092
rect 6092 5040 6144 5092
rect 8392 5083 8444 5092
rect 8392 5049 8401 5083
rect 8401 5049 8435 5083
rect 8435 5049 8444 5083
rect 8392 5040 8444 5049
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 8208 5015 8260 5024
rect 8208 4981 8217 5015
rect 8217 4981 8251 5015
rect 8251 4981 8260 5015
rect 8208 4972 8260 4981
rect 9772 4972 9824 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 3976 4768 4028 4820
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 5264 4768 5316 4820
rect 7104 4811 7156 4820
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 5356 4700 5408 4752
rect 7380 4700 7432 4752
rect 2780 4632 2832 4684
rect 7288 4675 7340 4684
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 10324 4632 10376 4684
rect 10692 4675 10744 4684
rect 10692 4641 10736 4675
rect 10736 4641 10744 4675
rect 10692 4632 10744 4641
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 8392 4564 8444 4616
rect 8852 4496 8904 4548
rect 2596 4428 2648 4480
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 5632 4428 5684 4437
rect 6092 4428 6144 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 2780 4224 2832 4276
rect 3424 4267 3476 4276
rect 3424 4233 3433 4267
rect 3433 4233 3467 4267
rect 3467 4233 3476 4267
rect 3424 4224 3476 4233
rect 4436 4224 4488 4276
rect 5356 4224 5408 4276
rect 8208 4224 8260 4276
rect 10324 4267 10376 4276
rect 2228 4020 2280 4072
rect 3240 4156 3292 4208
rect 4712 4156 4764 4208
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 7288 4156 7340 4208
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 3700 3995 3752 4004
rect 3700 3961 3709 3995
rect 3709 3961 3743 3995
rect 3743 3961 3752 3995
rect 3700 3952 3752 3961
rect 3792 3995 3844 4004
rect 3792 3961 3801 3995
rect 3801 3961 3835 3995
rect 3835 3961 3844 3995
rect 4344 3995 4396 4004
rect 3792 3952 3844 3961
rect 4344 3961 4353 3995
rect 4353 3961 4387 3995
rect 4387 3961 4396 3995
rect 4344 3952 4396 3961
rect 1400 3884 1452 3936
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 2136 3884 2188 3893
rect 5448 3952 5500 4004
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 6184 3952 6236 4004
rect 7380 3952 7432 4004
rect 10324 4233 10333 4267
rect 10333 4233 10367 4267
rect 10367 4233 10376 4267
rect 10324 4224 10376 4233
rect 10692 4224 10744 4276
rect 8852 4156 8904 4208
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 9588 4088 9640 4140
rect 10324 4020 10376 4072
rect 5540 3884 5592 3936
rect 8208 3884 8260 3936
rect 11060 3952 11112 4004
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 3792 3680 3844 3732
rect 5264 3680 5316 3732
rect 7380 3680 7432 3732
rect 8024 3680 8076 3732
rect 2596 3612 2648 3664
rect 4436 3655 4488 3664
rect 4436 3621 4439 3655
rect 4439 3621 4473 3655
rect 4473 3621 4488 3655
rect 4436 3612 4488 3621
rect 5448 3612 5500 3664
rect 6000 3655 6052 3664
rect 6000 3621 6009 3655
rect 6009 3621 6043 3655
rect 6043 3621 6052 3655
rect 6000 3612 6052 3621
rect 8208 3655 8260 3664
rect 8208 3621 8217 3655
rect 8217 3621 8251 3655
rect 8251 3621 8260 3655
rect 8208 3612 8260 3621
rect 9220 3612 9272 3664
rect 2320 3544 2372 3596
rect 3148 3544 3200 3596
rect 5264 3544 5316 3596
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 10140 3544 10192 3596
rect 11336 3544 11388 3596
rect 2504 3476 2556 3528
rect 2688 3476 2740 3528
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 9588 3476 9640 3528
rect 2780 3340 2832 3392
rect 4252 3340 4304 3392
rect 9312 3340 9364 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 2320 3136 2372 3188
rect 5264 3136 5316 3188
rect 6000 3136 6052 3188
rect 8208 3136 8260 3188
rect 9588 3136 9640 3188
rect 10140 3136 10192 3188
rect 11336 3136 11388 3188
rect 2596 3068 2648 3120
rect 8760 3111 8812 3120
rect 8760 3077 8769 3111
rect 8769 3077 8803 3111
rect 8803 3077 8812 3111
rect 8760 3068 8812 3077
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 5908 3000 5960 3052
rect 8024 3000 8076 3052
rect 1216 2932 1268 2984
rect 1676 2975 1728 2984
rect 1676 2941 1694 2975
rect 1694 2941 1728 2975
rect 1676 2932 1728 2941
rect 2780 2907 2832 2916
rect 2780 2873 2789 2907
rect 2789 2873 2823 2907
rect 2823 2873 2832 2907
rect 2780 2864 2832 2873
rect 3056 2864 3108 2916
rect 3516 2932 3568 2984
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 9864 3000 9916 3052
rect 6828 2932 6880 2941
rect 10784 2975 10836 2984
rect 10784 2941 10828 2975
rect 10828 2941 10836 2975
rect 10784 2932 10836 2941
rect 2320 2796 2372 2848
rect 4436 2864 4488 2916
rect 8300 2907 8352 2916
rect 8300 2873 8309 2907
rect 8309 2873 8343 2907
rect 8343 2873 8352 2907
rect 8300 2864 8352 2873
rect 4344 2796 4396 2848
rect 7012 2839 7064 2848
rect 7012 2805 7021 2839
rect 7021 2805 7055 2839
rect 7055 2805 7064 2839
rect 7012 2796 7064 2805
rect 10140 2796 10192 2848
rect 10324 2796 10376 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 2412 2592 2464 2644
rect 2872 2592 2924 2644
rect 4160 2592 4212 2644
rect 4344 2592 4396 2644
rect 4068 2524 4120 2576
rect 4988 2567 5040 2576
rect 4988 2533 4997 2567
rect 4997 2533 5031 2567
rect 5031 2533 5040 2567
rect 4988 2524 5040 2533
rect 6000 2592 6052 2644
rect 6184 2524 6236 2576
rect 7012 2567 7064 2576
rect 7012 2533 7021 2567
rect 7021 2533 7055 2567
rect 7055 2533 7064 2567
rect 7012 2524 7064 2533
rect 8208 2592 8260 2644
rect 9496 2592 9548 2644
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12072 2592 12124 2601
rect 10232 2456 10284 2508
rect 13176 2499 13228 2508
rect 13176 2465 13185 2499
rect 13185 2465 13219 2499
rect 13219 2465 13228 2499
rect 13176 2456 13228 2465
rect 2688 2388 2740 2440
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 4988 2388 5040 2440
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 11888 2320 11940 2372
rect 14188 2320 14240 2372
rect 8392 2252 8444 2304
rect 12348 2252 12400 2304
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 3884 1980 3936 2032
rect 4620 1980 4672 2032
rect 5172 552 5224 604
rect 5724 552 5776 604
<< metal2 >>
rect 386 39520 442 40000
rect 1214 39520 1270 40000
rect 2134 39522 2190 40000
rect 1412 39520 2190 39522
rect 3054 39520 3110 40000
rect 3882 39520 3938 40000
rect 4802 39522 4858 40000
rect 4802 39520 5028 39522
rect 5722 39520 5778 40000
rect 6550 39520 6606 40000
rect 7470 39520 7526 40000
rect 8390 39520 8446 40000
rect 9218 39520 9274 40000
rect 10138 39520 10194 40000
rect 11058 39520 11114 40000
rect 11886 39520 11942 40000
rect 12806 39520 12862 40000
rect 13726 39520 13782 40000
rect 14554 39520 14610 40000
rect 15474 39520 15530 40000
rect 400 35057 428 39520
rect 386 35048 442 35057
rect 386 34983 442 34992
rect 1228 34649 1256 39520
rect 1412 39494 2176 39520
rect 1214 34640 1270 34649
rect 1214 34575 1270 34584
rect 1412 19281 1440 39494
rect 3068 35601 3096 39520
rect 3896 37754 3924 39520
rect 4816 39494 5028 39520
rect 3896 37726 4016 37754
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3054 35592 3110 35601
rect 3054 35527 3110 35536
rect 3988 35193 4016 37726
rect 4066 37496 4122 37505
rect 4066 37431 4122 37440
rect 4080 37330 4108 37431
rect 4068 37324 4120 37330
rect 4068 37266 4120 37272
rect 3974 35184 4030 35193
rect 3974 35119 4030 35128
rect 4710 35048 4766 35057
rect 4710 34983 4766 34992
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 4158 34640 4214 34649
rect 4158 34575 4214 34584
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3240 28008 3292 28014
rect 3240 27950 3292 27956
rect 2872 26920 2924 26926
rect 2872 26862 2924 26868
rect 2688 25356 2740 25362
rect 2688 25298 2740 25304
rect 2700 25265 2728 25298
rect 2686 25256 2742 25265
rect 2686 25191 2742 25200
rect 2700 24954 2728 25191
rect 2688 24948 2740 24954
rect 2688 24890 2740 24896
rect 2884 22658 2912 26862
rect 3146 25800 3202 25809
rect 3146 25735 3202 25744
rect 3160 25430 3188 25735
rect 3148 25424 3200 25430
rect 2962 25392 3018 25401
rect 3148 25366 3200 25372
rect 2962 25327 2964 25336
rect 3016 25327 3018 25336
rect 2964 25298 3016 25304
rect 2976 24954 3004 25298
rect 2964 24948 3016 24954
rect 2964 24890 3016 24896
rect 2976 23186 3004 24890
rect 3146 24712 3202 24721
rect 3146 24647 3202 24656
rect 3056 24608 3108 24614
rect 3056 24550 3108 24556
rect 3068 24070 3096 24550
rect 3160 24274 3188 24647
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 3056 24064 3108 24070
rect 3056 24006 3108 24012
rect 2964 23180 3016 23186
rect 2964 23122 3016 23128
rect 2976 22778 3004 23122
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 2884 22630 3004 22658
rect 1398 19272 1454 19281
rect 1398 19207 1454 19216
rect 2870 19272 2926 19281
rect 2870 19207 2926 19216
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2778 19136 2834 19145
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 2056 18154 2084 18770
rect 2044 18148 2096 18154
rect 2044 18090 2096 18096
rect 1674 13968 1730 13977
rect 1674 13903 1730 13912
rect 386 8256 442 8265
rect 386 8191 442 8200
rect 400 480 428 8191
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1216 2984 1268 2990
rect 1216 2926 1268 2932
rect 1228 480 1256 2926
rect 1412 2553 1440 3878
rect 1688 2990 1716 13903
rect 2424 11218 2452 19110
rect 2778 19071 2834 19080
rect 2792 18970 2820 19071
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2792 18426 2820 18906
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2516 17542 2544 18158
rect 2884 18057 2912 19207
rect 2870 18048 2926 18057
rect 2870 17983 2926 17992
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2516 17105 2544 17478
rect 2502 17096 2558 17105
rect 2502 17031 2558 17040
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2516 14618 2544 14894
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2424 10470 2452 11154
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 9625 2452 10406
rect 2410 9616 2466 9625
rect 2410 9551 2466 9560
rect 2884 7528 2912 17983
rect 2976 13394 3004 22630
rect 3068 19242 3096 24006
rect 3160 23866 3188 24210
rect 3148 23860 3200 23866
rect 3148 23802 3200 23808
rect 3146 23760 3202 23769
rect 3146 23695 3202 23704
rect 3160 23594 3188 23695
rect 3148 23588 3200 23594
rect 3148 23530 3200 23536
rect 3252 19394 3280 27950
rect 4068 27872 4120 27878
rect 4068 27814 4120 27820
rect 3974 27432 4030 27441
rect 3974 27367 4030 27376
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3988 25945 4016 27367
rect 4080 27033 4108 27814
rect 4066 27024 4122 27033
rect 4066 26959 4122 26968
rect 4172 26926 4200 34575
rect 4724 33454 4752 34983
rect 4894 34776 4950 34785
rect 4894 34711 4950 34720
rect 4908 33658 4936 34711
rect 4896 33652 4948 33658
rect 4896 33594 4948 33600
rect 4712 33448 4764 33454
rect 4712 33390 4764 33396
rect 5000 29034 5028 39494
rect 5632 35624 5684 35630
rect 5632 35566 5684 35572
rect 5354 35048 5410 35057
rect 5354 34983 5410 34992
rect 5368 34202 5396 34983
rect 5540 34536 5592 34542
rect 5540 34478 5592 34484
rect 5356 34196 5408 34202
rect 5356 34138 5408 34144
rect 5264 34060 5316 34066
rect 5264 34002 5316 34008
rect 5276 33454 5304 34002
rect 5264 33448 5316 33454
rect 5262 33416 5264 33425
rect 5316 33416 5318 33425
rect 5262 33351 5318 33360
rect 5262 30424 5318 30433
rect 5262 30359 5318 30368
rect 5276 29170 5304 30359
rect 5356 29504 5408 29510
rect 5356 29446 5408 29452
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 5368 29073 5396 29446
rect 5354 29064 5410 29073
rect 4896 29028 4948 29034
rect 4896 28970 4948 28976
rect 4988 29028 5040 29034
rect 5354 28999 5356 29008
rect 4988 28970 5040 28976
rect 5408 28999 5410 29008
rect 5356 28970 5408 28976
rect 4908 28626 4936 28970
rect 4896 28620 4948 28626
rect 4896 28562 4948 28568
rect 4804 28416 4856 28422
rect 4804 28358 4856 28364
rect 4816 27674 4844 28358
rect 4908 27878 4936 28562
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5276 27946 5304 28358
rect 5368 28082 5396 28358
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 5264 27940 5316 27946
rect 5264 27882 5316 27888
rect 4896 27872 4948 27878
rect 4896 27814 4948 27820
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 4528 27532 4580 27538
rect 4528 27474 4580 27480
rect 4540 27441 4568 27474
rect 4526 27432 4582 27441
rect 4526 27367 4582 27376
rect 4540 27062 4568 27367
rect 4528 27056 4580 27062
rect 4528 26998 4580 27004
rect 4816 26994 4844 27610
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 4160 26920 4212 26926
rect 4160 26862 4212 26868
rect 4436 26784 4488 26790
rect 4436 26726 4488 26732
rect 4448 26450 4476 26726
rect 4620 26512 4672 26518
rect 4620 26454 4672 26460
rect 4436 26444 4488 26450
rect 4436 26386 4488 26392
rect 3974 25936 4030 25945
rect 3974 25871 4030 25880
rect 4632 25770 4660 26454
rect 4620 25764 4672 25770
rect 4620 25706 4672 25712
rect 3976 25696 4028 25702
rect 3976 25638 4028 25644
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3988 24614 4016 25638
rect 4632 25430 4660 25706
rect 4620 25424 4672 25430
rect 4620 25366 4672 25372
rect 4160 25220 4212 25226
rect 4160 25162 4212 25168
rect 4172 25106 4200 25162
rect 4080 25078 4200 25106
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 4080 23526 4108 25078
rect 4252 24744 4304 24750
rect 4252 24686 4304 24692
rect 4264 24274 4292 24686
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4264 24070 4292 24210
rect 4712 24200 4764 24206
rect 4342 24168 4398 24177
rect 4712 24142 4764 24148
rect 4342 24103 4398 24112
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 4264 23662 4292 24006
rect 4252 23656 4304 23662
rect 4252 23598 4304 23604
rect 3332 23520 3384 23526
rect 3332 23462 3384 23468
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 3344 22982 3372 23462
rect 3516 23112 3568 23118
rect 3516 23054 3568 23060
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3160 19366 3280 19394
rect 3056 19236 3108 19242
rect 3056 19178 3108 19184
rect 3160 18834 3188 19366
rect 3240 19304 3292 19310
rect 3238 19272 3240 19281
rect 3292 19272 3294 19281
rect 3238 19207 3294 19216
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3160 18426 3188 18770
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 3068 17270 3096 17682
rect 3056 17264 3108 17270
rect 3054 17232 3056 17241
rect 3108 17232 3110 17241
rect 3054 17167 3110 17176
rect 3160 14618 3188 18362
rect 3252 17814 3280 18566
rect 3344 17921 3372 22918
rect 3528 22778 3556 23054
rect 4264 22982 4292 23598
rect 4252 22976 4304 22982
rect 4252 22918 4304 22924
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 4066 22536 4122 22545
rect 4066 22471 4122 22480
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3804 21146 3832 21286
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3422 20360 3478 20369
rect 3988 20330 4016 20878
rect 3422 20295 3478 20304
rect 3976 20324 4028 20330
rect 3436 18970 3464 20295
rect 3976 20266 4028 20272
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 19961 3924 20198
rect 3882 19952 3938 19961
rect 3882 19887 3938 19896
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3436 18222 3464 18702
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3884 18216 3936 18222
rect 3988 18204 4016 20266
rect 4080 20074 4108 22471
rect 4264 21894 4292 22918
rect 4356 22574 4384 24103
rect 4724 23798 4752 24142
rect 4712 23792 4764 23798
rect 4712 23734 4764 23740
rect 4724 23526 4752 23734
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4344 22568 4396 22574
rect 4344 22510 4396 22516
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4448 21350 4476 22646
rect 4632 22642 4660 22918
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4632 22522 4660 22578
rect 4632 22494 4844 22522
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4344 21344 4396 21350
rect 4344 21286 4396 21292
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4250 20496 4306 20505
rect 4250 20431 4306 20440
rect 4264 20262 4292 20431
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4080 20058 4200 20074
rect 4080 20052 4212 20058
rect 4080 20046 4160 20052
rect 4160 19994 4212 20000
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4080 19310 4108 19858
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4172 18630 4200 19246
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4172 18290 4200 18566
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 3936 18176 4016 18204
rect 4264 18170 4292 20198
rect 3884 18158 3936 18164
rect 3330 17912 3386 17921
rect 3330 17847 3386 17856
rect 3240 17808 3292 17814
rect 3240 17750 3292 17756
rect 3238 17504 3294 17513
rect 3238 17439 3294 17448
rect 3252 16250 3280 17439
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2976 12986 3004 13330
rect 3344 12986 3372 17847
rect 3436 15094 3464 18158
rect 3896 17882 3924 18158
rect 4080 18142 4292 18170
rect 4080 18068 4108 18142
rect 3988 18040 4108 18068
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3436 13870 3464 15030
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3436 13462 3464 13806
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3436 13002 3464 13398
rect 3896 13297 3924 13670
rect 3882 13288 3938 13297
rect 3882 13223 3938 13232
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 2964 12980 3016 12986
rect 3332 12980 3384 12986
rect 3016 12940 3188 12968
rect 2964 12922 3016 12928
rect 3054 12472 3110 12481
rect 3054 12407 3056 12416
rect 3108 12407 3110 12416
rect 3056 12378 3108 12384
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3068 12209 3096 12242
rect 3054 12200 3110 12209
rect 3054 12135 3110 12144
rect 3068 11898 3096 12135
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2976 10810 3004 11154
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 3068 10418 3096 11018
rect 2608 7500 2912 7528
rect 2976 10390 3096 10418
rect 2608 6338 2636 7500
rect 2778 7440 2834 7449
rect 2778 7375 2834 7384
rect 2792 6474 2820 7375
rect 2976 6882 3004 10390
rect 3054 10296 3110 10305
rect 3054 10231 3110 10240
rect 3068 10130 3096 10231
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 3068 9382 3096 10066
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2700 6458 2820 6474
rect 2688 6452 2820 6458
rect 2740 6446 2820 6452
rect 2884 6854 3004 6882
rect 2688 6394 2740 6400
rect 2608 6310 2820 6338
rect 2504 6248 2556 6254
rect 2502 6216 2504 6225
rect 2556 6216 2558 6225
rect 2502 6151 2558 6160
rect 2516 5914 2544 6151
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2410 4992 2466 5001
rect 2410 4927 2466 4936
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 3777 2176 3878
rect 2134 3768 2190 3777
rect 2134 3703 2190 3712
rect 2240 3652 2268 4014
rect 2148 3624 2268 3652
rect 2318 3632 2374 3641
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1398 2544 1454 2553
rect 1398 2479 1454 2488
rect 2148 480 2176 3624
rect 2318 3567 2320 3576
rect 2372 3567 2374 3576
rect 2320 3538 2372 3544
rect 2332 3194 2360 3538
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2332 2689 2360 2790
rect 2318 2680 2374 2689
rect 2424 2650 2452 4927
rect 2792 4690 2820 6310
rect 2884 5137 2912 6854
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6458 3004 6666
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2870 5128 2926 5137
rect 2870 5063 2926 5072
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2608 3670 2636 4422
rect 2792 4282 2820 4626
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2504 3528 2556 3534
rect 2502 3496 2504 3505
rect 2556 3496 2558 3505
rect 2502 3431 2558 3440
rect 2608 3126 2636 3606
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2318 2615 2374 2624
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2700 2446 2728 3470
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2792 2922 2820 3334
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2884 2650 2912 5063
rect 2962 3768 3018 3777
rect 2962 3703 3018 3712
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2976 2446 3004 3703
rect 3068 3097 3096 9318
rect 3160 6905 3188 12940
rect 3436 12974 3556 13002
rect 3332 12922 3384 12928
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3238 9616 3294 9625
rect 3238 9551 3294 9560
rect 3146 6896 3202 6905
rect 3146 6831 3202 6840
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3160 3602 3188 6734
rect 3252 6458 3280 9551
rect 3344 9382 3372 12378
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 6730 3372 9318
rect 3436 7342 3464 12718
rect 3528 12442 3556 12974
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3988 11778 4016 18040
rect 4356 17898 4384 21286
rect 4448 21010 4476 21286
rect 4540 21146 4568 21966
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4632 21486 4660 21830
rect 4816 21554 4844 22494
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4620 21480 4672 21486
rect 4620 21422 4672 21428
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4632 21010 4660 21422
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4448 20262 4476 20946
rect 4908 20482 4936 27814
rect 5276 27674 5304 27882
rect 5264 27668 5316 27674
rect 5264 27610 5316 27616
rect 5276 26858 5304 27610
rect 5368 27606 5396 28018
rect 5356 27600 5408 27606
rect 5356 27542 5408 27548
rect 5356 27464 5408 27470
rect 5356 27406 5408 27412
rect 5368 27130 5396 27406
rect 5356 27124 5408 27130
rect 5356 27066 5408 27072
rect 5264 26852 5316 26858
rect 5264 26794 5316 26800
rect 5172 26784 5224 26790
rect 5172 26726 5224 26732
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4988 23248 5040 23254
rect 4988 23190 5040 23196
rect 5000 22778 5028 23190
rect 4988 22772 5040 22778
rect 4988 22714 5040 22720
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 5000 22506 5028 22578
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 5000 22166 5028 22442
rect 4988 22160 5040 22166
rect 4988 22102 5040 22108
rect 5000 21690 5028 22102
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 5092 21418 5120 23598
rect 5080 21412 5132 21418
rect 5080 21354 5132 21360
rect 4540 20454 4936 20482
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4448 18086 4476 18770
rect 4436 18080 4488 18086
rect 4434 18048 4436 18057
rect 4488 18048 4490 18057
rect 4434 17983 4490 17992
rect 4356 17870 4476 17898
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4172 17649 4200 17682
rect 4158 17640 4214 17649
rect 4158 17575 4214 17584
rect 4172 17338 4200 17575
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4448 16590 4476 17870
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4448 16114 4476 16526
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4160 15496 4212 15502
rect 4264 15473 4292 15982
rect 4160 15438 4212 15444
rect 4250 15464 4306 15473
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4080 14890 4108 15098
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4172 14414 4200 15438
rect 4250 15399 4306 15408
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4172 14074 4200 14350
rect 4264 14346 4292 15399
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4172 13818 4200 13874
rect 4080 13790 4200 13818
rect 4080 13530 4108 13790
rect 4356 13716 4384 14962
rect 4172 13688 4384 13716
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4172 12782 4200 13688
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4160 12776 4212 12782
rect 4080 12736 4160 12764
rect 4080 12442 4108 12736
rect 4160 12718 4212 12724
rect 4264 12442 4292 13194
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4356 12850 4384 13126
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 3896 11750 4016 11778
rect 3896 11082 3924 11750
rect 4080 11694 4108 12378
rect 4068 11688 4120 11694
rect 3974 11656 4030 11665
rect 4068 11630 4120 11636
rect 3974 11591 4030 11600
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3882 10704 3938 10713
rect 3882 10639 3938 10648
rect 3896 10470 3924 10639
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3896 10010 3924 10406
rect 3988 10266 4016 11591
rect 4080 11354 4108 11630
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10810 4108 10950
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4172 10674 4200 11154
rect 4264 11150 4292 11562
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4356 10810 4384 11222
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4172 10266 4200 10610
rect 4356 10538 4384 10746
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4068 10056 4120 10062
rect 3896 9982 4016 10010
rect 4068 9998 4120 10004
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3528 7342 3556 8026
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3988 7478 4016 9982
rect 4080 9654 4108 9998
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4448 8634 4476 16050
rect 4540 10305 4568 20454
rect 4804 20324 4856 20330
rect 4804 20266 4856 20272
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4632 17202 4660 20198
rect 4816 19990 4844 20266
rect 4908 20058 4936 20266
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 4908 19514 4936 19994
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4908 18222 4936 18566
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4816 17785 4844 17818
rect 4802 17776 4858 17785
rect 4802 17711 4858 17720
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4724 17134 4752 17478
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4724 16658 4752 17070
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4724 15706 4752 16594
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4724 15094 4752 15642
rect 4816 15570 4844 16526
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4908 15450 4936 18158
rect 5078 17912 5134 17921
rect 5078 17847 5134 17856
rect 5092 17746 5120 17847
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5092 17338 5120 17682
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 5000 16794 5028 17002
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5000 16114 5028 16730
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 4816 15422 4936 15450
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4632 14550 4660 14758
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4632 13530 4660 14486
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4724 13394 4752 14010
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4724 12646 4752 13330
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4618 12336 4674 12345
rect 4618 12271 4674 12280
rect 4632 11762 4660 12271
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4526 10296 4582 10305
rect 4526 10231 4582 10240
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4540 9994 4568 10066
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4540 9722 4568 9930
rect 4632 9897 4660 11698
rect 4724 10742 4752 12582
rect 4816 12481 4844 15422
rect 5092 15314 5120 17138
rect 4908 15286 5120 15314
rect 4802 12472 4858 12481
rect 4802 12407 4858 12416
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4816 11082 4844 12174
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4724 10198 4752 10474
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4618 9888 4674 9897
rect 4618 9823 4674 9832
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4264 8090 4292 8366
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3252 6254 3280 6394
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3436 5794 3464 7103
rect 3528 7002 3556 7278
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3528 5914 3556 6258
rect 3988 6254 4016 6938
rect 4080 6882 4108 7210
rect 4264 7206 4292 7822
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4080 6854 4200 6882
rect 4172 6662 4200 6854
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 4264 6202 4292 7142
rect 4356 6866 4384 8298
rect 4540 8265 4568 9658
rect 4632 9110 4660 9823
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4632 8566 4660 9046
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4724 8430 4752 8978
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4526 8256 4582 8265
rect 4526 8191 4582 8200
rect 4816 8090 4844 8910
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4434 7984 4490 7993
rect 4434 7919 4490 7928
rect 4448 7410 4476 7919
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 6322 4384 6802
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3436 5766 3556 5794
rect 3238 4720 3294 4729
rect 3238 4655 3294 4664
rect 3252 4214 3280 4655
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3238 3632 3294 3641
rect 3148 3596 3200 3602
rect 3238 3567 3294 3576
rect 3148 3538 3200 3544
rect 3054 3088 3110 3097
rect 3054 3023 3110 3032
rect 3252 2961 3280 3567
rect 3344 3058 3372 3839
rect 3436 3641 3464 4218
rect 3422 3632 3478 3641
rect 3422 3567 3478 3576
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3528 2990 3556 5766
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3988 5166 4016 6190
rect 4160 6180 4212 6186
rect 4264 6174 4384 6202
rect 4160 6122 4212 6128
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5302 4108 5510
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3988 4826 4016 5102
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3790 4176 3846 4185
rect 3790 4111 3846 4120
rect 3698 4040 3754 4049
rect 3804 4010 3832 4111
rect 3698 3975 3700 3984
rect 3752 3975 3754 3984
rect 3792 4004 3844 4010
rect 3700 3946 3752 3952
rect 3792 3946 3844 3952
rect 3804 3738 3832 3946
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 4172 3058 4200 6122
rect 4356 5778 4384 6174
rect 4448 5846 4476 7346
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6458 4568 6734
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5302 4384 5714
rect 4448 5370 4476 5782
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4356 4826 4384 5238
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4356 3777 4384 3946
rect 4342 3768 4398 3777
rect 4342 3703 4398 3712
rect 4448 3670 4476 4218
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 3516 2984 3568 2990
rect 3238 2952 3294 2961
rect 3056 2916 3108 2922
rect 3516 2926 3568 2932
rect 3238 2887 3294 2896
rect 3056 2858 3108 2864
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3068 480 3096 2858
rect 4172 2650 4200 2994
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4068 2576 4120 2582
rect 4264 2530 4292 3334
rect 4448 2922 4476 3606
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2650 4384 2790
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4120 2524 4292 2530
rect 4068 2518 4292 2524
rect 4080 2502 4292 2518
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 4632 2038 4660 7414
rect 4816 7410 4844 8026
rect 4908 7954 4936 15286
rect 5092 15201 5120 15286
rect 5078 15192 5134 15201
rect 5078 15127 5134 15136
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 5000 13870 5028 14282
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 5184 13705 5212 26726
rect 5276 26042 5304 26794
rect 5368 26518 5396 27066
rect 5552 27062 5580 34478
rect 5644 28150 5672 35566
rect 5632 28144 5684 28150
rect 5632 28086 5684 28092
rect 5736 28098 5764 39520
rect 6564 37754 6592 39520
rect 6564 37726 6868 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6000 37324 6052 37330
rect 6000 37266 6052 37272
rect 6012 35290 6040 37266
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6000 35284 6052 35290
rect 6000 35226 6052 35232
rect 5998 35184 6054 35193
rect 5998 35119 6054 35128
rect 6736 35148 6788 35154
rect 5816 34672 5868 34678
rect 5814 34640 5816 34649
rect 5868 34640 5870 34649
rect 5814 34575 5870 34584
rect 6012 32978 6040 35119
rect 6736 35090 6788 35096
rect 6748 34542 6776 35090
rect 6840 34626 6868 37726
rect 7484 36242 7512 39520
rect 7472 36236 7524 36242
rect 7472 36178 7524 36184
rect 7484 35834 7512 36178
rect 8300 36100 8352 36106
rect 8300 36042 8352 36048
rect 7472 35828 7524 35834
rect 7472 35770 7524 35776
rect 7012 35760 7064 35766
rect 7010 35728 7012 35737
rect 7064 35728 7066 35737
rect 7010 35663 7066 35672
rect 7484 35193 7512 35770
rect 8312 35562 8340 36042
rect 8300 35556 8352 35562
rect 8300 35498 8352 35504
rect 8312 35290 8340 35498
rect 8300 35284 8352 35290
rect 8300 35226 8352 35232
rect 7470 35184 7526 35193
rect 7288 35148 7340 35154
rect 7470 35119 7526 35128
rect 7288 35090 7340 35096
rect 6840 34598 6960 34626
rect 6736 34536 6788 34542
rect 6736 34478 6788 34484
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6368 34128 6420 34134
rect 6368 34070 6420 34076
rect 6184 33924 6236 33930
rect 6184 33866 6236 33872
rect 6092 33380 6144 33386
rect 6092 33322 6144 33328
rect 6000 32972 6052 32978
rect 6000 32914 6052 32920
rect 6012 32230 6040 32914
rect 6000 32224 6052 32230
rect 6000 32166 6052 32172
rect 5814 31920 5870 31929
rect 5814 31855 5816 31864
rect 5868 31855 5870 31864
rect 5816 31826 5868 31832
rect 5828 31482 5856 31826
rect 5816 31476 5868 31482
rect 5816 31418 5868 31424
rect 5828 28234 5856 31418
rect 5906 30696 5962 30705
rect 5906 30631 5962 30640
rect 5920 29170 5948 30631
rect 5908 29164 5960 29170
rect 5908 29106 5960 29112
rect 5828 28206 5948 28234
rect 5736 28070 5856 28098
rect 5724 27940 5776 27946
rect 5724 27882 5776 27888
rect 5632 27600 5684 27606
rect 5632 27542 5684 27548
rect 5540 27056 5592 27062
rect 5540 26998 5592 27004
rect 5644 26586 5672 27542
rect 5736 27470 5764 27882
rect 5724 27464 5776 27470
rect 5724 27406 5776 27412
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5356 26512 5408 26518
rect 5356 26454 5408 26460
rect 5448 26376 5500 26382
rect 5736 26330 5764 27406
rect 5828 27169 5856 28070
rect 5814 27160 5870 27169
rect 5814 27095 5870 27104
rect 5448 26318 5500 26324
rect 5264 26036 5316 26042
rect 5264 25978 5316 25984
rect 5460 25684 5488 26318
rect 5644 26314 5764 26330
rect 5632 26308 5764 26314
rect 5684 26302 5764 26308
rect 5632 26250 5684 26256
rect 5540 25696 5592 25702
rect 5460 25656 5540 25684
rect 5264 25424 5316 25430
rect 5264 25366 5316 25372
rect 5276 24614 5304 25366
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 5460 24342 5488 25656
rect 5540 25638 5592 25644
rect 5540 24744 5592 24750
rect 5540 24686 5592 24692
rect 5448 24336 5500 24342
rect 5448 24278 5500 24284
rect 5448 24132 5500 24138
rect 5448 24074 5500 24080
rect 5460 23662 5488 24074
rect 5552 24070 5580 24686
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5552 23662 5580 24006
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 5276 18630 5304 23462
rect 5448 23044 5500 23050
rect 5448 22986 5500 22992
rect 5460 22953 5488 22986
rect 5446 22944 5502 22953
rect 5368 22902 5446 22930
rect 5368 20534 5396 22902
rect 5446 22879 5502 22888
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5460 22234 5488 22714
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5552 22030 5580 23598
rect 5644 23118 5672 26250
rect 5828 24698 5856 27095
rect 5920 25401 5948 28206
rect 6012 27334 6040 32166
rect 6000 27328 6052 27334
rect 6104 27305 6132 33322
rect 6196 33114 6224 33866
rect 6380 33658 6408 34070
rect 6368 33652 6420 33658
rect 6368 33594 6420 33600
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6184 33108 6236 33114
rect 6184 33050 6236 33056
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6644 31884 6696 31890
rect 6644 31826 6696 31832
rect 6656 31142 6684 31826
rect 6644 31136 6696 31142
rect 6644 31078 6696 31084
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6656 30054 6684 31078
rect 6748 30705 6776 34478
rect 6828 32360 6880 32366
rect 6828 32302 6880 32308
rect 6840 31958 6868 32302
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6932 31793 6960 34598
rect 7300 34406 7328 35090
rect 8116 35080 8168 35086
rect 8114 35048 8116 35057
rect 8168 35048 8170 35057
rect 8404 35034 8432 39520
rect 9232 37210 9260 39520
rect 9232 37182 9352 37210
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 9324 36378 9352 37182
rect 9956 36576 10008 36582
rect 9956 36518 10008 36524
rect 9312 36372 9364 36378
rect 9312 36314 9364 36320
rect 8576 36304 8628 36310
rect 8576 36246 8628 36252
rect 8588 35562 8616 36246
rect 9588 36236 9640 36242
rect 9588 36178 9640 36184
rect 9772 36236 9824 36242
rect 9772 36178 9824 36184
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 9600 35834 9628 36178
rect 9588 35828 9640 35834
rect 9588 35770 9640 35776
rect 8760 35692 8812 35698
rect 8760 35634 8812 35640
rect 8576 35556 8628 35562
rect 8576 35498 8628 35504
rect 8588 35222 8616 35498
rect 8576 35216 8628 35222
rect 8576 35158 8628 35164
rect 8220 35018 8432 35034
rect 8114 34983 8170 34992
rect 8208 35012 8432 35018
rect 7564 34944 7616 34950
rect 7564 34886 7616 34892
rect 8024 34944 8076 34950
rect 8024 34886 8076 34892
rect 7576 34785 7604 34886
rect 7562 34776 7618 34785
rect 7562 34711 7618 34720
rect 7576 34678 7604 34711
rect 7564 34672 7616 34678
rect 7564 34614 7616 34620
rect 8036 34610 8064 34886
rect 8128 34746 8156 34983
rect 8260 35006 8432 35012
rect 8208 34954 8260 34960
rect 8116 34740 8168 34746
rect 8116 34682 8168 34688
rect 8024 34604 8076 34610
rect 8024 34546 8076 34552
rect 7932 34468 7984 34474
rect 7932 34410 7984 34416
rect 7288 34400 7340 34406
rect 7288 34342 7340 34348
rect 7300 33318 7328 34342
rect 7944 34134 7972 34410
rect 7932 34128 7984 34134
rect 7932 34070 7984 34076
rect 7564 33856 7616 33862
rect 7564 33798 7616 33804
rect 7576 33522 7604 33798
rect 7564 33516 7616 33522
rect 7564 33458 7616 33464
rect 7656 33380 7708 33386
rect 7656 33322 7708 33328
rect 7288 33312 7340 33318
rect 7288 33254 7340 33260
rect 7196 33040 7248 33046
rect 7196 32982 7248 32988
rect 7208 32298 7236 32982
rect 7196 32292 7248 32298
rect 7196 32234 7248 32240
rect 6918 31784 6974 31793
rect 6918 31719 6974 31728
rect 7300 31634 7328 33254
rect 7668 33114 7696 33322
rect 7944 33114 7972 34070
rect 8036 33522 8064 34546
rect 8588 34524 8616 35158
rect 8668 34536 8720 34542
rect 8588 34496 8668 34524
rect 8668 34478 8720 34484
rect 8300 33992 8352 33998
rect 8300 33934 8352 33940
rect 8024 33516 8076 33522
rect 8024 33458 8076 33464
rect 7656 33108 7708 33114
rect 7656 33050 7708 33056
rect 7932 33108 7984 33114
rect 7932 33050 7984 33056
rect 7472 32904 7524 32910
rect 7472 32846 7524 32852
rect 7116 31606 7328 31634
rect 7380 31680 7432 31686
rect 7484 31668 7512 32846
rect 7944 32570 7972 33050
rect 7932 32564 7984 32570
rect 7932 32506 7984 32512
rect 8036 32450 8064 33458
rect 8312 33114 8340 33934
rect 8300 33108 8352 33114
rect 8300 33050 8352 33056
rect 8576 32972 8628 32978
rect 8576 32914 8628 32920
rect 8588 32570 8616 32914
rect 8680 32570 8708 34478
rect 8772 33998 8800 35634
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8760 33992 8812 33998
rect 8760 33934 8812 33940
rect 8760 32768 8812 32774
rect 8760 32710 8812 32716
rect 8576 32564 8628 32570
rect 8576 32506 8628 32512
rect 8668 32564 8720 32570
rect 8668 32506 8720 32512
rect 7944 32422 8064 32450
rect 8482 32464 8538 32473
rect 7748 31816 7800 31822
rect 7748 31758 7800 31764
rect 7432 31640 7512 31668
rect 7380 31622 7432 31628
rect 6920 31272 6972 31278
rect 6920 31214 6972 31220
rect 6734 30696 6790 30705
rect 6734 30631 6790 30640
rect 6932 30598 6960 31214
rect 7012 30728 7064 30734
rect 7012 30670 7064 30676
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 7024 30433 7052 30670
rect 7010 30424 7066 30433
rect 7010 30359 7066 30368
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6656 29714 6684 29990
rect 6644 29708 6696 29714
rect 6644 29650 6696 29656
rect 6656 29102 6684 29650
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 6644 29096 6696 29102
rect 6644 29038 6696 29044
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6366 28656 6422 28665
rect 6656 28626 6684 29038
rect 6366 28591 6368 28600
rect 6420 28591 6422 28600
rect 6644 28620 6696 28626
rect 6368 28562 6420 28568
rect 6644 28562 6696 28568
rect 6380 27962 6408 28562
rect 6656 28218 6684 28562
rect 6748 28422 6776 29582
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 6736 28416 6788 28422
rect 6736 28358 6788 28364
rect 6644 28212 6696 28218
rect 6644 28154 6696 28160
rect 6840 28082 6868 28494
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6196 27934 6408 27962
rect 6196 27674 6224 27934
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6840 27674 6868 28018
rect 6184 27668 6236 27674
rect 6184 27610 6236 27616
rect 6828 27668 6880 27674
rect 6828 27610 6880 27616
rect 6000 27270 6052 27276
rect 6090 27296 6146 27305
rect 6090 27231 6146 27240
rect 6196 27010 6224 27610
rect 7116 27606 7144 31606
rect 7392 31346 7420 31622
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7760 30938 7788 31758
rect 7748 30932 7800 30938
rect 7748 30874 7800 30880
rect 7944 30734 7972 32422
rect 8772 32434 8800 32710
rect 8482 32399 8538 32408
rect 8760 32428 8812 32434
rect 8116 31884 8168 31890
rect 8116 31826 8168 31832
rect 8022 31784 8078 31793
rect 8022 31719 8078 31728
rect 7932 30728 7984 30734
rect 7932 30670 7984 30676
rect 7472 30184 7524 30190
rect 7472 30126 7524 30132
rect 7484 29850 7512 30126
rect 7564 30048 7616 30054
rect 7564 29990 7616 29996
rect 7472 29844 7524 29850
rect 7472 29786 7524 29792
rect 7196 29640 7248 29646
rect 7196 29582 7248 29588
rect 7208 29170 7236 29582
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 7208 28762 7236 29106
rect 7196 28756 7248 28762
rect 7196 28698 7248 28704
rect 7576 28626 7604 29990
rect 7944 29850 7972 30670
rect 7932 29844 7984 29850
rect 7932 29786 7984 29792
rect 7932 29096 7984 29102
rect 7746 29064 7802 29073
rect 7746 28999 7802 29008
rect 7930 29064 7932 29073
rect 7984 29064 7986 29073
rect 7930 28999 7986 29008
rect 7564 28620 7616 28626
rect 7564 28562 7616 28568
rect 7576 28218 7604 28562
rect 7564 28212 7616 28218
rect 7564 28154 7616 28160
rect 7760 28150 7788 28999
rect 7748 28144 7800 28150
rect 7748 28086 7800 28092
rect 7932 27940 7984 27946
rect 7932 27882 7984 27888
rect 6276 27600 6328 27606
rect 6276 27542 6328 27548
rect 7104 27600 7156 27606
rect 7380 27600 7432 27606
rect 7104 27542 7156 27548
rect 7378 27568 7380 27577
rect 7432 27568 7434 27577
rect 6288 27130 6316 27542
rect 7378 27503 7434 27512
rect 7392 27452 7420 27503
rect 7840 27464 7892 27470
rect 7194 27432 7250 27441
rect 7012 27396 7064 27402
rect 7392 27424 7512 27452
rect 7194 27367 7250 27376
rect 7012 27338 7064 27344
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6276 27124 6328 27130
rect 6276 27066 6328 27072
rect 6012 26982 6224 27010
rect 5906 25392 5962 25401
rect 5906 25327 5962 25336
rect 5908 25152 5960 25158
rect 5908 25094 5960 25100
rect 5920 24818 5948 25094
rect 6012 24818 6040 26982
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 6196 26518 6224 26862
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6184 26512 6236 26518
rect 6104 26472 6184 26500
rect 6104 25702 6132 26472
rect 6184 26454 6236 26460
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6472 26042 6500 26318
rect 6460 26036 6512 26042
rect 6460 25978 6512 25984
rect 6092 25696 6144 25702
rect 6092 25638 6144 25644
rect 6104 25498 6132 25638
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6092 25492 6144 25498
rect 6092 25434 6144 25440
rect 6656 24993 6684 27270
rect 6918 27024 6974 27033
rect 7024 26994 7052 27338
rect 6918 26959 6920 26968
rect 6972 26959 6974 26968
rect 7012 26988 7064 26994
rect 6920 26930 6972 26936
rect 7012 26930 7064 26936
rect 6932 26586 6960 26930
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6920 25968 6972 25974
rect 6918 25936 6920 25945
rect 6972 25936 6974 25945
rect 6918 25871 6974 25880
rect 7024 25786 7052 26930
rect 6932 25758 7052 25786
rect 6642 24984 6698 24993
rect 6642 24919 6698 24928
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 6000 24812 6052 24818
rect 6000 24754 6052 24760
rect 5828 24670 6224 24698
rect 5908 23588 5960 23594
rect 5908 23530 5960 23536
rect 5920 23322 5948 23530
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 5632 23112 5684 23118
rect 5632 23054 5684 23060
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5356 20528 5408 20534
rect 5356 20470 5408 20476
rect 5368 19922 5396 20470
rect 5460 20074 5488 21626
rect 6012 21350 6040 22034
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5460 20046 5580 20074
rect 5552 19990 5580 20046
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5552 19310 5580 19790
rect 5540 19304 5592 19310
rect 5644 19281 5672 21082
rect 6196 20505 6224 24670
rect 6644 24608 6696 24614
rect 6644 24550 6696 24556
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6276 24268 6328 24274
rect 6276 24210 6328 24216
rect 6288 23662 6316 24210
rect 6656 23866 6684 24550
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6276 23656 6328 23662
rect 6274 23624 6276 23633
rect 6328 23624 6330 23633
rect 6656 23594 6684 23802
rect 6840 23662 6868 24006
rect 6828 23656 6880 23662
rect 6828 23598 6880 23604
rect 6274 23559 6330 23568
rect 6644 23588 6696 23594
rect 6644 23530 6696 23536
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6656 23254 6684 23530
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 6656 22778 6684 23190
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6840 22234 6868 23598
rect 6932 22506 6960 25758
rect 7104 25424 7156 25430
rect 7104 25366 7156 25372
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7024 23186 7052 24754
rect 7116 24614 7144 25366
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7208 23202 7236 27367
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7300 24682 7328 25094
rect 7288 24676 7340 24682
rect 7288 24618 7340 24624
rect 7288 24336 7340 24342
rect 7288 24278 7340 24284
rect 7300 23322 7328 24278
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 7012 23180 7064 23186
rect 7208 23174 7328 23202
rect 7012 23122 7064 23128
rect 7194 22944 7250 22953
rect 7194 22879 7250 22888
rect 7208 22642 7236 22879
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7194 22536 7250 22545
rect 6920 22500 6972 22506
rect 7194 22471 7250 22480
rect 6920 22442 6972 22448
rect 6932 22234 6960 22442
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6748 21321 6776 21422
rect 6734 21312 6790 21321
rect 6289 21244 6585 21264
rect 6734 21247 6790 21256
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6840 21146 6868 22034
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6932 21622 6960 21966
rect 6920 21616 6972 21622
rect 6920 21558 6972 21564
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6288 20602 6316 20878
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 6182 20496 6238 20505
rect 6182 20431 6238 20440
rect 6656 20262 6684 21014
rect 7208 20874 7236 22471
rect 7196 20868 7248 20874
rect 7196 20810 7248 20816
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 20369 6960 20742
rect 6918 20360 6974 20369
rect 6918 20295 6920 20304
rect 6972 20295 6974 20304
rect 7012 20324 7064 20330
rect 6920 20266 6972 20272
rect 7012 20266 7064 20272
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6656 19990 6684 20198
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 5736 19514 5764 19926
rect 7024 19802 7052 20266
rect 7194 19952 7250 19961
rect 7194 19887 7250 19896
rect 7208 19854 7236 19887
rect 6932 19774 7052 19802
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 6932 19718 6960 19774
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5540 19246 5592 19252
rect 5630 19272 5686 19281
rect 5736 19242 5764 19450
rect 5998 19272 6054 19281
rect 5630 19207 5686 19216
rect 5724 19236 5776 19242
rect 5644 18816 5672 19207
rect 5998 19207 6054 19216
rect 5724 19178 5776 19184
rect 5736 18902 5764 19178
rect 5724 18896 5776 18902
rect 5776 18844 5856 18850
rect 5724 18838 5856 18844
rect 5736 18822 5856 18838
rect 5552 18788 5672 18816
rect 5552 18630 5580 18788
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5632 18692 5684 18698
rect 5632 18634 5684 18640
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5276 16250 5304 18362
rect 5552 18222 5580 18566
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5368 17513 5396 18090
rect 5552 17746 5580 18158
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5354 17504 5410 17513
rect 5354 17439 5410 17448
rect 5552 17338 5580 17682
rect 5644 17678 5672 18634
rect 5736 18154 5764 18702
rect 5828 18426 5856 18822
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5724 18148 5776 18154
rect 5724 18090 5776 18096
rect 5736 17882 5764 18090
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5828 17814 5856 18158
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5644 16794 5672 17614
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5276 15978 5304 16186
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5276 15638 5304 15914
rect 5908 15904 5960 15910
rect 5908 15846 5960 15852
rect 5920 15638 5948 15846
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5908 15632 5960 15638
rect 5908 15574 5960 15580
rect 5276 15162 5304 15574
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 15162 5580 15506
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5276 14929 5304 15098
rect 5262 14920 5318 14929
rect 5262 14855 5318 14864
rect 5170 13696 5226 13705
rect 5170 13631 5226 13640
rect 5276 13462 5304 14855
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 13938 5580 14214
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 4988 13252 5040 13258
rect 4988 13194 5040 13200
rect 5000 12850 5028 13194
rect 5276 13002 5304 13398
rect 5184 12974 5304 13002
rect 5184 12918 5212 12974
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 5000 11898 5028 12310
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11354 5120 11494
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5184 11218 5212 12854
rect 5644 12850 5672 15302
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5828 14278 5856 14826
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 14006 5856 14214
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12238 5672 12786
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5276 11665 5304 11698
rect 5262 11656 5318 11665
rect 5262 11591 5318 11600
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5448 11144 5500 11150
rect 5500 11092 5580 11098
rect 5448 11086 5580 11092
rect 5460 11070 5580 11086
rect 5552 10810 5580 11070
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10198 5396 10406
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5080 9512 5132 9518
rect 5078 9480 5080 9489
rect 5132 9480 5134 9489
rect 5368 9450 5396 10134
rect 5644 10062 5672 12174
rect 5828 11626 5856 13942
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5078 9415 5134 9424
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5368 9178 5396 9386
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8430 5396 8774
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5368 7954 5396 8366
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4908 7002 4936 7890
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4710 6896 4766 6905
rect 4710 6831 4766 6840
rect 4724 5522 4752 6831
rect 4804 5704 4856 5710
rect 4802 5672 4804 5681
rect 4856 5672 4858 5681
rect 4802 5607 4858 5616
rect 4908 5574 4936 6938
rect 5092 6934 5120 7210
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5080 6928 5132 6934
rect 4986 6896 5042 6905
rect 5080 6870 5132 6876
rect 4986 6831 5042 6840
rect 5000 6798 5028 6831
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5092 6390 5120 6870
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 4896 5568 4948 5574
rect 4724 5494 4844 5522
rect 4896 5510 4948 5516
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4724 4622 4752 5034
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4214 4752 4558
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 3884 2032 3936 2038
rect 3884 1974 3936 1980
rect 4620 2032 4672 2038
rect 4620 1974 4672 1980
rect 3896 480 3924 1974
rect 4816 480 4844 5494
rect 5184 3233 5212 6938
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 6458 5304 6598
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5460 6361 5488 7822
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5446 6352 5502 6361
rect 5446 6287 5502 6296
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5368 5914 5396 6122
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5276 5001 5304 5034
rect 5262 4992 5318 5001
rect 5262 4927 5318 4936
rect 5276 4826 5304 4927
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5368 4758 5396 5850
rect 5552 5114 5580 7142
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5460 5098 5580 5114
rect 5448 5092 5580 5098
rect 5500 5086 5580 5092
rect 5448 5034 5500 5040
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5368 4282 5396 4694
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5276 3738 5304 4082
rect 5460 4010 5488 5034
rect 5644 4570 5672 5578
rect 5552 4542 5672 4570
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5460 3670 5488 3946
rect 5552 3942 5580 4542
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5644 4185 5672 4422
rect 5630 4176 5686 4185
rect 5630 4111 5686 4120
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5170 3224 5226 3233
rect 5276 3194 5304 3538
rect 5736 3369 5764 10406
rect 5828 9654 5856 11562
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5920 7002 5948 14554
rect 6012 14074 6040 19207
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6196 17746 6224 18702
rect 6656 18358 6684 19110
rect 6932 18902 6960 19654
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 7024 19258 7052 19314
rect 7024 19242 7144 19258
rect 7024 19236 7156 19242
rect 7024 19230 7104 19236
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6656 17882 6684 18294
rect 6840 18222 6868 18566
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 7024 17785 7052 19230
rect 7104 19178 7156 19184
rect 7010 17776 7066 17785
rect 6184 17740 6236 17746
rect 7010 17711 7066 17720
rect 6184 17682 6236 17688
rect 6918 17232 6974 17241
rect 6918 17167 6920 17176
rect 6972 17167 6974 17176
rect 6920 17138 6972 17144
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 7208 16833 7236 17070
rect 7194 16824 7250 16833
rect 7194 16759 7196 16768
rect 7248 16759 7250 16768
rect 7196 16730 7248 16736
rect 6642 16688 6698 16697
rect 6092 16652 6144 16658
rect 6642 16623 6698 16632
rect 6092 16594 6144 16600
rect 6104 16250 6132 16594
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6472 15366 6500 15438
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6564 15162 6592 15574
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6656 15094 6684 16623
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 6920 15496 6972 15502
rect 6918 15464 6920 15473
rect 6972 15464 6974 15473
rect 6828 15428 6880 15434
rect 6918 15399 6974 15408
rect 6828 15370 6880 15376
rect 6644 15088 6696 15094
rect 6644 15030 6696 15036
rect 6734 15056 6790 15065
rect 6734 14991 6790 15000
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6748 14482 6776 14991
rect 6840 14822 6868 15370
rect 6932 15026 6960 15399
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14618 6868 14758
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6380 14074 6408 14418
rect 7024 14362 7052 15302
rect 6840 14346 7052 14362
rect 6828 14340 7052 14346
rect 6880 14334 7052 14340
rect 6828 14282 6880 14288
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 7116 13938 7144 15846
rect 7300 13977 7328 23174
rect 7380 22976 7432 22982
rect 7380 22918 7432 22924
rect 7392 22506 7420 22918
rect 7380 22500 7432 22506
rect 7380 22442 7432 22448
rect 7380 20868 7432 20874
rect 7380 20810 7432 20816
rect 7392 20466 7420 20810
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 7392 17814 7420 20402
rect 7380 17808 7432 17814
rect 7380 17750 7432 17756
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7392 15366 7420 15982
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7286 13968 7342 13977
rect 7104 13932 7156 13938
rect 7286 13903 7342 13912
rect 7104 13874 7156 13880
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6090 13696 6146 13705
rect 6012 13190 6040 13670
rect 6090 13631 6146 13640
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6012 12646 6040 13126
rect 6104 12889 6132 13631
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6828 13320 6880 13326
rect 6182 13288 6238 13297
rect 6828 13262 6880 13268
rect 6182 13223 6238 13232
rect 6196 12986 6224 13223
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6090 12880 6146 12889
rect 6090 12815 6146 12824
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 12442 6040 12582
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5920 5846 5948 6054
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5906 4040 5962 4049
rect 5906 3975 5908 3984
rect 5960 3975 5962 3984
rect 5908 3946 5960 3952
rect 6012 3670 6040 6598
rect 6104 6202 6132 12815
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6840 12238 6868 13262
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6840 11898 6868 12174
rect 7024 11898 7052 12310
rect 7102 12200 7158 12209
rect 7102 12135 7104 12144
rect 7156 12135 7158 12144
rect 7104 12106 7156 12112
rect 7392 11898 7420 12650
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7010 11792 7066 11801
rect 7010 11727 7066 11736
rect 6182 11656 6238 11665
rect 6182 11591 6238 11600
rect 6196 11218 6224 11591
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 10470 6224 11154
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6840 10146 6868 11018
rect 6840 10118 6960 10146
rect 6932 10062 6960 10118
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6550 9616 6606 9625
rect 6550 9551 6552 9560
rect 6604 9551 6606 9560
rect 6552 9522 6604 9528
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 8430 6224 8978
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 7993 6224 8366
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6656 8022 6684 8230
rect 6644 8016 6696 8022
rect 6182 7984 6238 7993
rect 6644 7958 6696 7964
rect 6182 7919 6238 7928
rect 6656 7546 6684 7958
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6748 6882 6776 8298
rect 6840 7886 6868 9998
rect 7024 7970 7052 11727
rect 7392 11626 7420 11834
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7392 11286 7420 11562
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7116 9042 7144 9386
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7024 7942 7144 7970
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6840 7478 6868 7822
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6748 6866 6960 6882
rect 6748 6860 6972 6866
rect 6748 6854 6920 6860
rect 6920 6802 6972 6808
rect 7024 6225 7052 7822
rect 7010 6216 7066 6225
rect 6104 6174 6684 6202
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6104 5098 6132 5646
rect 6196 5370 6224 5782
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6104 4486 6132 5034
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 3913 6132 4422
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6090 3904 6146 3913
rect 6090 3839 6146 3848
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 5908 3528 5960 3534
rect 5906 3496 5908 3505
rect 5960 3496 5962 3505
rect 5906 3431 5962 3440
rect 5722 3360 5778 3369
rect 5722 3295 5778 3304
rect 5170 3159 5226 3168
rect 5264 3188 5316 3194
rect 4986 2680 5042 2689
rect 4986 2615 5042 2624
rect 5000 2582 5028 2615
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 5000 2446 5028 2518
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5184 610 5212 3159
rect 5264 3130 5316 3136
rect 5920 3058 5948 3431
rect 6012 3194 6040 3606
rect 6196 3534 6224 3946
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6184 3528 6236 3534
rect 6656 3505 6684 6174
rect 7010 6151 7066 6160
rect 7116 5817 7144 7942
rect 7102 5808 7158 5817
rect 7208 5778 7236 9454
rect 7300 9110 7328 11086
rect 7392 10810 7420 11222
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7392 10538 7420 10746
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7392 10266 7420 10474
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7392 8362 7420 10202
rect 7484 9994 7512 27424
rect 7840 27406 7892 27412
rect 7852 27130 7880 27406
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7564 26444 7616 26450
rect 7564 26386 7616 26392
rect 7576 25702 7604 26386
rect 7656 26240 7708 26246
rect 7656 26182 7708 26188
rect 7668 25838 7696 26182
rect 7944 25974 7972 27882
rect 8036 26874 8064 31719
rect 8128 31142 8156 31826
rect 8300 31272 8352 31278
rect 8300 31214 8352 31220
rect 8116 31136 8168 31142
rect 8116 31078 8168 31084
rect 8208 30864 8260 30870
rect 8208 30806 8260 30812
rect 8220 30410 8248 30806
rect 8312 30546 8340 31214
rect 8392 30728 8444 30734
rect 8390 30696 8392 30705
rect 8444 30696 8446 30705
rect 8390 30631 8446 30640
rect 8392 30592 8444 30598
rect 8312 30540 8392 30546
rect 8312 30534 8444 30540
rect 8312 30518 8432 30534
rect 8220 30382 8340 30410
rect 8312 30054 8340 30382
rect 8404 30138 8432 30518
rect 8496 30326 8524 32399
rect 8760 32370 8812 32376
rect 8772 31958 8800 32370
rect 8760 31952 8812 31958
rect 8760 31894 8812 31900
rect 8864 31804 8892 34478
rect 9496 33992 9548 33998
rect 9496 33934 9548 33940
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9312 33448 9364 33454
rect 9312 33390 9364 33396
rect 9324 32774 9352 33390
rect 9404 33312 9456 33318
rect 9404 33254 9456 33260
rect 9416 33046 9444 33254
rect 9404 33040 9456 33046
rect 9404 32982 9456 32988
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8944 32496 8996 32502
rect 8942 32464 8944 32473
rect 8996 32464 8998 32473
rect 8942 32399 8998 32408
rect 8680 31776 8892 31804
rect 8680 31770 8708 31776
rect 8563 31742 8708 31770
rect 8563 31668 8591 31742
rect 8668 31680 8720 31686
rect 8563 31640 8616 31668
rect 8484 30320 8536 30326
rect 8484 30262 8536 30268
rect 8404 30110 8524 30138
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 8208 29708 8260 29714
rect 8208 29650 8260 29656
rect 8116 29028 8168 29034
rect 8116 28970 8168 28976
rect 8128 28694 8156 28970
rect 8220 28778 8248 29650
rect 8312 29306 8340 29990
rect 8392 29776 8444 29782
rect 8392 29718 8444 29724
rect 8300 29300 8352 29306
rect 8300 29242 8352 29248
rect 8220 28750 8340 28778
rect 8116 28688 8168 28694
rect 8312 28665 8340 28750
rect 8116 28630 8168 28636
rect 8298 28656 8354 28665
rect 8128 28150 8156 28630
rect 8298 28591 8300 28600
rect 8352 28591 8354 28600
rect 8300 28562 8352 28568
rect 8312 28531 8340 28562
rect 8404 28558 8432 29718
rect 8392 28552 8444 28558
rect 8392 28494 8444 28500
rect 8116 28144 8168 28150
rect 8116 28086 8168 28092
rect 8128 27946 8156 28086
rect 8404 28082 8432 28494
rect 8392 28076 8444 28082
rect 8392 28018 8444 28024
rect 8116 27940 8168 27946
rect 8116 27882 8168 27888
rect 8390 27568 8446 27577
rect 8390 27503 8392 27512
rect 8444 27503 8446 27512
rect 8392 27474 8444 27480
rect 8298 27160 8354 27169
rect 8298 27095 8354 27104
rect 8312 26926 8340 27095
rect 8404 27062 8432 27474
rect 8392 27056 8444 27062
rect 8392 26998 8444 27004
rect 8300 26920 8352 26926
rect 8036 26846 8248 26874
rect 8300 26862 8352 26868
rect 7932 25968 7984 25974
rect 7932 25910 7984 25916
rect 7656 25832 7708 25838
rect 7656 25774 7708 25780
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 7576 25265 7604 25638
rect 7562 25256 7618 25265
rect 7562 25191 7618 25200
rect 7576 23497 7604 25191
rect 7668 24682 7696 25774
rect 7944 25430 7972 25910
rect 7932 25424 7984 25430
rect 7932 25366 7984 25372
rect 7656 24676 7708 24682
rect 7656 24618 7708 24624
rect 7668 24138 7696 24618
rect 7932 24200 7984 24206
rect 7932 24142 7984 24148
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7668 23730 7696 24074
rect 7656 23724 7708 23730
rect 7656 23666 7708 23672
rect 7562 23488 7618 23497
rect 7562 23423 7618 23432
rect 7944 23322 7972 24142
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 7562 23080 7618 23089
rect 7562 23015 7618 23024
rect 7576 21554 7604 23015
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7760 20262 7788 20946
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7760 19394 7788 20198
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7852 19514 7880 19926
rect 7944 19786 7972 23258
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 8128 22778 8156 23122
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8128 21593 8156 22714
rect 8114 21584 8170 21593
rect 8114 21519 8170 21528
rect 7932 19780 7984 19786
rect 7932 19722 7984 19728
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7760 19366 7880 19394
rect 7944 19378 7972 19722
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7576 16658 7604 17002
rect 7760 16658 7788 17070
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 7576 15706 7604 16594
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7562 14920 7618 14929
rect 7562 14855 7618 14864
rect 7576 14550 7604 14855
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7576 14074 7604 14486
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7576 13841 7604 14010
rect 7562 13832 7618 13841
rect 7562 13767 7564 13776
rect 7616 13767 7618 13776
rect 7564 13738 7616 13744
rect 7576 13530 7604 13738
rect 7760 13530 7788 14418
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7668 11762 7696 12378
rect 7760 12306 7788 12582
rect 7852 12481 7880 19366
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7944 18698 7972 19314
rect 8024 18896 8076 18902
rect 8024 18838 8076 18844
rect 7932 18692 7984 18698
rect 7932 18634 7984 18640
rect 8036 18426 8064 18838
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 8220 17513 8248 26846
rect 8496 26772 8524 30110
rect 8588 29238 8616 31640
rect 8668 31622 8720 31628
rect 8680 31278 8708 31622
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9324 31346 9352 32710
rect 9416 32298 9444 32982
rect 9404 32292 9456 32298
rect 9404 32234 9456 32240
rect 9312 31340 9364 31346
rect 9312 31282 9364 31288
rect 8668 31272 8720 31278
rect 8668 31214 8720 31220
rect 8668 31136 8720 31142
rect 8668 31078 8720 31084
rect 8680 29714 8708 31078
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8760 30184 8812 30190
rect 8758 30152 8760 30161
rect 8812 30152 8814 30161
rect 8758 30087 8814 30096
rect 9416 30054 9444 32234
rect 9508 30938 9536 33934
rect 9496 30932 9548 30938
rect 9496 30874 9548 30880
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 9404 30048 9456 30054
rect 9404 29990 9456 29996
rect 8668 29708 8720 29714
rect 8668 29650 8720 29656
rect 8680 29306 8708 29650
rect 8852 29640 8904 29646
rect 8852 29582 8904 29588
rect 8668 29300 8720 29306
rect 8668 29242 8720 29248
rect 8576 29232 8628 29238
rect 8576 29174 8628 29180
rect 8576 29096 8628 29102
rect 8576 29038 8628 29044
rect 8312 26744 8524 26772
rect 8312 26450 8340 26744
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8312 26042 8340 26386
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 8312 24721 8340 25978
rect 8404 25906 8432 26318
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8404 25498 8432 25842
rect 8392 25492 8444 25498
rect 8392 25434 8444 25440
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8496 24954 8524 25230
rect 8484 24948 8536 24954
rect 8484 24890 8536 24896
rect 8298 24712 8354 24721
rect 8298 24647 8354 24656
rect 8392 24268 8444 24274
rect 8392 24210 8444 24216
rect 8404 23526 8432 24210
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8300 21480 8352 21486
rect 8404 21457 8432 23462
rect 8484 22976 8536 22982
rect 8484 22918 8536 22924
rect 8496 22574 8524 22918
rect 8484 22568 8536 22574
rect 8484 22510 8536 22516
rect 8300 21422 8352 21428
rect 8390 21448 8446 21457
rect 8312 21350 8340 21422
rect 8390 21383 8446 21392
rect 8300 21344 8352 21350
rect 8298 21312 8300 21321
rect 8352 21312 8354 21321
rect 8298 21247 8354 21256
rect 8312 20398 8340 21247
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8496 20346 8524 22510
rect 8588 21010 8616 29038
rect 8680 28694 8708 29242
rect 8864 29170 8892 29582
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 9324 28762 9352 29990
rect 9312 28756 9364 28762
rect 9312 28698 9364 28704
rect 8668 28688 8720 28694
rect 8668 28630 8720 28636
rect 8680 28218 8708 28630
rect 9404 28416 9456 28422
rect 9404 28358 9456 28364
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 9416 28014 9444 28358
rect 9404 28008 9456 28014
rect 9404 27950 9456 27956
rect 9416 27334 9444 27950
rect 9600 27441 9628 35770
rect 9784 35601 9812 36178
rect 9770 35592 9826 35601
rect 9770 35527 9826 35536
rect 9784 35494 9812 35527
rect 9772 35488 9824 35494
rect 9772 35430 9824 35436
rect 9680 33992 9732 33998
rect 9680 33934 9732 33940
rect 9692 33522 9720 33934
rect 9680 33516 9732 33522
rect 9680 33458 9732 33464
rect 9692 32026 9720 33458
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 9784 31906 9812 35430
rect 9968 35290 9996 36518
rect 9956 35284 10008 35290
rect 9956 35226 10008 35232
rect 9968 34610 9996 35226
rect 10152 34746 10180 39520
rect 10692 36576 10744 36582
rect 10692 36518 10744 36524
rect 10324 36032 10376 36038
rect 10324 35974 10376 35980
rect 10336 35698 10364 35974
rect 10324 35692 10376 35698
rect 10324 35634 10376 35640
rect 10416 35556 10468 35562
rect 10416 35498 10468 35504
rect 10140 34740 10192 34746
rect 10140 34682 10192 34688
rect 9956 34604 10008 34610
rect 9956 34546 10008 34552
rect 10232 34400 10284 34406
rect 10232 34342 10284 34348
rect 10048 34128 10100 34134
rect 10048 34070 10100 34076
rect 10060 33318 10088 34070
rect 10244 33658 10272 34342
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 10048 33312 10100 33318
rect 10048 33254 10100 33260
rect 10428 33114 10456 35498
rect 10600 35216 10652 35222
rect 10600 35158 10652 35164
rect 10612 34406 10640 35158
rect 10704 34785 10732 36518
rect 10784 35692 10836 35698
rect 10784 35634 10836 35640
rect 10690 34776 10746 34785
rect 10690 34711 10746 34720
rect 10600 34400 10652 34406
rect 10600 34342 10652 34348
rect 10416 33108 10468 33114
rect 10416 33050 10468 33056
rect 10416 32904 10468 32910
rect 10416 32846 10468 32852
rect 10232 32292 10284 32298
rect 10232 32234 10284 32240
rect 9692 31878 9812 31906
rect 10244 31890 10272 32234
rect 10428 32230 10456 32846
rect 10704 32586 10732 34711
rect 10796 34610 10824 35634
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 10784 34604 10836 34610
rect 10784 34546 10836 34552
rect 10796 33930 10824 34546
rect 10784 33924 10836 33930
rect 10784 33866 10836 33872
rect 10612 32558 10732 32586
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 10232 31884 10284 31890
rect 9692 29034 9720 31878
rect 10232 31826 10284 31832
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 10152 31278 10180 31758
rect 10244 31482 10272 31826
rect 10232 31476 10284 31482
rect 10232 31418 10284 31424
rect 10140 31272 10192 31278
rect 10140 31214 10192 31220
rect 9864 30864 9916 30870
rect 10152 30841 10180 31214
rect 9864 30806 9916 30812
rect 10138 30832 10194 30841
rect 9876 30138 9904 30806
rect 10138 30767 10194 30776
rect 9784 30122 9904 30138
rect 9956 30184 10008 30190
rect 9956 30126 10008 30132
rect 9772 30116 9904 30122
rect 9824 30110 9904 30116
rect 9772 30058 9824 30064
rect 9968 29510 9996 30126
rect 10416 30116 10468 30122
rect 10416 30058 10468 30064
rect 10428 29782 10456 30058
rect 10416 29776 10468 29782
rect 10416 29718 10468 29724
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9680 29028 9732 29034
rect 9680 28970 9732 28976
rect 9968 28762 9996 29446
rect 10428 29306 10456 29718
rect 10416 29300 10468 29306
rect 10416 29242 10468 29248
rect 10324 29028 10376 29034
rect 10324 28970 10376 28976
rect 10336 28914 10364 28970
rect 10414 28928 10470 28937
rect 10336 28886 10414 28914
rect 10414 28863 10470 28872
rect 9956 28756 10008 28762
rect 9956 28698 10008 28704
rect 10416 28552 10468 28558
rect 10416 28494 10468 28500
rect 10140 28008 10192 28014
rect 10140 27950 10192 27956
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 9772 27464 9824 27470
rect 9586 27432 9642 27441
rect 9772 27406 9824 27412
rect 9586 27367 9642 27376
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 8864 25498 8892 27270
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 9312 26036 9364 26042
rect 9312 25978 9364 25984
rect 8852 25492 8904 25498
rect 8852 25434 8904 25440
rect 8758 25392 8814 25401
rect 8758 25327 8814 25336
rect 8772 24410 8800 25327
rect 8864 24818 8892 25434
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 9218 24848 9274 24857
rect 8852 24812 8904 24818
rect 9218 24783 9274 24792
rect 8852 24754 8904 24760
rect 9232 24562 9260 24783
rect 9324 24682 9352 25978
rect 9312 24676 9364 24682
rect 9312 24618 9364 24624
rect 9232 24534 9352 24562
rect 8760 24404 8812 24410
rect 8760 24346 8812 24352
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8680 23594 8708 24074
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 8668 23588 8720 23594
rect 8668 23530 8720 23536
rect 8680 22545 8708 23530
rect 8942 23488 8998 23497
rect 8942 23423 8998 23432
rect 8956 23322 8984 23423
rect 8944 23316 8996 23322
rect 8944 23258 8996 23264
rect 8956 23202 8984 23258
rect 8864 23174 8984 23202
rect 8864 22574 8892 23174
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8852 22568 8904 22574
rect 8666 22536 8722 22545
rect 8852 22510 8904 22516
rect 8666 22471 8722 22480
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9140 22234 9168 22442
rect 9128 22228 9180 22234
rect 9128 22170 9180 22176
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8772 21622 8800 21966
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8760 21616 8812 21622
rect 8760 21558 8812 21564
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8760 20392 8812 20398
rect 8496 20318 8616 20346
rect 8760 20334 8812 20340
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8312 18970 8340 19790
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19378 8432 19654
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8392 19236 8444 19242
rect 8392 19178 8444 19184
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8206 17504 8262 17513
rect 8206 17439 8262 17448
rect 8312 17338 8340 17614
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8022 17096 8078 17105
rect 8312 17066 8340 17274
rect 8022 17031 8078 17040
rect 8300 17060 8352 17066
rect 8036 16794 8064 17031
rect 8300 17002 8352 17008
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8404 16674 8432 19178
rect 8496 18426 8524 20198
rect 8588 18766 8616 20318
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8496 17898 8524 18362
rect 8496 17870 8616 17898
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8496 16697 8524 17478
rect 8588 17202 8616 17870
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8220 16646 8432 16674
rect 8482 16688 8538 16697
rect 8036 15570 8064 16594
rect 8220 16590 8248 16646
rect 8482 16623 8538 16632
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8220 16250 8248 16526
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8116 15496 8168 15502
rect 8036 15444 8116 15450
rect 8036 15438 8168 15444
rect 8036 15422 8156 15438
rect 8220 15434 8248 16186
rect 8772 15978 8800 20334
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8956 18737 8984 19314
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9232 18873 9260 19246
rect 9218 18864 9274 18873
rect 9218 18799 9274 18808
rect 8942 18728 8998 18737
rect 8942 18663 8998 18672
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8864 17066 8892 17546
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8852 17060 8904 17066
rect 8852 17002 8904 17008
rect 8864 16046 8892 17002
rect 9140 16794 9168 17138
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8864 15638 8892 15982
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8208 15428 8260 15434
rect 7838 12472 7894 12481
rect 7838 12407 7894 12416
rect 7930 12336 7986 12345
rect 7748 12300 7800 12306
rect 7930 12271 7986 12280
rect 7748 12242 7800 12248
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7576 9926 7604 10542
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9586 7604 9862
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7668 8498 7696 8774
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7392 7546 7420 8298
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7392 7274 7420 7482
rect 7668 7410 7696 8026
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7392 6458 7420 7210
rect 7852 6934 7880 7210
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7392 6186 7420 6394
rect 7470 6352 7526 6361
rect 7470 6287 7472 6296
rect 7524 6287 7526 6296
rect 7472 6258 7524 6264
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7102 5743 7158 5752
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7102 5672 7158 5681
rect 6932 5522 6960 5646
rect 7102 5607 7158 5616
rect 6840 5494 6960 5522
rect 6840 5302 6868 5494
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6828 5160 6880 5166
rect 6826 5128 6828 5137
rect 6880 5128 6882 5137
rect 6826 5063 6882 5072
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7024 4185 7052 4966
rect 7116 4826 7144 5607
rect 7208 5370 7236 5714
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7010 4176 7066 4185
rect 7116 4146 7144 4762
rect 7300 4690 7328 5850
rect 7392 4758 7420 6122
rect 7380 4752 7432 4758
rect 7944 4729 7972 12271
rect 8036 11336 8064 15422
rect 8208 15370 8260 15376
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8128 15026 8156 15302
rect 8220 15162 8248 15370
rect 8298 15192 8354 15201
rect 8208 15156 8260 15162
rect 8298 15127 8300 15136
rect 8208 15098 8260 15104
rect 8352 15127 8354 15136
rect 8300 15098 8352 15104
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8312 14958 8340 15098
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8496 14482 8524 14758
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8680 14278 8708 14894
rect 8864 14618 8892 15574
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8220 13462 8248 14214
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8208 13456 8260 13462
rect 8128 13404 8208 13410
rect 8128 13398 8260 13404
rect 8128 13382 8248 13398
rect 8128 12986 8156 13382
rect 8312 12986 8340 13806
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8312 12714 8340 12922
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8220 11898 8248 12310
rect 8496 12170 8524 12854
rect 8588 12442 8616 13262
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8588 11354 8616 12174
rect 8680 11830 8708 14214
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8772 12850 8800 13126
rect 8864 12850 8892 13262
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8772 12170 8800 12786
rect 9324 12730 9352 24534
rect 9416 24177 9444 27270
rect 9784 27169 9812 27406
rect 9770 27160 9826 27169
rect 9600 27118 9770 27146
rect 9600 26518 9628 27118
rect 9770 27095 9826 27104
rect 9876 26994 9904 27542
rect 9864 26988 9916 26994
rect 9864 26930 9916 26936
rect 9678 26888 9734 26897
rect 9678 26823 9680 26832
rect 9732 26823 9734 26832
rect 9772 26852 9824 26858
rect 9680 26794 9732 26800
rect 9772 26794 9824 26800
rect 9692 26586 9720 26794
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9588 26512 9640 26518
rect 9588 26454 9640 26460
rect 9784 26058 9812 26794
rect 9876 26518 9904 26930
rect 10152 26874 10180 27950
rect 10324 27872 10376 27878
rect 10324 27814 10376 27820
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10244 27062 10272 27406
rect 10232 27056 10284 27062
rect 10232 26998 10284 27004
rect 10152 26846 10272 26874
rect 9864 26512 9916 26518
rect 9864 26454 9916 26460
rect 10138 26480 10194 26489
rect 9508 26042 9812 26058
rect 9876 26042 9904 26454
rect 10138 26415 10194 26424
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9496 26036 9812 26042
rect 9548 26030 9812 26036
rect 9864 26036 9916 26042
rect 9496 25978 9548 25984
rect 9864 25978 9916 25984
rect 9968 25498 9996 26318
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 10060 25838 10088 26182
rect 10048 25832 10100 25838
rect 10046 25800 10048 25809
rect 10100 25800 10102 25809
rect 10046 25735 10102 25744
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 10152 25362 10180 26415
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 10048 24948 10100 24954
rect 10048 24890 10100 24896
rect 9494 24848 9550 24857
rect 9494 24783 9496 24792
rect 9548 24783 9550 24792
rect 9496 24754 9548 24760
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9402 24168 9458 24177
rect 9402 24103 9458 24112
rect 9692 23594 9720 24210
rect 9862 24168 9918 24177
rect 9862 24103 9864 24112
rect 9916 24103 9918 24112
rect 9864 24074 9916 24080
rect 9680 23588 9732 23594
rect 9680 23530 9732 23536
rect 9864 23520 9916 23526
rect 9862 23488 9864 23497
rect 9916 23488 9918 23497
rect 9862 23423 9918 23432
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9692 23089 9720 23122
rect 9678 23080 9734 23089
rect 9678 23015 9734 23024
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 9680 22568 9732 22574
rect 9586 22536 9642 22545
rect 9680 22510 9732 22516
rect 9586 22471 9642 22480
rect 9508 22030 9536 22061
rect 9496 22024 9548 22030
rect 9494 21992 9496 22001
rect 9548 21992 9550 22001
rect 9494 21927 9550 21936
rect 9508 21690 9536 21927
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 9508 21146 9536 21626
rect 9600 21554 9628 22471
rect 9692 21894 9720 22510
rect 9876 22001 9904 22578
rect 10060 22234 10088 24890
rect 10152 24410 10180 25298
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 10244 24290 10272 26846
rect 10152 24262 10272 24290
rect 10048 22228 10100 22234
rect 10048 22170 10100 22176
rect 9862 21992 9918 22001
rect 9862 21927 9918 21936
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9692 21486 9720 21830
rect 9680 21480 9732 21486
rect 9600 21428 9680 21434
rect 9600 21422 9732 21428
rect 9600 21406 9720 21422
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9600 20777 9628 21406
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9784 20806 9812 21286
rect 9680 20800 9732 20806
rect 9586 20768 9642 20777
rect 9680 20742 9732 20748
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9586 20703 9642 20712
rect 9600 20262 9628 20703
rect 9692 20398 9720 20742
rect 9784 20602 9812 20742
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9692 19922 9720 20334
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9956 19780 10008 19786
rect 9956 19722 10008 19728
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9600 18426 9628 18906
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9784 18222 9812 18770
rect 9876 18698 9904 19246
rect 9968 19242 9996 19722
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9968 18970 9996 19178
rect 10060 18970 10088 19858
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9876 18358 9904 18634
rect 10152 18426 10180 24262
rect 10232 23656 10284 23662
rect 10230 23624 10232 23633
rect 10284 23624 10286 23633
rect 10230 23559 10286 23568
rect 10244 23322 10272 23559
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10244 22234 10272 22510
rect 10232 22228 10284 22234
rect 10232 22170 10284 22176
rect 10244 21146 10272 22170
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 10336 19854 10364 27814
rect 10428 24342 10456 28494
rect 10612 25786 10640 32558
rect 10692 32360 10744 32366
rect 10692 32302 10744 32308
rect 10704 31958 10732 32302
rect 10692 31952 10744 31958
rect 10690 31920 10692 31929
rect 10744 31920 10746 31929
rect 10690 31855 10746 31864
rect 10796 31346 10824 33866
rect 10980 33862 11008 35022
rect 11072 34746 11100 39520
rect 11900 37754 11928 39520
rect 12346 38176 12402 38185
rect 12346 38111 12402 38120
rect 11900 37726 12020 37754
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11242 35184 11298 35193
rect 11242 35119 11298 35128
rect 11060 34740 11112 34746
rect 11060 34682 11112 34688
rect 11060 34128 11112 34134
rect 11060 34070 11112 34076
rect 10968 33856 11020 33862
rect 10968 33798 11020 33804
rect 10876 33380 10928 33386
rect 10876 33322 10928 33328
rect 10888 33114 10916 33322
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 10980 33017 11008 33798
rect 11072 33318 11100 34070
rect 11152 33448 11204 33454
rect 11150 33416 11152 33425
rect 11204 33416 11206 33425
rect 11150 33351 11206 33360
rect 11060 33312 11112 33318
rect 11060 33254 11112 33260
rect 11072 33046 11100 33254
rect 11060 33040 11112 33046
rect 10966 33008 11022 33017
rect 11060 32982 11112 32988
rect 10966 32943 11022 32952
rect 11256 31890 11284 35119
rect 11520 35080 11572 35086
rect 11520 35022 11572 35028
rect 11336 33992 11388 33998
rect 11336 33934 11388 33940
rect 11348 32774 11376 33934
rect 11532 33561 11560 35022
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11992 33658 12020 37726
rect 12072 35148 12124 35154
rect 12072 35090 12124 35096
rect 12084 34542 12112 35090
rect 12072 34536 12124 34542
rect 12072 34478 12124 34484
rect 12084 34082 12112 34478
rect 12084 34066 12204 34082
rect 12084 34060 12216 34066
rect 12084 34054 12164 34060
rect 11980 33652 12032 33658
rect 11980 33594 12032 33600
rect 11518 33552 11574 33561
rect 11518 33487 11574 33496
rect 11532 32994 11560 33487
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11704 33040 11756 33046
rect 11440 32966 11652 32994
rect 11704 32982 11756 32988
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11440 32348 11468 32966
rect 11624 32910 11652 32966
rect 11520 32904 11572 32910
rect 11520 32846 11572 32852
rect 11612 32904 11664 32910
rect 11612 32846 11664 32852
rect 11348 32320 11468 32348
rect 11244 31884 11296 31890
rect 11244 31826 11296 31832
rect 10784 31340 10836 31346
rect 10784 31282 10836 31288
rect 10796 30938 10824 31282
rect 10968 31204 11020 31210
rect 10968 31146 11020 31152
rect 10784 30932 10836 30938
rect 10784 30874 10836 30880
rect 10980 29850 11008 31146
rect 11256 31142 11284 31826
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 11348 30734 11376 32320
rect 11532 32026 11560 32846
rect 11716 32570 11744 32982
rect 11704 32564 11756 32570
rect 11704 32506 11756 32512
rect 12084 32473 12112 34054
rect 12164 34002 12216 34008
rect 12256 33448 12308 33454
rect 12256 33390 12308 33396
rect 12070 32464 12126 32473
rect 12070 32399 12126 32408
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 11520 31136 11572 31142
rect 11520 31078 11572 31084
rect 11428 30864 11480 30870
rect 11428 30806 11480 30812
rect 11336 30728 11388 30734
rect 11058 30696 11114 30705
rect 11336 30670 11388 30676
rect 11058 30631 11114 30640
rect 11072 30122 11100 30631
rect 11348 30258 11376 30670
rect 11440 30394 11468 30806
rect 11428 30388 11480 30394
rect 11428 30330 11480 30336
rect 11336 30252 11388 30258
rect 11336 30194 11388 30200
rect 11060 30116 11112 30122
rect 11060 30058 11112 30064
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 10692 29640 10744 29646
rect 10692 29582 10744 29588
rect 10704 28966 10732 29582
rect 11058 29064 11114 29073
rect 11058 28999 11114 29008
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10704 28082 10732 28902
rect 11072 28218 11100 28999
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10692 28076 10744 28082
rect 10692 28018 10744 28024
rect 11256 27878 11284 28562
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 11426 27568 11482 27577
rect 11532 27554 11560 31078
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11980 29776 12032 29782
rect 11980 29718 12032 29724
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 11900 29306 11928 29582
rect 11888 29300 11940 29306
rect 11888 29242 11940 29248
rect 11992 29102 12020 29718
rect 11980 29096 12032 29102
rect 11980 29038 12032 29044
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11482 27526 11560 27554
rect 11980 27600 12032 27606
rect 11980 27542 12032 27548
rect 12084 27554 12112 32399
rect 12164 32224 12216 32230
rect 12164 32166 12216 32172
rect 12176 31793 12204 32166
rect 12162 31784 12218 31793
rect 12162 31719 12218 31728
rect 12164 31204 12216 31210
rect 12164 31146 12216 31152
rect 12176 30734 12204 31146
rect 12164 30728 12216 30734
rect 12164 30670 12216 30676
rect 12176 30161 12204 30670
rect 12162 30152 12218 30161
rect 12162 30087 12218 30096
rect 12176 29646 12204 30087
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 11426 27503 11482 27512
rect 11058 27024 11114 27033
rect 11058 26959 11114 26968
rect 11336 26988 11388 26994
rect 11072 26926 11100 26959
rect 11336 26930 11388 26936
rect 11060 26920 11112 26926
rect 11060 26862 11112 26868
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 11072 26382 11100 26726
rect 11348 26518 11376 26930
rect 11336 26512 11388 26518
rect 11336 26454 11388 26460
rect 11440 26466 11468 27503
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 11532 26586 11560 27406
rect 11992 27130 12020 27542
rect 12084 27526 12204 27554
rect 12072 27464 12124 27470
rect 12072 27406 12124 27412
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 11992 26790 12020 27066
rect 12084 26858 12112 27406
rect 12072 26852 12124 26858
rect 12072 26794 12124 26800
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11520 26580 11572 26586
rect 11520 26522 11572 26528
rect 11060 26376 11112 26382
rect 11060 26318 11112 26324
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 11058 26208 11114 26217
rect 11058 26143 11114 26152
rect 10968 25832 11020 25838
rect 10508 25764 10560 25770
rect 10612 25758 10732 25786
rect 10968 25774 11020 25780
rect 10508 25706 10560 25712
rect 10520 25430 10548 25706
rect 10508 25424 10560 25430
rect 10508 25366 10560 25372
rect 10520 24954 10548 25366
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10598 24712 10654 24721
rect 10598 24647 10654 24656
rect 10416 24336 10468 24342
rect 10416 24278 10468 24284
rect 10428 23730 10456 24278
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 10416 23588 10468 23594
rect 10416 23530 10468 23536
rect 10428 22642 10456 23530
rect 10508 23520 10560 23526
rect 10508 23462 10560 23468
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10428 20398 10456 21014
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10428 19922 10456 20334
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10322 19680 10378 19689
rect 10322 19615 10378 19624
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 9772 18216 9824 18222
rect 9586 18184 9642 18193
rect 9772 18158 9824 18164
rect 9586 18119 9588 18128
rect 9640 18119 9642 18128
rect 9588 18090 9640 18096
rect 9600 17882 9628 18090
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9600 17202 9628 17818
rect 9784 17814 9812 18158
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9876 17610 9904 18294
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9692 17066 9720 17478
rect 9876 17338 9904 17546
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9416 16114 9444 16730
rect 9494 16688 9550 16697
rect 9494 16623 9550 16632
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9402 16008 9458 16017
rect 9402 15943 9404 15952
rect 9456 15943 9458 15952
rect 9404 15914 9456 15920
rect 9508 15722 9536 16623
rect 9600 15994 9628 16934
rect 9692 16658 9720 17002
rect 9770 16824 9826 16833
rect 9770 16759 9826 16768
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9692 16130 9720 16594
rect 9784 16522 9812 16759
rect 9954 16688 10010 16697
rect 9954 16623 9956 16632
rect 10008 16623 10010 16632
rect 9956 16594 10008 16600
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9784 16250 9812 16458
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9692 16102 9812 16130
rect 9600 15966 9720 15994
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9416 15706 9536 15722
rect 9416 15700 9548 15706
rect 9416 15694 9496 15700
rect 9416 15162 9444 15694
rect 9496 15642 9548 15648
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9508 14618 9536 15506
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9600 14482 9628 15846
rect 9692 15570 9720 15966
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9784 15162 9812 16102
rect 10048 15632 10100 15638
rect 10048 15574 10100 15580
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 10060 14822 10088 15574
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9692 14618 9720 14758
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 14074 9628 14418
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9692 13938 9720 14554
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9692 13841 9720 13874
rect 9678 13832 9734 13841
rect 9678 13767 9734 13776
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 8864 12702 9352 12730
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8576 11348 8628 11354
rect 8036 11308 8248 11336
rect 8114 11248 8170 11257
rect 8114 11183 8170 11192
rect 8128 11014 8156 11183
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10198 8156 10950
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8128 9722 8156 10134
rect 8220 9722 8248 11308
rect 8576 11290 8628 11296
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10810 8432 10950
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8312 9042 8340 9658
rect 8404 9654 8432 9998
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8392 9512 8444 9518
rect 8390 9480 8392 9489
rect 8444 9480 8446 9489
rect 8680 9450 8708 11766
rect 8772 11121 8800 12106
rect 8758 11112 8814 11121
rect 8758 11047 8814 11056
rect 8772 10198 8800 11047
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8864 9518 8892 12702
rect 9600 12442 9628 13262
rect 10060 12850 10088 13398
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9508 11354 9536 11562
rect 9968 11558 9996 12242
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 11830 10088 12038
rect 10152 11898 10180 12242
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9864 11280 9916 11286
rect 9862 11248 9864 11257
rect 9916 11248 9918 11257
rect 9862 11183 9918 11192
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 9876 10810 9904 11183
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9324 10266 9352 10474
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8390 9415 8446 9424
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8312 8634 8340 8978
rect 8588 8820 8616 9318
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8668 8832 8720 8838
rect 8588 8792 8668 8820
rect 8668 8774 8720 8780
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8680 8430 8708 8774
rect 8772 8430 8800 8842
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8772 8022 8800 8366
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 6730 8156 7822
rect 8220 7546 8248 7958
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8772 7206 8800 7958
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8220 5914 8248 6802
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8588 6458 8616 6598
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8772 5914 8800 6598
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9324 6186 9352 7822
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 9324 5574 9352 6122
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 8772 5234 8800 5510
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8220 4826 8248 4966
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 7380 4694 7432 4700
rect 7930 4720 7986 4729
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7300 4214 7328 4626
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7010 4111 7066 4120
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7286 4040 7342 4049
rect 7392 4010 7420 4694
rect 7930 4655 7986 4664
rect 8220 4282 8248 4762
rect 8404 4622 8432 5034
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 7286 3975 7342 3984
rect 7380 4004 7432 4010
rect 6184 3470 6236 3476
rect 6642 3496 6698 3505
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6012 2650 6040 3130
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6196 2582 6224 3470
rect 6642 3431 6698 3440
rect 6656 2961 6684 3431
rect 6826 3088 6882 3097
rect 6826 3023 6882 3032
rect 6840 2990 6868 3023
rect 6828 2984 6880 2990
rect 6642 2952 6698 2961
rect 6828 2926 6880 2932
rect 7010 2952 7066 2961
rect 6642 2887 6698 2896
rect 7010 2887 7066 2896
rect 7024 2854 7052 2887
rect 7012 2848 7064 2854
rect 6734 2816 6790 2825
rect 6656 2774 6734 2802
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 6656 1714 6684 2774
rect 7012 2790 7064 2796
rect 6734 2751 6790 2760
rect 7010 2680 7066 2689
rect 7010 2615 7066 2624
rect 7024 2582 7052 2615
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 7300 2446 7328 3975
rect 7380 3946 7432 3952
rect 7392 3738 7420 3946
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7470 3360 7526 3369
rect 7470 3295 7526 3304
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 6564 1686 6684 1714
rect 5172 604 5224 610
rect 5172 546 5224 552
rect 5724 604 5776 610
rect 5724 546 5776 552
rect 5736 480 5764 546
rect 6564 480 6592 1686
rect 7484 480 7512 3295
rect 8036 3058 8064 3674
rect 8220 3670 8248 3878
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8220 3194 8248 3606
rect 8208 3188 8260 3194
rect 8260 3148 8340 3176
rect 8208 3130 8260 3136
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8220 2650 8248 3130
rect 8312 2922 8340 3148
rect 8772 3126 8800 5170
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8864 4214 8892 4490
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9232 3670 9260 4082
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8404 480 8432 2246
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 9324 1714 9352 3334
rect 9416 3108 9444 10678
rect 9494 10568 9550 10577
rect 9494 10503 9496 10512
rect 9548 10503 9550 10512
rect 9496 10474 9548 10480
rect 9586 10160 9642 10169
rect 9586 10095 9642 10104
rect 9772 10124 9824 10130
rect 9600 9586 9628 10095
rect 9772 10066 9824 10072
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9784 9382 9812 10066
rect 9968 10033 9996 11494
rect 10060 11286 10088 11766
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10060 10674 10088 11222
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10336 10606 10364 19615
rect 10428 19514 10456 19858
rect 10520 19786 10548 23462
rect 10612 22710 10640 24647
rect 10600 22704 10652 22710
rect 10600 22646 10652 22652
rect 10704 22080 10732 25758
rect 10980 25498 11008 25774
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10796 23526 10824 24754
rect 10968 24744 11020 24750
rect 10968 24686 11020 24692
rect 10980 24342 11008 24686
rect 10968 24336 11020 24342
rect 10966 24304 10968 24313
rect 11020 24304 11022 24313
rect 10966 24239 11022 24248
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10888 23730 10916 24006
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 11072 22522 11100 26143
rect 11164 24857 11192 26318
rect 11348 26042 11376 26454
rect 11440 26438 11560 26466
rect 11336 26036 11388 26042
rect 11336 25978 11388 25984
rect 11150 24848 11206 24857
rect 11150 24783 11206 24792
rect 11164 24206 11192 24783
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11256 24342 11284 24550
rect 11244 24336 11296 24342
rect 11244 24278 11296 24284
rect 11532 24290 11560 26438
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 11992 25702 12020 26318
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11992 25498 12020 25638
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 11796 25424 11848 25430
rect 11796 25366 11848 25372
rect 11808 24954 11836 25366
rect 11980 25288 12032 25294
rect 11980 25230 12032 25236
rect 11796 24948 11848 24954
rect 11796 24890 11848 24896
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11164 23798 11192 24142
rect 11256 23866 11284 24278
rect 11532 24262 11652 24290
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11152 23792 11204 23798
rect 11152 23734 11204 23740
rect 11334 23624 11390 23633
rect 11334 23559 11390 23568
rect 11244 23248 11296 23254
rect 11244 23190 11296 23196
rect 10888 22494 11100 22522
rect 10704 22052 10824 22080
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10704 19922 10732 20266
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10508 19780 10560 19786
rect 10508 19722 10560 19728
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10428 18902 10456 19450
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10416 18896 10468 18902
rect 10468 18844 10548 18850
rect 10416 18838 10548 18844
rect 10428 18822 10548 18838
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10428 18222 10456 18702
rect 10520 18426 10548 18822
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10612 17882 10640 18906
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10506 17640 10562 17649
rect 10506 17575 10562 17584
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 9954 10024 10010 10033
rect 9954 9959 10010 9968
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7410 9536 7686
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9784 7313 9812 9318
rect 9968 7954 9996 9959
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9968 7546 9996 7890
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9770 7304 9826 7313
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9680 7268 9732 7274
rect 9770 7239 9826 7248
rect 9680 7210 9732 7216
rect 9508 7002 9536 7210
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9692 6730 9720 7210
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 6610 9720 6666
rect 9600 6582 9720 6610
rect 9600 4146 9628 6582
rect 9692 6458 9720 6582
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9876 6390 9904 6870
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10152 6746 10180 9386
rect 10244 6905 10272 9658
rect 10230 6896 10286 6905
rect 10230 6831 10286 6840
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 10060 6322 10088 6734
rect 10152 6718 10272 6746
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9692 6225 9720 6258
rect 9678 6216 9734 6225
rect 9678 6151 9734 6160
rect 9678 5808 9734 5817
rect 9678 5743 9680 5752
rect 9732 5743 9734 5752
rect 9680 5714 9732 5720
rect 9692 5370 9720 5714
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9692 4321 9720 5306
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9678 4312 9734 4321
rect 9678 4247 9734 4256
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3528 9640 3534
rect 9692 3505 9720 3538
rect 9588 3470 9640 3476
rect 9678 3496 9734 3505
rect 9600 3194 9628 3470
rect 9678 3431 9734 3440
rect 9588 3188 9640 3194
rect 9784 3176 9812 4966
rect 9876 3641 9904 5102
rect 9862 3632 9918 3641
rect 9862 3567 9918 3576
rect 10140 3596 10192 3602
rect 9640 3148 9812 3176
rect 9588 3130 9640 3136
rect 9416 3080 9536 3108
rect 9508 2650 9536 3080
rect 9876 3058 9904 3567
rect 10140 3538 10192 3544
rect 10152 3194 10180 3538
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9232 1686 9352 1714
rect 9232 480 9260 1686
rect 10152 480 10180 2790
rect 10244 2514 10272 6718
rect 10336 4690 10364 10542
rect 10428 9722 10456 16526
rect 10520 12714 10548 17575
rect 10612 17134 10640 17818
rect 10704 17814 10732 18022
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10612 16658 10640 17070
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 13802 10640 14758
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10612 13462 10640 13738
rect 10704 13734 10732 14214
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10704 12782 10732 13670
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10704 12442 10732 12718
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10612 10810 10640 11086
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10796 10130 10824 22052
rect 10888 20534 10916 22494
rect 11256 22438 11284 23190
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 10980 22234 11008 22374
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 11072 21978 11100 22374
rect 10980 21962 11100 21978
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 10968 21956 11100 21962
rect 11020 21950 11100 21956
rect 10968 21898 11020 21904
rect 11164 21690 11192 21966
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11150 21448 11206 21457
rect 11150 21383 11206 21392
rect 11164 21146 11192 21383
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11164 20777 11192 20946
rect 11150 20768 11206 20777
rect 11150 20703 11206 20712
rect 10876 20528 10928 20534
rect 10876 20470 10928 20476
rect 10888 20058 10916 20470
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10888 19514 10916 19994
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10888 19310 10916 19450
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 11242 18864 11298 18873
rect 11242 18799 11244 18808
rect 11296 18799 11298 18808
rect 11244 18770 11296 18776
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10968 17536 11020 17542
rect 11072 17524 11100 18022
rect 11020 17496 11100 17524
rect 10968 17478 11020 17484
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16794 10916 17070
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10966 16552 11022 16561
rect 10966 16487 11022 16496
rect 10980 16250 11008 16487
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11072 16130 11100 16934
rect 11164 16697 11192 18566
rect 11256 18426 11284 18770
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11256 17134 11284 17614
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11150 16688 11206 16697
rect 11150 16623 11206 16632
rect 10888 16102 11100 16130
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11152 16108 11204 16114
rect 10888 15065 10916 16102
rect 11152 16050 11204 16056
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10980 15586 11008 15914
rect 11164 15706 11192 16050
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 10980 15558 11100 15586
rect 11072 15162 11100 15558
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10874 15056 10930 15065
rect 10874 14991 10930 15000
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10888 11665 10916 14826
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10980 14074 11008 14214
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10980 11694 11008 11834
rect 10968 11688 11020 11694
rect 10874 11656 10930 11665
rect 10968 11630 11020 11636
rect 10874 11591 10930 11600
rect 10980 10713 11008 11630
rect 10966 10704 11022 10713
rect 10966 10639 11022 10648
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 11256 9081 11284 16118
rect 11348 14890 11376 23559
rect 11428 23316 11480 23322
rect 11428 23258 11480 23264
rect 11440 22778 11468 23258
rect 11532 23118 11560 24142
rect 11624 23594 11652 24262
rect 11992 24070 12020 25230
rect 12084 24206 12112 26794
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 12176 23633 12204 27526
rect 12268 26926 12296 33390
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 12162 23624 12218 23633
rect 11612 23588 11664 23594
rect 12162 23559 12218 23568
rect 11612 23530 11664 23536
rect 12164 23520 12216 23526
rect 12070 23488 12126 23497
rect 11992 23446 12070 23474
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11520 23112 11572 23118
rect 11520 23054 11572 23060
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 11440 21350 11468 22034
rect 11886 21992 11942 22001
rect 11886 21927 11888 21936
rect 11940 21927 11942 21936
rect 11888 21898 11940 21904
rect 11900 21418 11928 21898
rect 11520 21412 11572 21418
rect 11520 21354 11572 21360
rect 11888 21412 11940 21418
rect 11888 21354 11940 21360
rect 11428 21344 11480 21350
rect 11426 21312 11428 21321
rect 11480 21312 11482 21321
rect 11426 21247 11482 21256
rect 11532 20874 11560 21354
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11992 21078 12020 23446
rect 12164 23462 12216 23468
rect 12070 23423 12126 23432
rect 12072 22228 12124 22234
rect 12072 22170 12124 22176
rect 12084 22098 12112 22170
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12084 21146 12112 22034
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 11980 21072 12032 21078
rect 11980 21014 12032 21020
rect 11612 21004 11664 21010
rect 11612 20946 11664 20952
rect 11520 20868 11572 20874
rect 11520 20810 11572 20816
rect 11624 20806 11652 20946
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11978 20768 12034 20777
rect 11624 20330 11652 20742
rect 11978 20703 12034 20712
rect 11992 20602 12020 20703
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11612 20324 11664 20330
rect 11612 20266 11664 20272
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11532 19514 11560 19858
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11428 18692 11480 18698
rect 11428 18634 11480 18640
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11348 14006 11376 14418
rect 11336 14000 11388 14006
rect 11334 13968 11336 13977
rect 11388 13968 11390 13977
rect 11334 13903 11390 13912
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11348 12918 11376 13330
rect 11336 12912 11388 12918
rect 11334 12880 11336 12889
rect 11388 12880 11390 12889
rect 11334 12815 11390 12824
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11242 9072 11298 9081
rect 11242 9007 11298 9016
rect 10690 4720 10746 4729
rect 10324 4684 10376 4690
rect 10690 4655 10692 4664
rect 10324 4626 10376 4632
rect 10744 4655 10746 4664
rect 10692 4626 10744 4632
rect 10336 4282 10364 4626
rect 10704 4282 10732 4626
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10336 4078 10364 4218
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10782 3088 10838 3097
rect 10782 3023 10838 3032
rect 10796 2990 10824 3023
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10336 2689 10364 2790
rect 10322 2680 10378 2689
rect 10322 2615 10378 2624
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 11072 480 11100 3946
rect 11348 3602 11376 12650
rect 11440 11898 11468 18634
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11532 17746 11560 18226
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11532 17338 11560 17682
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11992 16182 12020 20266
rect 12084 20262 12112 20810
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 12084 18442 12112 20198
rect 12176 18578 12204 23462
rect 12268 18698 12296 26862
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12176 18550 12296 18578
rect 12084 18414 12204 18442
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11992 15638 12020 15914
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11716 14890 11744 15438
rect 11808 15162 11836 15574
rect 11992 15502 12020 15574
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11808 14958 11836 15098
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 12176 12753 12204 18414
rect 12162 12744 12218 12753
rect 12162 12679 12218 12688
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11440 10810 11468 11222
rect 11612 11144 11664 11150
rect 11610 11112 11612 11121
rect 11664 11112 11666 11121
rect 11520 11076 11572 11082
rect 11610 11047 11666 11056
rect 11520 11018 11572 11024
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11440 10577 11468 10746
rect 11426 10568 11482 10577
rect 11426 10503 11482 10512
rect 11532 10470 11560 11018
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 10169 11560 10406
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11518 10160 11574 10169
rect 11518 10095 11574 10104
rect 11992 9654 12020 12310
rect 12268 12306 12296 18550
rect 12360 16810 12388 38111
rect 12532 34944 12584 34950
rect 12532 34886 12584 34892
rect 12438 34776 12494 34785
rect 12438 34711 12494 34720
rect 12452 34542 12480 34711
rect 12440 34536 12492 34542
rect 12440 34478 12492 34484
rect 12544 33522 12572 34886
rect 12820 34649 12848 39520
rect 13740 35737 13768 39520
rect 14568 37754 14596 39520
rect 14568 37726 14688 37754
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 13726 35728 13782 35737
rect 13726 35663 13782 35672
rect 14660 35465 14688 37726
rect 13174 35456 13230 35465
rect 13174 35391 13230 35400
rect 14646 35456 14702 35465
rect 14646 35391 14702 35400
rect 13188 35290 13216 35391
rect 13176 35284 13228 35290
rect 13176 35226 13228 35232
rect 13084 35148 13136 35154
rect 13084 35090 13136 35096
rect 12806 34640 12862 34649
rect 12806 34575 12862 34584
rect 13096 34542 13124 35090
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 13634 34504 13690 34513
rect 12806 33552 12862 33561
rect 12532 33516 12584 33522
rect 12806 33487 12808 33496
rect 12532 33458 12584 33464
rect 12860 33487 12862 33496
rect 12808 33458 12860 33464
rect 12544 33114 12572 33458
rect 12532 33108 12584 33114
rect 12532 33050 12584 33056
rect 12438 33008 12494 33017
rect 13096 32978 13124 34478
rect 13634 34439 13690 34448
rect 13174 34232 13230 34241
rect 13174 34167 13176 34176
rect 13228 34167 13230 34176
rect 13176 34138 13228 34144
rect 13452 34060 13504 34066
rect 13452 34002 13504 34008
rect 13464 33658 13492 34002
rect 13452 33652 13504 33658
rect 13452 33594 13504 33600
rect 12438 32943 12494 32952
rect 13084 32972 13136 32978
rect 12452 32570 12480 32943
rect 13084 32914 13136 32920
rect 12440 32564 12492 32570
rect 12440 32506 12492 32512
rect 13096 32230 13124 32914
rect 13084 32224 13136 32230
rect 13084 32166 13136 32172
rect 12714 30832 12770 30841
rect 12714 30767 12770 30776
rect 12532 27328 12584 27334
rect 12532 27270 12584 27276
rect 12440 26512 12492 26518
rect 12440 26454 12492 26460
rect 12452 25702 12480 26454
rect 12544 25906 12572 27270
rect 12728 26874 12756 30767
rect 12806 27568 12862 27577
rect 12806 27503 12808 27512
rect 12860 27503 12862 27512
rect 12808 27474 12860 27480
rect 12820 27130 12848 27474
rect 12990 27160 13046 27169
rect 12808 27124 12860 27130
rect 12990 27095 13046 27104
rect 12808 27066 12860 27072
rect 12728 26846 12848 26874
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12624 26580 12676 26586
rect 12624 26522 12676 26528
rect 12636 25906 12664 26522
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 12544 25498 12572 25842
rect 12440 25492 12492 25498
rect 12440 25434 12492 25440
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12452 23746 12480 25434
rect 12728 25362 12756 26726
rect 12820 26382 12848 26846
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12912 26489 12940 26522
rect 12898 26480 12954 26489
rect 12898 26415 12954 26424
rect 12808 26376 12860 26382
rect 12808 26318 12860 26324
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12532 24880 12584 24886
rect 12532 24822 12584 24828
rect 12544 24750 12572 24822
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12900 24744 12952 24750
rect 12900 24686 12952 24692
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12544 24313 12572 24550
rect 12912 24410 12940 24686
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 12530 24304 12586 24313
rect 12530 24239 12586 24248
rect 12624 24268 12676 24274
rect 12624 24210 12676 24216
rect 12530 23760 12586 23769
rect 12452 23718 12530 23746
rect 12530 23695 12586 23704
rect 12544 22778 12572 23695
rect 12636 23662 12664 24210
rect 12912 24177 12940 24346
rect 13004 24342 13032 27095
rect 12992 24336 13044 24342
rect 12992 24278 13044 24284
rect 12898 24168 12954 24177
rect 12898 24103 12954 24112
rect 12624 23656 12676 23662
rect 12622 23624 12624 23633
rect 12676 23624 12678 23633
rect 12622 23559 12678 23568
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 12544 22166 12572 22510
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 12624 21616 12676 21622
rect 12622 21584 12624 21593
rect 12676 21584 12678 21593
rect 12622 21519 12678 21528
rect 13096 20210 13124 32166
rect 13648 27130 13676 34439
rect 15488 34241 15516 39520
rect 15474 34232 15530 34241
rect 15474 34167 15530 34176
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 13636 27124 13688 27130
rect 13636 27066 13688 27072
rect 13266 26888 13322 26897
rect 13266 26823 13322 26832
rect 13280 25498 13308 26823
rect 13360 26512 13412 26518
rect 13360 26454 13412 26460
rect 13372 25702 13400 26454
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 13360 25696 13412 25702
rect 13360 25638 13412 25644
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13372 24886 13400 25638
rect 13452 25356 13504 25362
rect 13452 25298 13504 25304
rect 13464 25265 13492 25298
rect 13450 25256 13506 25265
rect 13450 25191 13506 25200
rect 13464 24954 13492 25191
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 13452 24948 13504 24954
rect 13452 24890 13504 24896
rect 13360 24880 13412 24886
rect 13360 24822 13412 24828
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 13452 22568 13504 22574
rect 13450 22536 13452 22545
rect 13504 22536 13506 22545
rect 13450 22471 13506 22480
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 13004 20182 13124 20210
rect 12438 18728 12494 18737
rect 12438 18663 12494 18672
rect 12452 18222 12480 18663
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12622 18184 12678 18193
rect 12622 18119 12678 18128
rect 12636 18086 12664 18119
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12820 17338 12848 17682
rect 13004 17649 13032 20182
rect 13082 19952 13138 19961
rect 13082 19887 13138 19896
rect 13096 18834 13124 19887
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13096 17746 13124 18770
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12990 17640 13046 17649
rect 12900 17604 12952 17610
rect 12990 17575 13046 17584
rect 12900 17546 12952 17552
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12360 16794 12480 16810
rect 12360 16788 12492 16794
rect 12360 16782 12440 16788
rect 12440 16730 12492 16736
rect 12820 16726 12848 17274
rect 12912 16998 12940 17546
rect 13096 17270 13124 17682
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12808 16720 12860 16726
rect 12912 16697 12940 16934
rect 12808 16662 12860 16668
rect 12898 16688 12954 16697
rect 12440 16652 12492 16658
rect 12898 16623 12954 16632
rect 13544 16652 13596 16658
rect 12440 16594 12492 16600
rect 13544 16594 13596 16600
rect 12346 16008 12402 16017
rect 12346 15943 12402 15952
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12268 11558 12296 12242
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11428 7336 11480 7342
rect 11426 7304 11428 7313
rect 11480 7304 11482 7313
rect 11426 7239 11482 7248
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11348 3194 11376 3538
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11348 2825 11376 3130
rect 11334 2816 11390 2825
rect 11334 2751 11390 2760
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 12084 2650 12112 11494
rect 12360 5273 12388 15943
rect 12452 15910 12480 16594
rect 13556 16250 13584 16594
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 12374 12480 15846
rect 13556 15638 13584 16186
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 12346 5264 12402 5273
rect 12346 5199 12402 5208
rect 13174 4312 13230 4321
rect 13174 4247 13230 4256
rect 12806 2952 12862 2961
rect 12806 2887 12862 2896
rect 12346 2816 12402 2825
rect 12346 2751 12402 2760
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11900 480 11928 2314
rect 12360 2310 12388 2751
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12820 480 12848 2887
rect 13188 2514 13216 4247
rect 13726 4176 13782 4185
rect 13726 4111 13782 4120
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 13740 480 13768 4111
rect 13832 1873 13860 9590
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 15474 2816 15530 2825
rect 15474 2751 15530 2760
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 13818 1864 13874 1873
rect 13818 1799 13874 1808
rect 14200 1170 14228 2314
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14200 1142 14596 1170
rect 14568 480 14596 1142
rect 15488 480 15516 2751
rect 386 0 442 480
rect 1214 0 1270 480
rect 2134 0 2190 480
rect 3054 0 3110 480
rect 3882 0 3938 480
rect 4802 0 4858 480
rect 5722 0 5778 480
rect 6550 0 6606 480
rect 7470 0 7526 480
rect 8390 0 8446 480
rect 9218 0 9274 480
rect 10138 0 10194 480
rect 11058 0 11114 480
rect 11886 0 11942 480
rect 12806 0 12862 480
rect 13726 0 13782 480
rect 14554 0 14610 480
rect 15474 0 15530 480
<< via2 >>
rect 386 34992 442 35048
rect 1214 34584 1270 34640
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3054 35536 3110 35592
rect 4066 37440 4122 37496
rect 3974 35128 4030 35184
rect 4710 34992 4766 35048
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 4158 34584 4214 34640
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 2686 25200 2742 25256
rect 3146 25744 3202 25800
rect 2962 25356 3018 25392
rect 2962 25336 2964 25356
rect 2964 25336 3016 25356
rect 3016 25336 3018 25356
rect 3146 24656 3202 24712
rect 1398 19216 1454 19272
rect 2870 19216 2926 19272
rect 1674 13912 1730 13968
rect 386 8200 442 8256
rect 2778 19080 2834 19136
rect 2870 17992 2926 18048
rect 2502 17040 2558 17096
rect 2410 9560 2466 9616
rect 3146 23704 3202 23760
rect 3974 27376 4030 27432
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 4066 26968 4122 27024
rect 4894 34720 4950 34776
rect 5354 34992 5410 35048
rect 5262 33396 5264 33416
rect 5264 33396 5316 33416
rect 5316 33396 5318 33416
rect 5262 33360 5318 33396
rect 5262 30368 5318 30424
rect 5354 29028 5410 29064
rect 5354 29008 5356 29028
rect 5356 29008 5408 29028
rect 5408 29008 5410 29028
rect 4526 27376 4582 27432
rect 3974 25880 4030 25936
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 4342 24112 4398 24168
rect 3238 19252 3240 19272
rect 3240 19252 3292 19272
rect 3292 19252 3294 19272
rect 3238 19216 3294 19252
rect 3054 17212 3056 17232
rect 3056 17212 3108 17232
rect 3108 17212 3110 17232
rect 3054 17176 3110 17212
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 4066 22480 4122 22536
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3422 20304 3478 20360
rect 3882 19896 3938 19952
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 4250 20440 4306 20496
rect 3330 17856 3386 17912
rect 3238 17448 3294 17504
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3882 13232 3938 13288
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3054 12436 3110 12472
rect 3054 12416 3056 12436
rect 3056 12416 3108 12436
rect 3108 12416 3110 12436
rect 3054 12144 3110 12200
rect 2778 7384 2834 7440
rect 3054 10240 3110 10296
rect 2502 6196 2504 6216
rect 2504 6196 2556 6216
rect 2556 6196 2558 6216
rect 2502 6160 2558 6196
rect 2410 4936 2466 4992
rect 2134 3712 2190 3768
rect 1398 2488 1454 2544
rect 2318 3596 2374 3632
rect 2318 3576 2320 3596
rect 2320 3576 2372 3596
rect 2372 3576 2374 3596
rect 2318 2624 2374 2680
rect 2870 5072 2926 5128
rect 2502 3476 2504 3496
rect 2504 3476 2556 3496
rect 2556 3476 2558 3496
rect 2502 3440 2558 3476
rect 2962 3712 3018 3768
rect 3238 9560 3294 9616
rect 3146 6840 3202 6896
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 4434 18028 4436 18048
rect 4436 18028 4488 18048
rect 4488 18028 4490 18048
rect 4434 17992 4490 18028
rect 4158 17584 4214 17640
rect 4250 15408 4306 15464
rect 3974 11600 4030 11656
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3882 10648 3938 10704
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 4802 17720 4858 17776
rect 5078 17856 5134 17912
rect 4618 12280 4674 12336
rect 4526 10240 4582 10296
rect 4802 12416 4858 12472
rect 4618 9832 4674 9888
rect 3422 7112 3478 7168
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 4526 8200 4582 8256
rect 4434 7928 4490 7984
rect 3238 4664 3294 4720
rect 3330 3848 3386 3904
rect 3238 3576 3294 3632
rect 3054 3032 3110 3088
rect 3422 3576 3478 3632
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3790 4120 3846 4176
rect 3698 4004 3754 4040
rect 3698 3984 3700 4004
rect 3700 3984 3752 4004
rect 3752 3984 3754 4004
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 4342 3712 4398 3768
rect 3238 2896 3294 2952
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 5078 15136 5134 15192
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 5998 35128 6054 35184
rect 5814 34620 5816 34640
rect 5816 34620 5868 34640
rect 5868 34620 5870 34640
rect 5814 34584 5870 34620
rect 7010 35708 7012 35728
rect 7012 35708 7064 35728
rect 7064 35708 7066 35728
rect 7010 35672 7066 35708
rect 7470 35128 7526 35184
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 5814 31884 5870 31920
rect 5814 31864 5816 31884
rect 5816 31864 5868 31884
rect 5868 31864 5870 31884
rect 5906 30640 5962 30696
rect 5814 27104 5870 27160
rect 5446 22888 5502 22944
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 8114 35028 8116 35048
rect 8116 35028 8168 35048
rect 8168 35028 8170 35048
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8114 34992 8170 35028
rect 7562 34720 7618 34776
rect 6918 31728 6974 31784
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 6734 30640 6790 30696
rect 7010 30368 7066 30424
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6366 28620 6422 28656
rect 6366 28600 6368 28620
rect 6368 28600 6420 28620
rect 6420 28600 6422 28620
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6090 27240 6146 27296
rect 8482 32408 8538 32464
rect 8022 31728 8078 31784
rect 7746 29008 7802 29064
rect 7930 29044 7932 29064
rect 7932 29044 7984 29064
rect 7984 29044 7986 29064
rect 7930 29008 7986 29044
rect 7378 27548 7380 27568
rect 7380 27548 7432 27568
rect 7432 27548 7434 27568
rect 7378 27512 7434 27548
rect 7194 27376 7250 27432
rect 5906 25336 5962 25392
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6918 26988 6974 27024
rect 6918 26968 6920 26988
rect 6920 26968 6972 26988
rect 6972 26968 6974 26988
rect 6918 25916 6920 25936
rect 6920 25916 6972 25936
rect 6972 25916 6974 25936
rect 6918 25880 6974 25916
rect 6642 24928 6698 24984
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6274 23604 6276 23624
rect 6276 23604 6328 23624
rect 6328 23604 6330 23624
rect 6274 23568 6330 23604
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 7194 22888 7250 22944
rect 7194 22480 7250 22536
rect 6734 21256 6790 21312
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6182 20440 6238 20496
rect 6918 20324 6974 20360
rect 6918 20304 6920 20324
rect 6920 20304 6972 20324
rect 6972 20304 6974 20324
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 7194 19896 7250 19952
rect 5630 19216 5686 19272
rect 5998 19216 6054 19272
rect 5354 17448 5410 17504
rect 5262 14864 5318 14920
rect 5170 13640 5226 13696
rect 5262 11600 5318 11656
rect 5078 9460 5080 9480
rect 5080 9460 5132 9480
rect 5132 9460 5134 9480
rect 5078 9424 5134 9460
rect 4710 6840 4766 6896
rect 4802 5652 4804 5672
rect 4804 5652 4856 5672
rect 4856 5652 4858 5672
rect 4802 5616 4858 5652
rect 4986 6840 5042 6896
rect 5446 6296 5502 6352
rect 5262 4936 5318 4992
rect 5630 4120 5686 4176
rect 5170 3168 5226 3224
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 7010 17720 7066 17776
rect 6918 17196 6974 17232
rect 6918 17176 6920 17196
rect 6920 17176 6972 17196
rect 6972 17176 6974 17196
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 7194 16788 7250 16824
rect 7194 16768 7196 16788
rect 7196 16768 7248 16788
rect 7248 16768 7250 16788
rect 6642 16632 6698 16688
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6918 15444 6920 15464
rect 6920 15444 6972 15464
rect 6972 15444 6974 15464
rect 6918 15408 6974 15444
rect 6734 15000 6790 15056
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 7286 13912 7342 13968
rect 6090 13640 6146 13696
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6182 13232 6238 13288
rect 6090 12824 6146 12880
rect 5906 4004 5962 4040
rect 5906 3984 5908 4004
rect 5908 3984 5960 4004
rect 5960 3984 5962 4004
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 7102 12164 7158 12200
rect 7102 12144 7104 12164
rect 7104 12144 7156 12164
rect 7156 12144 7158 12164
rect 7010 11736 7066 11792
rect 6182 11600 6238 11656
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6550 9580 6606 9616
rect 6550 9560 6552 9580
rect 6552 9560 6604 9580
rect 6604 9560 6606 9580
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6182 7928 6238 7984
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6090 3848 6146 3904
rect 5906 3476 5908 3496
rect 5908 3476 5960 3496
rect 5960 3476 5962 3496
rect 5906 3440 5962 3476
rect 5722 3304 5778 3360
rect 4986 2624 5042 2680
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 7010 6160 7066 6216
rect 7102 5752 7158 5808
rect 8390 30676 8392 30696
rect 8392 30676 8444 30696
rect 8444 30676 8446 30696
rect 8390 30640 8446 30676
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8942 32444 8944 32464
rect 8944 32444 8996 32464
rect 8996 32444 8998 32464
rect 8942 32408 8998 32444
rect 8298 28620 8354 28656
rect 8298 28600 8300 28620
rect 8300 28600 8352 28620
rect 8352 28600 8354 28620
rect 8390 27532 8446 27568
rect 8390 27512 8392 27532
rect 8392 27512 8444 27532
rect 8444 27512 8446 27532
rect 8298 27104 8354 27160
rect 7562 25200 7618 25256
rect 7562 23432 7618 23488
rect 7562 23024 7618 23080
rect 8114 21528 8170 21584
rect 7562 14864 7618 14920
rect 7562 13796 7618 13832
rect 7562 13776 7564 13796
rect 7564 13776 7616 13796
rect 7616 13776 7618 13796
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8758 30132 8760 30152
rect 8760 30132 8812 30152
rect 8812 30132 8814 30152
rect 8758 30096 8814 30132
rect 8298 24656 8354 24712
rect 8390 21392 8446 21448
rect 8298 21292 8300 21312
rect 8300 21292 8352 21312
rect 8352 21292 8354 21312
rect 8298 21256 8354 21292
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 9770 35536 9826 35592
rect 10690 34720 10746 34776
rect 10138 30776 10194 30832
rect 10414 28872 10470 28928
rect 9586 27376 9642 27432
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8758 25336 8814 25392
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 9218 24792 9274 24848
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8942 23432 8998 23488
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8666 22480 8722 22536
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8206 17448 8262 17504
rect 8022 17040 8078 17096
rect 8482 16632 8538 16688
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 9218 18808 9274 18864
rect 8942 18672 8998 18728
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 7838 12416 7894 12472
rect 7930 12280 7986 12336
rect 7470 6316 7526 6352
rect 7470 6296 7472 6316
rect 7472 6296 7524 6316
rect 7524 6296 7526 6316
rect 7102 5616 7158 5672
rect 6826 5108 6828 5128
rect 6828 5108 6880 5128
rect 6880 5108 6882 5128
rect 6826 5072 6882 5108
rect 7010 4120 7066 4176
rect 8298 15156 8354 15192
rect 8298 15136 8300 15156
rect 8300 15136 8352 15156
rect 8352 15136 8354 15156
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 9770 27104 9826 27160
rect 9678 26852 9734 26888
rect 9678 26832 9680 26852
rect 9680 26832 9732 26852
rect 9732 26832 9734 26852
rect 10138 26424 10194 26480
rect 10046 25780 10048 25800
rect 10048 25780 10100 25800
rect 10100 25780 10102 25800
rect 10046 25744 10102 25780
rect 9494 24812 9550 24848
rect 9494 24792 9496 24812
rect 9496 24792 9548 24812
rect 9548 24792 9550 24812
rect 9402 24112 9458 24168
rect 9862 24132 9918 24168
rect 9862 24112 9864 24132
rect 9864 24112 9916 24132
rect 9916 24112 9918 24132
rect 9862 23468 9864 23488
rect 9864 23468 9916 23488
rect 9916 23468 9918 23488
rect 9862 23432 9918 23468
rect 9678 23024 9734 23080
rect 9586 22480 9642 22536
rect 9494 21972 9496 21992
rect 9496 21972 9548 21992
rect 9548 21972 9550 21992
rect 9494 21936 9550 21972
rect 9862 21936 9918 21992
rect 9586 20712 9642 20768
rect 10230 23604 10232 23624
rect 10232 23604 10284 23624
rect 10284 23604 10286 23624
rect 10230 23568 10286 23604
rect 10690 31900 10692 31920
rect 10692 31900 10744 31920
rect 10744 31900 10746 31920
rect 10690 31864 10746 31900
rect 12346 38120 12402 38176
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11242 35128 11298 35184
rect 11150 33396 11152 33416
rect 11152 33396 11204 33416
rect 11204 33396 11206 33416
rect 11150 33360 11206 33396
rect 10966 32952 11022 33008
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11518 33496 11574 33552
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 12070 32408 12126 32464
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11058 30640 11114 30696
rect 11058 29008 11114 29064
rect 11426 27512 11482 27568
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 12162 31728 12218 31784
rect 12162 30096 12218 30152
rect 11058 26968 11114 27024
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11058 26152 11114 26208
rect 10598 24656 10654 24712
rect 10322 19624 10378 19680
rect 9586 18148 9642 18184
rect 9586 18128 9588 18148
rect 9588 18128 9640 18148
rect 9640 18128 9642 18148
rect 9494 16632 9550 16688
rect 9402 15972 9458 16008
rect 9402 15952 9404 15972
rect 9404 15952 9456 15972
rect 9456 15952 9458 15972
rect 9770 16768 9826 16824
rect 9954 16652 10010 16688
rect 9954 16632 9956 16652
rect 9956 16632 10008 16652
rect 10008 16632 10010 16652
rect 9678 13776 9734 13832
rect 8114 11192 8170 11248
rect 8390 9460 8392 9480
rect 8392 9460 8444 9480
rect 8444 9460 8446 9480
rect 8390 9424 8446 9460
rect 8758 11056 8814 11112
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 9862 11228 9864 11248
rect 9864 11228 9916 11248
rect 9916 11228 9918 11248
rect 9862 11192 9918 11228
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 7286 3984 7342 4040
rect 7930 4664 7986 4720
rect 6642 3440 6698 3496
rect 6826 3032 6882 3088
rect 6642 2896 6698 2952
rect 7010 2896 7066 2952
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 6734 2760 6790 2816
rect 7010 2624 7066 2680
rect 7470 3304 7526 3360
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 9494 10532 9550 10568
rect 9494 10512 9496 10532
rect 9496 10512 9548 10532
rect 9548 10512 9550 10532
rect 9586 10104 9642 10160
rect 10966 24284 10968 24304
rect 10968 24284 11020 24304
rect 11020 24284 11022 24304
rect 10966 24248 11022 24284
rect 11150 24792 11206 24848
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11334 23568 11390 23624
rect 10506 17584 10562 17640
rect 9954 9968 10010 10024
rect 9770 7248 9826 7304
rect 10230 6840 10286 6896
rect 9678 6160 9734 6216
rect 9678 5772 9734 5808
rect 9678 5752 9680 5772
rect 9680 5752 9732 5772
rect 9732 5752 9734 5772
rect 9678 4256 9734 4312
rect 9678 3440 9734 3496
rect 9862 3576 9918 3632
rect 11150 21392 11206 21448
rect 11150 20712 11206 20768
rect 11242 18828 11298 18864
rect 11242 18808 11244 18828
rect 11244 18808 11296 18828
rect 11296 18808 11298 18828
rect 10966 16496 11022 16552
rect 11150 16632 11206 16688
rect 10874 15000 10930 15056
rect 10874 11600 10930 11656
rect 10966 10648 11022 10704
rect 12162 23568 12218 23624
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11886 21956 11942 21992
rect 11886 21936 11888 21956
rect 11888 21936 11940 21956
rect 11940 21936 11942 21956
rect 11426 21292 11428 21312
rect 11428 21292 11480 21312
rect 11480 21292 11482 21312
rect 11426 21256 11482 21292
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 12070 23432 12126 23488
rect 11978 20712 12034 20768
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11334 13948 11336 13968
rect 11336 13948 11388 13968
rect 11388 13948 11390 13968
rect 11334 13912 11390 13948
rect 11334 12860 11336 12880
rect 11336 12860 11388 12880
rect 11388 12860 11390 12880
rect 11334 12824 11390 12860
rect 11242 9016 11298 9072
rect 10690 4684 10746 4720
rect 10690 4664 10692 4684
rect 10692 4664 10744 4684
rect 10744 4664 10746 4684
rect 10782 3032 10838 3088
rect 10322 2624 10378 2680
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 12162 12688 12218 12744
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11610 11092 11612 11112
rect 11612 11092 11664 11112
rect 11664 11092 11666 11112
rect 11610 11056 11666 11092
rect 11426 10512 11482 10568
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11518 10104 11574 10160
rect 12438 34720 12494 34776
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 13726 35672 13782 35728
rect 13174 35400 13230 35456
rect 14646 35400 14702 35456
rect 12806 34584 12862 34640
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 12806 33516 12862 33552
rect 12806 33496 12808 33516
rect 12808 33496 12860 33516
rect 12860 33496 12862 33516
rect 12438 32952 12494 33008
rect 13634 34448 13690 34504
rect 13174 34196 13230 34232
rect 13174 34176 13176 34196
rect 13176 34176 13228 34196
rect 13228 34176 13230 34196
rect 12714 30776 12770 30832
rect 12806 27532 12862 27568
rect 12806 27512 12808 27532
rect 12808 27512 12860 27532
rect 12860 27512 12862 27532
rect 12990 27104 13046 27160
rect 12898 26424 12954 26480
rect 12530 24248 12586 24304
rect 12530 23704 12586 23760
rect 12898 24112 12954 24168
rect 12622 23604 12624 23624
rect 12624 23604 12676 23624
rect 12676 23604 12678 23624
rect 12622 23568 12678 23604
rect 12622 21564 12624 21584
rect 12624 21564 12676 21584
rect 12676 21564 12678 21584
rect 12622 21528 12678 21564
rect 15474 34176 15530 34232
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 13266 26832 13322 26888
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 13450 25200 13506 25256
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 13450 22516 13452 22536
rect 13452 22516 13504 22536
rect 13504 22516 13506 22536
rect 13450 22480 13506 22516
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 12438 18672 12494 18728
rect 12622 18128 12678 18184
rect 13082 19896 13138 19952
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 12990 17584 13046 17640
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 12898 16632 12954 16688
rect 12346 15952 12402 16008
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11426 7284 11428 7304
rect 11428 7284 11480 7304
rect 11480 7284 11482 7304
rect 11426 7248 11482 7284
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11334 2760 11390 2816
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 12346 5208 12402 5264
rect 13174 4256 13230 4312
rect 12806 2896 12862 2952
rect 12346 2760 12402 2816
rect 13726 4120 13782 4176
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 15474 2760 15530 2816
rect 13818 1808 13874 1864
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
<< metal3 >>
rect 12341 38178 12407 38181
rect 15520 38178 16000 38208
rect 12341 38176 16000 38178
rect 12341 38120 12346 38176
rect 12402 38120 16000 38176
rect 12341 38118 16000 38120
rect 12341 38115 12407 38118
rect 15520 38088 16000 38118
rect 6277 37568 6597 37569
rect 0 37498 480 37528
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 4061 37498 4127 37501
rect 0 37496 4127 37498
rect 0 37440 4066 37496
rect 4122 37440 4127 37496
rect 0 37438 4127 37440
rect 0 37408 480 37438
rect 4061 37435 4127 37438
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 7005 35730 7071 35733
rect 13721 35730 13787 35733
rect 7005 35728 13787 35730
rect 7005 35672 7010 35728
rect 7066 35672 13726 35728
rect 13782 35672 13787 35728
rect 7005 35670 13787 35672
rect 7005 35667 7071 35670
rect 13721 35667 13787 35670
rect 3049 35594 3115 35597
rect 9765 35594 9831 35597
rect 3049 35592 9831 35594
rect 3049 35536 3054 35592
rect 3110 35536 9770 35592
rect 9826 35536 9831 35592
rect 3049 35534 9831 35536
rect 3049 35531 3115 35534
rect 9765 35531 9831 35534
rect 13169 35458 13235 35461
rect 14641 35458 14707 35461
rect 13169 35456 14707 35458
rect 13169 35400 13174 35456
rect 13230 35400 14646 35456
rect 14702 35400 14707 35456
rect 13169 35398 14707 35400
rect 13169 35395 13235 35398
rect 14641 35395 14707 35398
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 3969 35186 4035 35189
rect 5993 35186 6059 35189
rect 3969 35184 6059 35186
rect 3969 35128 3974 35184
rect 4030 35128 5998 35184
rect 6054 35128 6059 35184
rect 3969 35126 6059 35128
rect 3969 35123 4035 35126
rect 5993 35123 6059 35126
rect 7465 35186 7531 35189
rect 11237 35186 11303 35189
rect 7465 35184 11303 35186
rect 7465 35128 7470 35184
rect 7526 35128 11242 35184
rect 11298 35128 11303 35184
rect 7465 35126 11303 35128
rect 7465 35123 7531 35126
rect 11237 35123 11303 35126
rect 381 35050 447 35053
rect 4705 35050 4771 35053
rect 381 35048 4771 35050
rect 381 34992 386 35048
rect 442 34992 4710 35048
rect 4766 34992 4771 35048
rect 381 34990 4771 34992
rect 381 34987 447 34990
rect 4705 34987 4771 34990
rect 5349 35050 5415 35053
rect 8109 35050 8175 35053
rect 5349 35048 8175 35050
rect 5349 34992 5354 35048
rect 5410 34992 8114 35048
rect 8170 34992 8175 35048
rect 5349 34990 8175 34992
rect 5349 34987 5415 34990
rect 8109 34987 8175 34990
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 4889 34778 4955 34781
rect 7557 34778 7623 34781
rect 4889 34776 7623 34778
rect 4889 34720 4894 34776
rect 4950 34720 7562 34776
rect 7618 34720 7623 34776
rect 4889 34718 7623 34720
rect 4889 34715 4955 34718
rect 7557 34715 7623 34718
rect 10685 34778 10751 34781
rect 12433 34778 12499 34781
rect 10685 34776 12499 34778
rect 10685 34720 10690 34776
rect 10746 34720 12438 34776
rect 12494 34720 12499 34776
rect 10685 34718 12499 34720
rect 10685 34715 10751 34718
rect 12433 34715 12499 34718
rect 1209 34642 1275 34645
rect 4153 34642 4219 34645
rect 1209 34640 4219 34642
rect 1209 34584 1214 34640
rect 1270 34584 4158 34640
rect 4214 34584 4219 34640
rect 1209 34582 4219 34584
rect 1209 34579 1275 34582
rect 4153 34579 4219 34582
rect 5809 34642 5875 34645
rect 12801 34642 12867 34645
rect 5809 34640 12867 34642
rect 5809 34584 5814 34640
rect 5870 34584 12806 34640
rect 12862 34584 12867 34640
rect 5809 34582 12867 34584
rect 5809 34579 5875 34582
rect 12801 34579 12867 34582
rect 13629 34506 13695 34509
rect 15520 34506 16000 34536
rect 13629 34504 16000 34506
rect 13629 34448 13634 34504
rect 13690 34448 16000 34504
rect 13629 34446 16000 34448
rect 13629 34443 13695 34446
rect 15520 34416 16000 34446
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 13169 34234 13235 34237
rect 15469 34234 15535 34237
rect 13169 34232 15535 34234
rect 13169 34176 13174 34232
rect 13230 34176 15474 34232
rect 15530 34176 15535 34232
rect 13169 34174 15535 34176
rect 13169 34171 13235 34174
rect 15469 34171 15535 34174
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 11513 33554 11579 33557
rect 12801 33554 12867 33557
rect 11513 33552 12867 33554
rect 11513 33496 11518 33552
rect 11574 33496 12806 33552
rect 12862 33496 12867 33552
rect 11513 33494 12867 33496
rect 11513 33491 11579 33494
rect 12801 33491 12867 33494
rect 5257 33418 5323 33421
rect 11145 33418 11211 33421
rect 5257 33416 11211 33418
rect 5257 33360 5262 33416
rect 5318 33360 11150 33416
rect 11206 33360 11211 33416
rect 5257 33358 11211 33360
rect 5257 33355 5323 33358
rect 11145 33355 11211 33358
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 10961 33010 11027 33013
rect 12433 33010 12499 33013
rect 10961 33008 12499 33010
rect 10961 32952 10966 33008
rect 11022 32952 12438 33008
rect 12494 32952 12499 33008
rect 10961 32950 12499 32952
rect 10961 32947 11027 32950
rect 12433 32947 12499 32950
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 0 32466 480 32496
rect 8477 32466 8543 32469
rect 0 32464 8543 32466
rect 0 32408 8482 32464
rect 8538 32408 8543 32464
rect 0 32406 8543 32408
rect 0 32376 480 32406
rect 8477 32403 8543 32406
rect 8937 32466 9003 32469
rect 12065 32466 12131 32469
rect 8937 32464 12131 32466
rect 8937 32408 8942 32464
rect 8998 32408 12070 32464
rect 12126 32408 12131 32464
rect 8937 32406 12131 32408
rect 8937 32403 9003 32406
rect 12065 32403 12131 32406
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 5809 31922 5875 31925
rect 10685 31922 10751 31925
rect 5809 31920 10751 31922
rect 5809 31864 5814 31920
rect 5870 31864 10690 31920
rect 10746 31864 10751 31920
rect 5809 31862 10751 31864
rect 5809 31859 5875 31862
rect 10685 31859 10751 31862
rect 6913 31786 6979 31789
rect 8017 31786 8083 31789
rect 12157 31786 12223 31789
rect 6913 31784 12223 31786
rect 6913 31728 6918 31784
rect 6974 31728 8022 31784
rect 8078 31728 12162 31784
rect 12218 31728 12223 31784
rect 6913 31726 12223 31728
rect 6913 31723 6979 31726
rect 8017 31723 8083 31726
rect 12157 31723 12223 31726
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 10133 30834 10199 30837
rect 12709 30834 12775 30837
rect 15520 30834 16000 30864
rect 10133 30832 12775 30834
rect 10133 30776 10138 30832
rect 10194 30776 12714 30832
rect 12770 30776 12775 30832
rect 10133 30774 12775 30776
rect 10133 30771 10199 30774
rect 12709 30771 12775 30774
rect 13862 30774 16000 30834
rect 5901 30698 5967 30701
rect 6729 30698 6795 30701
rect 8385 30698 8451 30701
rect 5901 30696 8451 30698
rect 5901 30640 5906 30696
rect 5962 30640 6734 30696
rect 6790 30640 8390 30696
rect 8446 30640 8451 30696
rect 5901 30638 8451 30640
rect 5901 30635 5967 30638
rect 6729 30635 6795 30638
rect 8385 30635 8451 30638
rect 11053 30698 11119 30701
rect 13862 30698 13922 30774
rect 15520 30744 16000 30774
rect 11053 30696 13922 30698
rect 11053 30640 11058 30696
rect 11114 30640 13922 30696
rect 11053 30638 13922 30640
rect 11053 30635 11119 30638
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 5257 30426 5323 30429
rect 7005 30426 7071 30429
rect 5257 30424 7071 30426
rect 5257 30368 5262 30424
rect 5318 30368 7010 30424
rect 7066 30368 7071 30424
rect 5257 30366 7071 30368
rect 5257 30363 5323 30366
rect 7005 30363 7071 30366
rect 8753 30154 8819 30157
rect 12157 30154 12223 30157
rect 8753 30152 12223 30154
rect 8753 30096 8758 30152
rect 8814 30096 12162 30152
rect 12218 30096 12223 30152
rect 8753 30094 12223 30096
rect 8753 30091 8819 30094
rect 12157 30091 12223 30094
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 5349 29066 5415 29069
rect 7741 29066 7807 29069
rect 5349 29064 7807 29066
rect 5349 29008 5354 29064
rect 5410 29008 7746 29064
rect 7802 29008 7807 29064
rect 5349 29006 7807 29008
rect 5349 29003 5415 29006
rect 7741 29003 7807 29006
rect 7925 29066 7991 29069
rect 11053 29066 11119 29069
rect 7925 29064 11119 29066
rect 7925 29008 7930 29064
rect 7986 29008 11058 29064
rect 11114 29008 11119 29064
rect 7925 29006 11119 29008
rect 7925 29003 7991 29006
rect 11053 29003 11119 29006
rect 10409 28932 10475 28933
rect 10358 28930 10364 28932
rect 10318 28870 10364 28930
rect 10428 28928 10475 28932
rect 10470 28872 10475 28928
rect 10358 28868 10364 28870
rect 10428 28868 10475 28872
rect 10409 28867 10475 28868
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 6361 28658 6427 28661
rect 8293 28658 8359 28661
rect 6361 28656 8359 28658
rect 6361 28600 6366 28656
rect 6422 28600 8298 28656
rect 8354 28600 8359 28656
rect 6361 28598 8359 28600
rect 6361 28595 6427 28598
rect 8293 28595 8359 28598
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 7373 27570 7439 27573
rect 8385 27570 8451 27573
rect 7373 27568 8451 27570
rect 7373 27512 7378 27568
rect 7434 27512 8390 27568
rect 8446 27512 8451 27568
rect 7373 27510 8451 27512
rect 7373 27507 7439 27510
rect 8385 27507 8451 27510
rect 11421 27570 11487 27573
rect 12801 27570 12867 27573
rect 11421 27568 12867 27570
rect 11421 27512 11426 27568
rect 11482 27512 12806 27568
rect 12862 27512 12867 27568
rect 11421 27510 12867 27512
rect 11421 27507 11487 27510
rect 12801 27507 12867 27510
rect 0 27434 480 27464
rect 3969 27434 4035 27437
rect 0 27432 4035 27434
rect 0 27376 3974 27432
rect 4030 27376 4035 27432
rect 0 27374 4035 27376
rect 0 27344 480 27374
rect 3969 27371 4035 27374
rect 4521 27434 4587 27437
rect 7189 27434 7255 27437
rect 9581 27434 9647 27437
rect 4521 27432 9647 27434
rect 4521 27376 4526 27432
rect 4582 27376 7194 27432
rect 7250 27376 9586 27432
rect 9642 27376 9647 27432
rect 4521 27374 9647 27376
rect 4521 27371 4587 27374
rect 7189 27371 7255 27374
rect 9581 27371 9647 27374
rect 6085 27300 6151 27301
rect 6085 27298 6132 27300
rect 6040 27296 6132 27298
rect 6196 27298 6202 27300
rect 15520 27298 16000 27328
rect 6040 27240 6090 27296
rect 6040 27238 6132 27240
rect 6085 27236 6132 27238
rect 6196 27238 8770 27298
rect 6196 27236 6202 27238
rect 6085 27235 6151 27236
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 5809 27162 5875 27165
rect 8293 27162 8359 27165
rect 5809 27160 8359 27162
rect 5809 27104 5814 27160
rect 5870 27104 8298 27160
rect 8354 27104 8359 27160
rect 5809 27102 8359 27104
rect 5809 27099 5875 27102
rect 8293 27099 8359 27102
rect 4061 27026 4127 27029
rect 6913 27026 6979 27029
rect 4061 27024 6979 27026
rect 4061 26968 4066 27024
rect 4122 26968 6918 27024
rect 6974 26968 6979 27024
rect 4061 26966 6979 26968
rect 8710 27026 8770 27238
rect 14782 27238 16000 27298
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 9765 27162 9831 27165
rect 12985 27162 13051 27165
rect 9765 27160 13051 27162
rect 9765 27104 9770 27160
rect 9826 27104 12990 27160
rect 13046 27104 13051 27160
rect 9765 27102 13051 27104
rect 9765 27099 9831 27102
rect 12985 27099 13051 27102
rect 11053 27026 11119 27029
rect 8710 27024 11119 27026
rect 8710 26968 11058 27024
rect 11114 26968 11119 27024
rect 8710 26966 11119 26968
rect 4061 26963 4127 26966
rect 6913 26963 6979 26966
rect 11053 26963 11119 26966
rect 9673 26890 9739 26893
rect 13261 26890 13327 26893
rect 9673 26888 13327 26890
rect 9673 26832 9678 26888
rect 9734 26832 13266 26888
rect 13322 26832 13327 26888
rect 9673 26830 13327 26832
rect 9673 26827 9739 26830
rect 13261 26827 13327 26830
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 10133 26482 10199 26485
rect 12893 26482 12959 26485
rect 10133 26480 12959 26482
rect 10133 26424 10138 26480
rect 10194 26424 12898 26480
rect 12954 26424 12959 26480
rect 10133 26422 12959 26424
rect 10133 26419 10199 26422
rect 12893 26419 12959 26422
rect 14782 26346 14842 27238
rect 15520 27208 16000 27238
rect 11102 26286 14842 26346
rect 11102 26213 11162 26286
rect 11053 26208 11162 26213
rect 11053 26152 11058 26208
rect 11114 26152 11162 26208
rect 11053 26150 11162 26152
rect 11053 26147 11119 26150
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 3969 25938 4035 25941
rect 6913 25938 6979 25941
rect 3969 25936 6979 25938
rect 3969 25880 3974 25936
rect 4030 25880 6918 25936
rect 6974 25880 6979 25936
rect 3969 25878 6979 25880
rect 3969 25875 4035 25878
rect 6913 25875 6979 25878
rect 3141 25802 3207 25805
rect 10041 25802 10107 25805
rect 3141 25800 10107 25802
rect 3141 25744 3146 25800
rect 3202 25744 10046 25800
rect 10102 25744 10107 25800
rect 3141 25742 10107 25744
rect 3141 25739 3207 25742
rect 10041 25739 10107 25742
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 2957 25394 3023 25397
rect 5901 25394 5967 25397
rect 8753 25394 8819 25397
rect 2957 25392 8819 25394
rect 2957 25336 2962 25392
rect 3018 25336 5906 25392
rect 5962 25336 8758 25392
rect 8814 25336 8819 25392
rect 2957 25334 8819 25336
rect 2957 25331 3023 25334
rect 5901 25331 5967 25334
rect 8753 25331 8819 25334
rect 2681 25258 2747 25261
rect 7557 25258 7623 25261
rect 13445 25258 13511 25261
rect 2681 25256 7623 25258
rect 2681 25200 2686 25256
rect 2742 25200 7562 25256
rect 7618 25200 7623 25256
rect 2681 25198 7623 25200
rect 2681 25195 2747 25198
rect 7557 25195 7623 25198
rect 8710 25256 13511 25258
rect 8710 25200 13450 25256
rect 13506 25200 13511 25256
rect 8710 25198 13511 25200
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 6637 24986 6703 24989
rect 8710 24986 8770 25198
rect 13445 25195 13511 25198
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 6637 24984 8770 24986
rect 6637 24928 6642 24984
rect 6698 24928 8770 24984
rect 6637 24926 8770 24928
rect 6637 24923 6703 24926
rect 8710 24850 8770 24926
rect 9213 24850 9279 24853
rect 8710 24848 9279 24850
rect 8710 24792 9218 24848
rect 9274 24792 9279 24848
rect 8710 24790 9279 24792
rect 9213 24787 9279 24790
rect 9489 24850 9555 24853
rect 11145 24850 11211 24853
rect 9489 24848 11211 24850
rect 9489 24792 9494 24848
rect 9550 24792 11150 24848
rect 11206 24792 11211 24848
rect 9489 24790 11211 24792
rect 9489 24787 9555 24790
rect 11145 24787 11211 24790
rect 3141 24714 3207 24717
rect 8293 24714 8359 24717
rect 10593 24714 10659 24717
rect 3141 24712 10659 24714
rect 3141 24656 3146 24712
rect 3202 24656 8298 24712
rect 8354 24656 10598 24712
rect 10654 24656 10659 24712
rect 3141 24654 10659 24656
rect 3141 24651 3207 24654
rect 8293 24651 8359 24654
rect 10593 24651 10659 24654
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 10961 24306 11027 24309
rect 12525 24306 12591 24309
rect 10961 24304 12591 24306
rect 10961 24248 10966 24304
rect 11022 24248 12530 24304
rect 12586 24248 12591 24304
rect 10961 24246 12591 24248
rect 10961 24243 11027 24246
rect 12525 24243 12591 24246
rect 4337 24170 4403 24173
rect 9397 24170 9463 24173
rect 9857 24170 9923 24173
rect 12893 24170 12959 24173
rect 4337 24168 12959 24170
rect 4337 24112 4342 24168
rect 4398 24112 9402 24168
rect 9458 24112 9862 24168
rect 9918 24112 12898 24168
rect 12954 24112 12959 24168
rect 4337 24110 12959 24112
rect 4337 24107 4403 24110
rect 9397 24107 9463 24110
rect 9857 24107 9923 24110
rect 12893 24107 12959 24110
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 3141 23762 3207 23765
rect 12525 23762 12591 23765
rect 3141 23760 12591 23762
rect 3141 23704 3146 23760
rect 3202 23704 12530 23760
rect 12586 23704 12591 23760
rect 3141 23702 12591 23704
rect 3141 23699 3207 23702
rect 12525 23699 12591 23702
rect 6269 23626 6335 23629
rect 10225 23626 10291 23629
rect 6269 23624 10291 23626
rect 6269 23568 6274 23624
rect 6330 23568 10230 23624
rect 10286 23568 10291 23624
rect 6269 23566 10291 23568
rect 6269 23563 6335 23566
rect 10225 23563 10291 23566
rect 11329 23626 11395 23629
rect 12157 23626 12223 23629
rect 12617 23626 12683 23629
rect 15520 23626 16000 23656
rect 11329 23624 12683 23626
rect 11329 23568 11334 23624
rect 11390 23568 12162 23624
rect 12218 23568 12622 23624
rect 12678 23568 12683 23624
rect 11329 23566 12683 23568
rect 11329 23563 11395 23566
rect 12157 23563 12223 23566
rect 12617 23563 12683 23566
rect 13862 23566 16000 23626
rect 7557 23490 7623 23493
rect 8937 23490 9003 23493
rect 9857 23490 9923 23493
rect 7557 23488 9923 23490
rect 7557 23432 7562 23488
rect 7618 23432 8942 23488
rect 8998 23432 9862 23488
rect 9918 23432 9923 23488
rect 7557 23430 9923 23432
rect 7557 23427 7623 23430
rect 8937 23427 9003 23430
rect 9857 23427 9923 23430
rect 12065 23490 12131 23493
rect 13862 23490 13922 23566
rect 15520 23536 16000 23566
rect 12065 23488 13922 23490
rect 12065 23432 12070 23488
rect 12126 23432 13922 23488
rect 12065 23430 13922 23432
rect 12065 23427 12131 23430
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 7557 23082 7623 23085
rect 9673 23082 9739 23085
rect 7557 23080 9739 23082
rect 7557 23024 7562 23080
rect 7618 23024 9678 23080
rect 9734 23024 9739 23080
rect 7557 23022 9739 23024
rect 7557 23019 7623 23022
rect 9673 23019 9739 23022
rect 5441 22946 5507 22949
rect 7189 22946 7255 22949
rect 5441 22944 7255 22946
rect 5441 22888 5446 22944
rect 5502 22888 7194 22944
rect 7250 22888 7255 22944
rect 5441 22886 7255 22888
rect 5441 22883 5507 22886
rect 7189 22883 7255 22886
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 0 22538 480 22568
rect 4061 22538 4127 22541
rect 0 22536 4127 22538
rect 0 22480 4066 22536
rect 4122 22480 4127 22536
rect 0 22478 4127 22480
rect 0 22448 480 22478
rect 4061 22475 4127 22478
rect 7189 22538 7255 22541
rect 8661 22538 8727 22541
rect 7189 22536 8727 22538
rect 7189 22480 7194 22536
rect 7250 22480 8666 22536
rect 8722 22480 8727 22536
rect 7189 22478 8727 22480
rect 7189 22475 7255 22478
rect 8661 22475 8727 22478
rect 9581 22538 9647 22541
rect 13445 22538 13511 22541
rect 9581 22536 13511 22538
rect 9581 22480 9586 22536
rect 9642 22480 13450 22536
rect 13506 22480 13511 22536
rect 9581 22478 13511 22480
rect 9581 22475 9647 22478
rect 13445 22475 13511 22478
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 9489 21994 9555 21997
rect 9857 21994 9923 21997
rect 11881 21994 11947 21997
rect 9489 21992 11947 21994
rect 9489 21936 9494 21992
rect 9550 21936 9862 21992
rect 9918 21936 11886 21992
rect 11942 21936 11947 21992
rect 9489 21934 11947 21936
rect 9489 21931 9555 21934
rect 9857 21931 9923 21934
rect 11881 21931 11947 21934
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 8109 21586 8175 21589
rect 12617 21586 12683 21589
rect 8109 21584 12683 21586
rect 8109 21528 8114 21584
rect 8170 21528 12622 21584
rect 12678 21528 12683 21584
rect 8109 21526 12683 21528
rect 8109 21523 8175 21526
rect 12617 21523 12683 21526
rect 8385 21450 8451 21453
rect 11145 21450 11211 21453
rect 8385 21448 11211 21450
rect 8385 21392 8390 21448
rect 8446 21392 11150 21448
rect 11206 21392 11211 21448
rect 8385 21390 11211 21392
rect 8385 21387 8451 21390
rect 11145 21387 11211 21390
rect 6729 21314 6795 21317
rect 8293 21314 8359 21317
rect 11421 21314 11487 21317
rect 6729 21312 11487 21314
rect 6729 21256 6734 21312
rect 6790 21256 8298 21312
rect 8354 21256 11426 21312
rect 11482 21256 11487 21312
rect 6729 21254 11487 21256
rect 6729 21251 6795 21254
rect 8293 21251 8359 21254
rect 11421 21251 11487 21254
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 9581 20770 9647 20773
rect 11145 20770 11211 20773
rect 11973 20770 12039 20773
rect 9581 20768 12039 20770
rect 9581 20712 9586 20768
rect 9642 20712 11150 20768
rect 11206 20712 11978 20768
rect 12034 20712 12039 20768
rect 9581 20710 12039 20712
rect 9581 20707 9647 20710
rect 11145 20707 11211 20710
rect 11973 20707 12039 20710
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 4245 20498 4311 20501
rect 6177 20498 6243 20501
rect 4245 20496 6243 20498
rect 4245 20440 4250 20496
rect 4306 20440 6182 20496
rect 6238 20440 6243 20496
rect 4245 20438 6243 20440
rect 4245 20435 4311 20438
rect 6177 20435 6243 20438
rect 3417 20362 3483 20365
rect 6913 20362 6979 20365
rect 3417 20360 6979 20362
rect 3417 20304 3422 20360
rect 3478 20304 6918 20360
rect 6974 20304 6979 20360
rect 3417 20302 6979 20304
rect 3417 20299 3483 20302
rect 6913 20299 6979 20302
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 3877 19954 3943 19957
rect 7189 19954 7255 19957
rect 3877 19952 7255 19954
rect 3877 19896 3882 19952
rect 3938 19896 7194 19952
rect 7250 19896 7255 19952
rect 3877 19894 7255 19896
rect 3877 19891 3943 19894
rect 7189 19891 7255 19894
rect 13077 19954 13143 19957
rect 15520 19954 16000 19984
rect 13077 19952 16000 19954
rect 13077 19896 13082 19952
rect 13138 19896 16000 19952
rect 13077 19894 16000 19896
rect 13077 19891 13143 19894
rect 15520 19864 16000 19894
rect 10317 19684 10383 19685
rect 10317 19682 10364 19684
rect 10272 19680 10364 19682
rect 10272 19624 10322 19680
rect 10272 19622 10364 19624
rect 10317 19620 10364 19622
rect 10428 19620 10434 19684
rect 10317 19619 10383 19620
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 1393 19274 1459 19277
rect 2865 19274 2931 19277
rect 1393 19272 2931 19274
rect 1393 19216 1398 19272
rect 1454 19216 2870 19272
rect 2926 19216 2931 19272
rect 1393 19214 2931 19216
rect 1393 19211 1459 19214
rect 2865 19211 2931 19214
rect 3233 19274 3299 19277
rect 5625 19274 5691 19277
rect 3233 19272 5691 19274
rect 3233 19216 3238 19272
rect 3294 19216 5630 19272
rect 5686 19216 5691 19272
rect 3233 19214 5691 19216
rect 3233 19211 3299 19214
rect 5625 19211 5691 19214
rect 5993 19274 6059 19277
rect 6126 19274 6132 19276
rect 5993 19272 6132 19274
rect 5993 19216 5998 19272
rect 6054 19216 6132 19272
rect 5993 19214 6132 19216
rect 5993 19211 6059 19214
rect 6126 19212 6132 19214
rect 6196 19212 6202 19276
rect 2773 19138 2839 19141
rect 3236 19138 3296 19211
rect 2773 19136 3296 19138
rect 2773 19080 2778 19136
rect 2834 19080 3296 19136
rect 2773 19078 3296 19080
rect 2773 19075 2839 19078
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 9213 18866 9279 18869
rect 11237 18866 11303 18869
rect 9213 18864 11303 18866
rect 9213 18808 9218 18864
rect 9274 18808 11242 18864
rect 11298 18808 11303 18864
rect 9213 18806 11303 18808
rect 9213 18803 9279 18806
rect 11237 18803 11303 18806
rect 8937 18730 9003 18733
rect 12433 18730 12499 18733
rect 8937 18728 12499 18730
rect 8937 18672 8942 18728
rect 8998 18672 12438 18728
rect 12494 18672 12499 18728
rect 8937 18670 12499 18672
rect 8937 18667 9003 18670
rect 12433 18667 12499 18670
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 9581 18186 9647 18189
rect 12617 18186 12683 18189
rect 9581 18184 12683 18186
rect 9581 18128 9586 18184
rect 9642 18128 12622 18184
rect 12678 18128 12683 18184
rect 9581 18126 12683 18128
rect 9581 18123 9647 18126
rect 12617 18123 12683 18126
rect 2865 18050 2931 18053
rect 4429 18050 4495 18053
rect 2865 18048 4495 18050
rect 2865 17992 2870 18048
rect 2926 17992 4434 18048
rect 4490 17992 4495 18048
rect 2865 17990 4495 17992
rect 2865 17987 2931 17990
rect 4429 17987 4495 17990
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 3325 17914 3391 17917
rect 5073 17914 5139 17917
rect 3325 17912 5139 17914
rect 3325 17856 3330 17912
rect 3386 17856 5078 17912
rect 5134 17856 5139 17912
rect 3325 17854 5139 17856
rect 3325 17851 3391 17854
rect 5073 17851 5139 17854
rect 4797 17778 4863 17781
rect 7005 17778 7071 17781
rect 4797 17776 7071 17778
rect 4797 17720 4802 17776
rect 4858 17720 7010 17776
rect 7066 17720 7071 17776
rect 4797 17718 7071 17720
rect 4797 17715 4863 17718
rect 7005 17715 7071 17718
rect 4153 17642 4219 17645
rect 10501 17642 10567 17645
rect 12985 17642 13051 17645
rect 4153 17640 13051 17642
rect 4153 17584 4158 17640
rect 4214 17584 10506 17640
rect 10562 17584 12990 17640
rect 13046 17584 13051 17640
rect 4153 17582 13051 17584
rect 4153 17579 4219 17582
rect 10501 17579 10567 17582
rect 12985 17579 13051 17582
rect 0 17506 480 17536
rect 3233 17506 3299 17509
rect 0 17504 3299 17506
rect 0 17448 3238 17504
rect 3294 17448 3299 17504
rect 0 17446 3299 17448
rect 0 17416 480 17446
rect 3233 17443 3299 17446
rect 5349 17506 5415 17509
rect 7046 17506 7052 17508
rect 5349 17504 7052 17506
rect 5349 17448 5354 17504
rect 5410 17448 7052 17504
rect 5349 17446 7052 17448
rect 5349 17443 5415 17446
rect 7046 17444 7052 17446
rect 7116 17506 7122 17508
rect 8201 17506 8267 17509
rect 7116 17504 8267 17506
rect 7116 17448 8206 17504
rect 8262 17448 8267 17504
rect 7116 17446 8267 17448
rect 7116 17444 7122 17446
rect 8201 17443 8267 17446
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 3049 17234 3115 17237
rect 6913 17234 6979 17237
rect 3049 17232 6979 17234
rect 3049 17176 3054 17232
rect 3110 17176 6918 17232
rect 6974 17176 6979 17232
rect 3049 17174 6979 17176
rect 3049 17171 3115 17174
rect 6913 17171 6979 17174
rect 2497 17098 2563 17101
rect 8017 17098 8083 17101
rect 2497 17096 8083 17098
rect 2497 17040 2502 17096
rect 2558 17040 8022 17096
rect 8078 17040 8083 17096
rect 2497 17038 8083 17040
rect 2497 17035 2563 17038
rect 8017 17035 8083 17038
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 7189 16826 7255 16829
rect 9765 16826 9831 16829
rect 7189 16824 9831 16826
rect 7189 16768 7194 16824
rect 7250 16768 9770 16824
rect 9826 16768 9831 16824
rect 7189 16766 9831 16768
rect 7189 16763 7255 16766
rect 9765 16763 9831 16766
rect 6637 16690 6703 16693
rect 8477 16690 8543 16693
rect 6637 16688 8543 16690
rect 6637 16632 6642 16688
rect 6698 16632 8482 16688
rect 8538 16632 8543 16688
rect 6637 16630 8543 16632
rect 6637 16627 6703 16630
rect 8477 16627 8543 16630
rect 9489 16690 9555 16693
rect 9949 16690 10015 16693
rect 11145 16690 11211 16693
rect 9489 16688 11211 16690
rect 9489 16632 9494 16688
rect 9550 16632 9954 16688
rect 10010 16632 11150 16688
rect 11206 16632 11211 16688
rect 9489 16630 11211 16632
rect 9489 16627 9555 16630
rect 9949 16627 10015 16630
rect 11145 16627 11211 16630
rect 12893 16690 12959 16693
rect 12893 16688 13002 16690
rect 12893 16632 12898 16688
rect 12954 16632 13002 16688
rect 12893 16627 13002 16632
rect 10961 16554 11027 16557
rect 12942 16554 13002 16627
rect 10961 16552 14842 16554
rect 10961 16496 10966 16552
rect 11022 16496 14842 16552
rect 10961 16494 14842 16496
rect 10961 16491 11027 16494
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 14782 16282 14842 16494
rect 15520 16282 16000 16312
rect 14782 16222 16000 16282
rect 15520 16192 16000 16222
rect 9397 16010 9463 16013
rect 12341 16010 12407 16013
rect 9397 16008 12407 16010
rect 9397 15952 9402 16008
rect 9458 15952 12346 16008
rect 12402 15952 12407 16008
rect 9397 15950 12407 15952
rect 9397 15947 9463 15950
rect 12341 15947 12407 15950
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 4245 15466 4311 15469
rect 6913 15466 6979 15469
rect 4245 15464 6979 15466
rect 4245 15408 4250 15464
rect 4306 15408 6918 15464
rect 6974 15408 6979 15464
rect 4245 15406 6979 15408
rect 4245 15403 4311 15406
rect 6913 15403 6979 15406
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 5073 15194 5139 15197
rect 8293 15194 8359 15197
rect 5073 15192 8359 15194
rect 5073 15136 5078 15192
rect 5134 15136 8298 15192
rect 8354 15136 8359 15192
rect 5073 15134 8359 15136
rect 5073 15131 5139 15134
rect 8293 15131 8359 15134
rect 6729 15058 6795 15061
rect 10869 15058 10935 15061
rect 6729 15056 10935 15058
rect 6729 15000 6734 15056
rect 6790 15000 10874 15056
rect 10930 15000 10935 15056
rect 6729 14998 10935 15000
rect 6729 14995 6795 14998
rect 10869 14995 10935 14998
rect 5257 14922 5323 14925
rect 7557 14922 7623 14925
rect 5257 14920 7623 14922
rect 5257 14864 5262 14920
rect 5318 14864 7562 14920
rect 7618 14864 7623 14920
rect 5257 14862 7623 14864
rect 5257 14859 5323 14862
rect 7557 14859 7623 14862
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 1669 13970 1735 13973
rect 7281 13970 7347 13973
rect 11329 13970 11395 13973
rect 1669 13968 11395 13970
rect 1669 13912 1674 13968
rect 1730 13912 7286 13968
rect 7342 13912 11334 13968
rect 11390 13912 11395 13968
rect 1669 13910 11395 13912
rect 1669 13907 1735 13910
rect 7281 13907 7347 13910
rect 11329 13907 11395 13910
rect 7557 13834 7623 13837
rect 9673 13834 9739 13837
rect 7557 13832 9739 13834
rect 7557 13776 7562 13832
rect 7618 13776 9678 13832
rect 9734 13776 9739 13832
rect 7557 13774 9739 13776
rect 7557 13771 7623 13774
rect 9673 13771 9739 13774
rect 5165 13698 5231 13701
rect 6085 13698 6151 13701
rect 5165 13696 6151 13698
rect 5165 13640 5170 13696
rect 5226 13640 6090 13696
rect 6146 13640 6151 13696
rect 5165 13638 6151 13640
rect 5165 13635 5231 13638
rect 6085 13635 6151 13638
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3877 13290 3943 13293
rect 6177 13290 6243 13293
rect 3877 13288 6243 13290
rect 3877 13232 3882 13288
rect 3938 13232 6182 13288
rect 6238 13232 6243 13288
rect 3877 13230 6243 13232
rect 3877 13227 3943 13230
rect 6177 13227 6243 13230
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 6085 12882 6151 12885
rect 11329 12882 11395 12885
rect 6085 12880 11395 12882
rect 6085 12824 6090 12880
rect 6146 12824 11334 12880
rect 11390 12824 11395 12880
rect 6085 12822 11395 12824
rect 6085 12819 6151 12822
rect 11329 12819 11395 12822
rect 12157 12746 12223 12749
rect 15520 12746 16000 12776
rect 12157 12744 16000 12746
rect 12157 12688 12162 12744
rect 12218 12688 16000 12744
rect 12157 12686 16000 12688
rect 12157 12683 12223 12686
rect 15520 12656 16000 12686
rect 6277 12544 6597 12545
rect 0 12474 480 12504
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 3049 12474 3115 12477
rect 0 12472 3115 12474
rect 0 12416 3054 12472
rect 3110 12416 3115 12472
rect 0 12414 3115 12416
rect 0 12384 480 12414
rect 3049 12411 3115 12414
rect 4797 12474 4863 12477
rect 7833 12474 7899 12477
rect 4797 12472 4906 12474
rect 4797 12416 4802 12472
rect 4858 12416 4906 12472
rect 4797 12411 4906 12416
rect 4613 12338 4679 12341
rect 4846 12338 4906 12411
rect 4613 12336 4906 12338
rect 4613 12280 4618 12336
rect 4674 12280 4906 12336
rect 4613 12278 4906 12280
rect 7790 12472 7899 12474
rect 7790 12416 7838 12472
rect 7894 12416 7899 12472
rect 7790 12411 7899 12416
rect 7790 12338 7850 12411
rect 7925 12338 7991 12341
rect 7790 12336 7991 12338
rect 7790 12280 7930 12336
rect 7986 12280 7991 12336
rect 7790 12278 7991 12280
rect 4613 12275 4679 12278
rect 7925 12275 7991 12278
rect 3049 12202 3115 12205
rect 7097 12202 7163 12205
rect 3049 12200 7163 12202
rect 3049 12144 3054 12200
rect 3110 12144 7102 12200
rect 7158 12144 7163 12200
rect 3049 12142 7163 12144
rect 3049 12139 3115 12142
rect 7097 12139 7163 12142
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 7005 11796 7071 11797
rect 7005 11792 7052 11796
rect 7116 11794 7122 11796
rect 7005 11736 7010 11792
rect 7005 11732 7052 11736
rect 7116 11734 7162 11794
rect 7116 11732 7122 11734
rect 7005 11731 7071 11732
rect 3969 11658 4035 11661
rect 5257 11658 5323 11661
rect 3969 11656 5323 11658
rect 3969 11600 3974 11656
rect 4030 11600 5262 11656
rect 5318 11600 5323 11656
rect 3969 11598 5323 11600
rect 3969 11595 4035 11598
rect 5257 11595 5323 11598
rect 6177 11658 6243 11661
rect 10869 11658 10935 11661
rect 6177 11656 10935 11658
rect 6177 11600 6182 11656
rect 6238 11600 10874 11656
rect 10930 11600 10935 11656
rect 6177 11598 10935 11600
rect 6177 11595 6243 11598
rect 10869 11595 10935 11598
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 8109 11250 8175 11253
rect 9857 11250 9923 11253
rect 8109 11248 9923 11250
rect 8109 11192 8114 11248
rect 8170 11192 9862 11248
rect 9918 11192 9923 11248
rect 8109 11190 9923 11192
rect 8109 11187 8175 11190
rect 9857 11187 9923 11190
rect 8753 11114 8819 11117
rect 11605 11114 11671 11117
rect 8753 11112 11671 11114
rect 8753 11056 8758 11112
rect 8814 11056 11610 11112
rect 11666 11056 11671 11112
rect 8753 11054 11671 11056
rect 8753 11051 8819 11054
rect 11605 11051 11671 11054
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 3877 10706 3943 10709
rect 10961 10706 11027 10709
rect 3877 10704 11027 10706
rect 3877 10648 3882 10704
rect 3938 10648 10966 10704
rect 11022 10648 11027 10704
rect 3877 10646 11027 10648
rect 3877 10643 3943 10646
rect 10961 10643 11027 10646
rect 9489 10570 9555 10573
rect 11421 10570 11487 10573
rect 9489 10568 11487 10570
rect 9489 10512 9494 10568
rect 9550 10512 11426 10568
rect 11482 10512 11487 10568
rect 9489 10510 11487 10512
rect 9489 10507 9555 10510
rect 11421 10507 11487 10510
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 3049 10298 3115 10301
rect 4521 10298 4587 10301
rect 3049 10296 4587 10298
rect 3049 10240 3054 10296
rect 3110 10240 4526 10296
rect 4582 10240 4587 10296
rect 3049 10238 4587 10240
rect 3049 10235 3115 10238
rect 4521 10235 4587 10238
rect 9581 10162 9647 10165
rect 11513 10162 11579 10165
rect 9581 10160 11579 10162
rect 9581 10104 9586 10160
rect 9642 10104 11518 10160
rect 11574 10104 11579 10160
rect 9581 10102 11579 10104
rect 9581 10099 9647 10102
rect 11513 10099 11579 10102
rect 9949 10026 10015 10029
rect 7422 10024 10015 10026
rect 7422 9968 9954 10024
rect 10010 9968 10015 10024
rect 7422 9966 10015 9968
rect 4613 9890 4679 9893
rect 7422 9890 7482 9966
rect 9949 9963 10015 9966
rect 4613 9888 7482 9890
rect 4613 9832 4618 9888
rect 4674 9832 7482 9888
rect 4613 9830 7482 9832
rect 4613 9827 4679 9830
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 2405 9618 2471 9621
rect 3233 9618 3299 9621
rect 6545 9618 6611 9621
rect 2405 9616 6611 9618
rect 2405 9560 2410 9616
rect 2466 9560 3238 9616
rect 3294 9560 6550 9616
rect 6606 9560 6611 9616
rect 2405 9558 6611 9560
rect 2405 9555 2471 9558
rect 3233 9555 3299 9558
rect 6545 9555 6611 9558
rect 5073 9482 5139 9485
rect 8385 9482 8451 9485
rect 5073 9480 8451 9482
rect 5073 9424 5078 9480
rect 5134 9424 8390 9480
rect 8446 9424 8451 9480
rect 5073 9422 8451 9424
rect 5073 9419 5139 9422
rect 8385 9419 8451 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 11237 9074 11303 9077
rect 15520 9074 16000 9104
rect 11237 9072 16000 9074
rect 11237 9016 11242 9072
rect 11298 9016 16000 9072
rect 11237 9014 16000 9016
rect 11237 9011 11303 9014
rect 15520 8984 16000 9014
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 381 8258 447 8261
rect 4521 8258 4587 8261
rect 381 8256 4587 8258
rect 381 8200 386 8256
rect 442 8200 4526 8256
rect 4582 8200 4587 8256
rect 381 8198 4587 8200
rect 381 8195 447 8198
rect 4521 8195 4587 8198
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 4429 7986 4495 7989
rect 6177 7986 6243 7989
rect 4429 7984 6243 7986
rect 4429 7928 4434 7984
rect 4490 7928 6182 7984
rect 6238 7928 6243 7984
rect 4429 7926 6243 7928
rect 4429 7923 4495 7926
rect 6177 7923 6243 7926
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 0 7442 480 7472
rect 2773 7442 2839 7445
rect 0 7440 2839 7442
rect 0 7384 2778 7440
rect 2834 7384 2839 7440
rect 0 7382 2839 7384
rect 0 7352 480 7382
rect 2773 7379 2839 7382
rect 9765 7306 9831 7309
rect 11421 7306 11487 7309
rect 6134 7304 11487 7306
rect 6134 7248 9770 7304
rect 9826 7248 11426 7304
rect 11482 7248 11487 7304
rect 6134 7246 11487 7248
rect 3417 7170 3483 7173
rect 6134 7170 6194 7246
rect 9765 7243 9831 7246
rect 11421 7243 11487 7246
rect 3417 7168 6194 7170
rect 3417 7112 3422 7168
rect 3478 7112 6194 7168
rect 3417 7110 6194 7112
rect 3417 7107 3483 7110
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 3141 6898 3207 6901
rect 4705 6898 4771 6901
rect 3141 6896 4771 6898
rect 3141 6840 3146 6896
rect 3202 6840 4710 6896
rect 4766 6840 4771 6896
rect 3141 6838 4771 6840
rect 3141 6835 3207 6838
rect 4705 6835 4771 6838
rect 4981 6898 5047 6901
rect 10225 6898 10291 6901
rect 4981 6896 10291 6898
rect 4981 6840 4986 6896
rect 5042 6840 10230 6896
rect 10286 6840 10291 6896
rect 4981 6838 10291 6840
rect 4981 6835 5047 6838
rect 10225 6835 10291 6838
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 5441 6354 5507 6357
rect 7465 6354 7531 6357
rect 5441 6352 7531 6354
rect 5441 6296 5446 6352
rect 5502 6296 7470 6352
rect 7526 6296 7531 6352
rect 5441 6294 7531 6296
rect 5441 6291 5507 6294
rect 7465 6291 7531 6294
rect 2497 6218 2563 6221
rect 7005 6218 7071 6221
rect 9673 6218 9739 6221
rect 2497 6216 9739 6218
rect 2497 6160 2502 6216
rect 2558 6160 7010 6216
rect 7066 6160 9678 6216
rect 9734 6160 9739 6216
rect 2497 6158 9739 6160
rect 2497 6155 2563 6158
rect 7005 6155 7071 6158
rect 9673 6155 9739 6158
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 7097 5810 7163 5813
rect 9673 5810 9739 5813
rect 7097 5808 9739 5810
rect 7097 5752 7102 5808
rect 7158 5752 9678 5808
rect 9734 5752 9739 5808
rect 7097 5750 9739 5752
rect 7097 5747 7163 5750
rect 9673 5747 9739 5750
rect 4797 5674 4863 5677
rect 7097 5674 7163 5677
rect 4797 5672 7163 5674
rect 4797 5616 4802 5672
rect 4858 5616 7102 5672
rect 7158 5616 7163 5672
rect 4797 5614 7163 5616
rect 4797 5611 4863 5614
rect 7097 5611 7163 5614
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 15520 5402 16000 5432
rect 14782 5342 16000 5402
rect 12341 5266 12407 5269
rect 14782 5266 14842 5342
rect 15520 5312 16000 5342
rect 12341 5264 14842 5266
rect 12341 5208 12346 5264
rect 12402 5208 14842 5264
rect 12341 5206 14842 5208
rect 12341 5203 12407 5206
rect 2865 5130 2931 5133
rect 6821 5130 6887 5133
rect 2865 5128 6887 5130
rect 2865 5072 2870 5128
rect 2926 5072 6826 5128
rect 6882 5072 6887 5128
rect 2865 5070 6887 5072
rect 2865 5067 2931 5070
rect 6821 5067 6887 5070
rect 2405 4994 2471 4997
rect 5257 4994 5323 4997
rect 2405 4992 5323 4994
rect 2405 4936 2410 4992
rect 2466 4936 5262 4992
rect 5318 4936 5323 4992
rect 2405 4934 5323 4936
rect 2405 4931 2471 4934
rect 5257 4931 5323 4934
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 3233 4722 3299 4725
rect 7925 4722 7991 4725
rect 10685 4722 10751 4725
rect 3233 4720 10751 4722
rect 3233 4664 3238 4720
rect 3294 4664 7930 4720
rect 7986 4664 10690 4720
rect 10746 4664 10751 4720
rect 3233 4662 10751 4664
rect 3233 4659 3299 4662
rect 7925 4659 7991 4662
rect 10685 4659 10751 4662
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 9673 4314 9739 4317
rect 13169 4314 13235 4317
rect 9673 4312 13235 4314
rect 9673 4256 9678 4312
rect 9734 4256 13174 4312
rect 13230 4256 13235 4312
rect 9673 4254 13235 4256
rect 9673 4251 9739 4254
rect 13169 4251 13235 4254
rect 3785 4178 3851 4181
rect 5625 4178 5691 4181
rect 3785 4176 5691 4178
rect 3785 4120 3790 4176
rect 3846 4120 5630 4176
rect 5686 4120 5691 4176
rect 3785 4118 5691 4120
rect 3785 4115 3851 4118
rect 5625 4115 5691 4118
rect 7005 4178 7071 4181
rect 13721 4178 13787 4181
rect 7005 4176 13787 4178
rect 7005 4120 7010 4176
rect 7066 4120 13726 4176
rect 13782 4120 13787 4176
rect 7005 4118 13787 4120
rect 7005 4115 7071 4118
rect 13721 4115 13787 4118
rect 3693 4042 3759 4045
rect 5901 4042 5967 4045
rect 7281 4042 7347 4045
rect 3693 4040 5967 4042
rect 3693 3984 3698 4040
rect 3754 3984 5906 4040
rect 5962 3984 5967 4040
rect 3693 3982 5967 3984
rect 3693 3979 3759 3982
rect 5901 3979 5967 3982
rect 6134 4040 7347 4042
rect 6134 3984 7286 4040
rect 7342 3984 7347 4040
rect 6134 3982 7347 3984
rect 6134 3909 6194 3982
rect 7281 3979 7347 3982
rect 3325 3906 3391 3909
rect 6085 3906 6194 3909
rect 3325 3904 6194 3906
rect 3325 3848 3330 3904
rect 3386 3848 6090 3904
rect 6146 3848 6194 3904
rect 3325 3846 6194 3848
rect 3325 3843 3391 3846
rect 6085 3843 6151 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 2129 3770 2195 3773
rect 2957 3770 3023 3773
rect 4337 3770 4403 3773
rect 2129 3768 4403 3770
rect 2129 3712 2134 3768
rect 2190 3712 2962 3768
rect 3018 3712 4342 3768
rect 4398 3712 4403 3768
rect 2129 3710 4403 3712
rect 2129 3707 2195 3710
rect 2957 3707 3023 3710
rect 4337 3707 4403 3710
rect 2313 3634 2379 3637
rect 3233 3634 3299 3637
rect 2313 3632 3299 3634
rect 2313 3576 2318 3632
rect 2374 3576 3238 3632
rect 3294 3576 3299 3632
rect 2313 3574 3299 3576
rect 2313 3571 2379 3574
rect 3233 3571 3299 3574
rect 3417 3634 3483 3637
rect 9857 3634 9923 3637
rect 3417 3632 9923 3634
rect 3417 3576 3422 3632
rect 3478 3576 9862 3632
rect 9918 3576 9923 3632
rect 3417 3574 9923 3576
rect 3417 3571 3483 3574
rect 9857 3571 9923 3574
rect 2497 3498 2563 3501
rect 5901 3498 5967 3501
rect 2497 3496 5967 3498
rect 2497 3440 2502 3496
rect 2558 3440 5906 3496
rect 5962 3440 5967 3496
rect 2497 3438 5967 3440
rect 2497 3435 2563 3438
rect 5901 3435 5967 3438
rect 6637 3498 6703 3501
rect 9673 3498 9739 3501
rect 6637 3496 9739 3498
rect 6637 3440 6642 3496
rect 6698 3440 9678 3496
rect 9734 3440 9739 3496
rect 6637 3438 9739 3440
rect 6637 3435 6703 3438
rect 9673 3435 9739 3438
rect 5717 3362 5783 3365
rect 7465 3362 7531 3365
rect 5717 3360 7531 3362
rect 5717 3304 5722 3360
rect 5778 3304 7470 3360
rect 7526 3304 7531 3360
rect 5717 3302 7531 3304
rect 5717 3299 5783 3302
rect 7465 3299 7531 3302
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 5165 3226 5231 3229
rect 5165 3224 7160 3226
rect 5165 3168 5170 3224
rect 5226 3168 7160 3224
rect 5165 3166 7160 3168
rect 5165 3163 5231 3166
rect 3049 3090 3115 3093
rect 6821 3090 6887 3093
rect 3049 3088 6887 3090
rect 3049 3032 3054 3088
rect 3110 3032 6826 3088
rect 6882 3032 6887 3088
rect 3049 3030 6887 3032
rect 7100 3090 7160 3166
rect 10777 3090 10843 3093
rect 7100 3088 10843 3090
rect 7100 3032 10782 3088
rect 10838 3032 10843 3088
rect 7100 3030 10843 3032
rect 3049 3027 3115 3030
rect 6821 3027 6887 3030
rect 10777 3027 10843 3030
rect 3233 2954 3299 2957
rect 6637 2954 6703 2957
rect 3233 2952 6703 2954
rect 3233 2896 3238 2952
rect 3294 2896 6642 2952
rect 6698 2896 6703 2952
rect 3233 2894 6703 2896
rect 3233 2891 3299 2894
rect 6637 2891 6703 2894
rect 7005 2954 7071 2957
rect 12801 2954 12867 2957
rect 7005 2952 12867 2954
rect 7005 2896 7010 2952
rect 7066 2896 12806 2952
rect 12862 2896 12867 2952
rect 7005 2894 12867 2896
rect 7005 2891 7071 2894
rect 12801 2891 12867 2894
rect 6729 2818 6795 2821
rect 11329 2818 11395 2821
rect 6729 2816 11395 2818
rect 6729 2760 6734 2816
rect 6790 2760 11334 2816
rect 11390 2760 11395 2816
rect 6729 2758 11395 2760
rect 6729 2755 6795 2758
rect 11329 2755 11395 2758
rect 12341 2818 12407 2821
rect 15469 2818 15535 2821
rect 12341 2816 15535 2818
rect 12341 2760 12346 2816
rect 12402 2760 15474 2816
rect 15530 2760 15535 2816
rect 12341 2758 15535 2760
rect 12341 2755 12407 2758
rect 15469 2755 15535 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 2313 2682 2379 2685
rect 4981 2682 5047 2685
rect 2313 2680 5047 2682
rect 2313 2624 2318 2680
rect 2374 2624 4986 2680
rect 5042 2624 5047 2680
rect 2313 2622 5047 2624
rect 2313 2619 2379 2622
rect 4981 2619 5047 2622
rect 7005 2682 7071 2685
rect 10317 2682 10383 2685
rect 7005 2680 10383 2682
rect 7005 2624 7010 2680
rect 7066 2624 10322 2680
rect 10378 2624 10383 2680
rect 7005 2622 10383 2624
rect 7005 2619 7071 2622
rect 10317 2619 10383 2622
rect 0 2546 480 2576
rect 1393 2546 1459 2549
rect 0 2544 1459 2546
rect 0 2488 1398 2544
rect 1454 2488 1459 2544
rect 0 2486 1459 2488
rect 0 2456 480 2486
rect 1393 2483 1459 2486
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 13813 1866 13879 1869
rect 15520 1866 16000 1896
rect 13813 1864 16000 1866
rect 13813 1808 13818 1864
rect 13874 1808 16000 1864
rect 13813 1806 16000 1808
rect 13813 1803 13879 1806
rect 15520 1776 16000 1806
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 10364 28928 10428 28932
rect 10364 28872 10414 28928
rect 10414 28872 10428 28928
rect 10364 28868 10428 28872
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 6132 27296 6196 27300
rect 6132 27240 6146 27296
rect 6146 27240 6196 27296
rect 6132 27236 6196 27240
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 10364 19680 10428 19684
rect 10364 19624 10378 19680
rect 10378 19624 10428 19680
rect 10364 19620 10428 19624
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6132 19212 6196 19276
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 7052 17444 7116 17508
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 7052 11792 7116 11796
rect 7052 11736 7066 11792
rect 7066 11736 7116 11792
rect 7052 11732 7116 11736
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6131 27300 6197 27301
rect 6131 27236 6132 27300
rect 6196 27236 6197 27300
rect 6131 27235 6197 27236
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 6134 19277 6194 27235
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6131 19276 6197 19277
rect 6131 19212 6132 19276
rect 6196 19212 6197 19276
rect 6131 19211 6197 19212
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 10363 28932 10429 28933
rect 10363 28868 10364 28932
rect 10428 28868 10429 28932
rect 10363 28867 10429 28868
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 10366 19685 10426 28867
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 10363 19684 10429 19685
rect 10363 19620 10364 19684
rect 10428 19620 10429 19684
rect 10363 19619 10429 19620
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 7051 17508 7117 17509
rect 7051 17444 7052 17508
rect 7116 17444 7117 17508
rect 7051 17443 7117 17444
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 7054 11797 7114 17443
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 7051 11796 7117 11797
rect 7051 11732 7052 11796
rect 7116 11732 7117 11796
rect 7051 11731 7117 11732
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_8
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_12
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_50
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_44
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _183_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_77
timestamp 1586364061
transform 1 0 8188 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_70
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_89
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_94 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_92 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_104
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_108
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _180_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_123 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _181_
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_135
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_135 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_139
timestamp 1586364061
transform 1 0 13892 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 406 592
use scs8hd_conb_1  _172_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_29
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_43
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_108
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_120
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_132
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_8
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_41
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_76
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_58
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_82
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_86
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_8  FILLER_4_96
timestamp 1586364061
transform 1 0 9936 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_nor2_4  _074_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _182_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_17
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 774 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_47
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_75
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_79
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_90
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_96
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_108
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_97
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_11
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _069_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_37
timestamp 1586364061
transform 1 0 4508 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_60
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_21
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_29
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_114
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_126
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_102
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_43
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_47
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _083_
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_37
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_conb_1  _173_
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_82
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_71
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_24
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_28
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_84
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_120
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_28
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_119
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_131
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_103
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_38
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_54
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_73
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_35
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_39
timestamp 1586364061
transform 1 0 4692 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_54
timestamp 1586364061
transform 1 0 6072 0 -1 13600
box -38 -48 774 592
use scs8hd_conb_1  _174_
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_65
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_69
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_73
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_8  _146_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_127
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_58
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_82
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_87
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_104
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_11
timestamp 1586364061
transform 1 0 2116 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_16
timestamp 1586364061
transform 1 0 2576 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_28
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_59
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_63
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_78
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_115
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_127
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_139
timestamp 1586364061
transform 1 0 13892 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_46
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_88
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 314 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _175_
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_or3_4  _082_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_123
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_23
timestamp 1586364061
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_30
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_49
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_25_55
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_nor3_4  _144_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__144__C
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 406 592
use scs8hd_conb_1  _171_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_137
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 590 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 4232 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_43
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 866 592
use scs8hd_or3_4  _110_
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_or3_4  _118_
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 866 592
use scs8hd_nor3_4  _143_
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use scs8hd_or3_4  _068_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_95
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 866 592
use scs8hd_inv_8  _152_
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use scs8hd_decap_4  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 13156 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_129
timestamp 1586364061
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_133
timestamp 1586364061
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_145
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_16
timestamp 1586364061
transform 1 0 2576 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_35
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_39
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_119
timestamp 1586364061
transform 1 0 12052 0 -1 17952
box -38 -48 774 592
use scs8hd_or3_4  _153_
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_136
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 590 592
use scs8hd_decap_3  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 866 592
use scs8hd_buf_1  _119_
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_17
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_81
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_or4_4  _135_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_85
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _067_
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_102
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_109
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_113
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_117
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_130
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_142
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_4  FILLER_30_12
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_16
timestamp 1586364061
transform 1 0 2576 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_40
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_59
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_76
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 406 592
use scs8hd_or3_4  _066_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_87
timestamp 1586364061
transform 1 0 9108 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_119
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_131
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_143
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_26
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_30
timestamp 1586364061
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_45
timestamp 1586364061
transform 1 0 5244 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_50
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_54
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_58
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 130 592
use scs8hd_or2_4  _100_
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _126_
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_90
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_103
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_107
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_111
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_115
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_conb_1  _176_
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_37
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_41
timestamp 1586364061
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_45
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_76
timestamp 1586364061
transform 1 0 8096 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 774 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_115
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_127
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 4140 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_48
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_54
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_42
timestamp 1586364061
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_54
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_58
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_72
timestamp 1586364061
transform 1 0 7728 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_75
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_83
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_79
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _148_
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 866 592
use scs8hd_or3_4  _154_
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 866 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__C
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_88
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_92
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_89
timestamp 1586364061
transform 1 0 9292 0 -1 21216
box -38 -48 130 592
use scs8hd_or3_4  _167_
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_105
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_109
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_106
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_116
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_123
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_135
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_143
timestamp 1586364061
transform 1 0 14260 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_30
timestamp 1586364061
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_43
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_or3_4  _157_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_or3_4  _062_
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_or3_4  _149_
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_105
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _150_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_113
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_126
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_130
timestamp 1586364061
transform 1 0 13064 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_142
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4508 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_48
timestamp 1586364061
transform 1 0 5520 0 -1 22304
box -38 -48 774 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_65
timestamp 1586364061
transform 1 0 7084 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_69
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_8  _147_
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_73
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 9844 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 22304
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 774 592
use scs8hd_or3_4  _164_
timestamp 1586364061
transform 1 0 11776 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_buf_1  _073_
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_22
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4600 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_30
timestamp 1586364061
transform 1 0 3864 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_34
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_49
timestamp 1586364061
transform 1 0 5612 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 8096 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_78
timestamp 1586364061
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use scs8hd_or3_4  _161_
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_88
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_105
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_117
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_buf_1  _063_
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_137
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_141
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_145
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 2944 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 4232 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_29
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_36
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_49
timestamp 1586364061
transform 1 0 5612 0 -1 23392
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 23392
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_1  _151_
timestamp 1586364061
transform 1 0 8096 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_72
timestamp 1586364061
transform 1 0 7728 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_79
timestamp 1586364061
transform 1 0 8372 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_83
timestamp 1586364061
transform 1 0 8740 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 8924 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_87
timestamp 1586364061
transform 1 0 9108 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_91
timestamp 1586364061
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_96
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_100
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 774 592
use scs8hd_conb_1  _170_
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_128
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_19
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 2944 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 2576 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 866 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_36
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_29
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_41
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 5980 0 -1 24480
box -38 -48 314 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_46
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_50
timestamp 1586364061
transform 1 0 5704 0 -1 24480
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_60
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_1  _168_
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_73
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_77
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_73
timestamp 1586364061
transform 1 0 7820 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_88
timestamp 1586364061
transform 1 0 9200 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_90
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_96
timestamp 1586364061
transform 1 0 9936 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_94
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _162_
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 10120 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_107
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_100
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_104
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_121
timestamp 1586364061
transform 1 0 12236 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_39_139
timestamp 1586364061
transform 1 0 13892 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_145
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_41_11
timestamp 1586364061
transform 1 0 2116 0 1 24480
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 2392 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 2760 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_16
timestamp 1586364061
transform 1 0 2576 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_20
timestamp 1586364061
transform 1 0 2944 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_24
timestamp 1586364061
transform 1 0 3312 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4876 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_36
timestamp 1586364061
transform 1 0 4416 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 130 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_43
timestamp 1586364061
transform 1 0 5060 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_78
timestamp 1586364061
transform 1 0 8280 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_92
timestamp 1586364061
transform 1 0 9568 0 1 24480
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_113
timestamp 1586364061
transform 1 0 11500 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_137
timestamp 1586364061
transform 1 0 13708 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_41_145
timestamp 1586364061
transform 1 0 14444 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_11
timestamp 1586364061
transform 1 0 2116 0 -1 25568
box -38 -48 314 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 2392 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_8  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4232 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_36
timestamp 1586364061
transform 1 0 4416 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_52
timestamp 1586364061
transform 1 0 5888 0 -1 25568
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_58
timestamp 1586364061
transform 1 0 6440 0 -1 25568
box -38 -48 130 592
use scs8hd_conb_1  _177_
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_72
timestamp 1586364061
transform 1 0 7728 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_76
timestamp 1586364061
transform 1 0 8096 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_83
timestamp 1586364061
transform 1 0 8740 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_91
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 25568
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_42_108
timestamp 1586364061
transform 1 0 11040 0 -1 25568
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 25568
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_127
timestamp 1586364061
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_131
timestamp 1586364061
transform 1 0 13156 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_8  FILLER_42_138
timestamp 1586364061
transform 1 0 13800 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4232 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_30
timestamp 1586364061
transform 1 0 3864 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6072 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_45
timestamp 1586364061
transform 1 0 5244 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_49
timestamp 1586364061
transform 1 0 5612 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_53
timestamp 1586364061
transform 1 0 5980 0 1 25568
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 7360 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_56
timestamp 1586364061
transform 1 0 6256 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_60
timestamp 1586364061
transform 1 0 6624 0 1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_43_65
timestamp 1586364061
transform 1 0 7084 0 1 25568
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8280 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 7728 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_70
timestamp 1586364061
transform 1 0 7544 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_89
timestamp 1586364061
transform 1 0 9292 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_93
timestamp 1586364061
transform 1 0 9660 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10028 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_108
timestamp 1586364061
transform 1 0 11040 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_112
timestamp 1586364061
transform 1 0 11408 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_116
timestamp 1586364061
transform 1 0 11776 0 1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 13432 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_132
timestamp 1586364061
transform 1 0 13248 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_136
timestamp 1586364061
transform 1 0 13616 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_144
timestamp 1586364061
transform 1 0 14352 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4324 0 -1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_46
timestamp 1586364061
transform 1 0 5336 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_50
timestamp 1586364061
transform 1 0 5704 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_63
timestamp 1586364061
transform 1 0 6900 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_67
timestamp 1586364061
transform 1 0 7268 0 -1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 7820 0 -1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_44_71
timestamp 1586364061
transform 1 0 7636 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_82
timestamp 1586364061
transform 1 0 8648 0 -1 26656
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_88
timestamp 1586364061
transform 1 0 9200 0 -1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_102
timestamp 1586364061
transform 1 0 10488 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_106
timestamp 1586364061
transform 1 0 10856 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_119
timestamp 1586364061
transform 1 0 12052 0 -1 26656
box -38 -48 406 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 12788 0 -1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_44_125
timestamp 1586364061
transform 1 0 12604 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_136
timestamp 1586364061
transform 1 0 13616 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_144
timestamp 1586364061
transform 1 0 14352 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3036 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3496 0 1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 590 592
use scs8hd_fill_2  FILLER_45_24
timestamp 1586364061
transform 1 0 3312 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_28
timestamp 1586364061
transform 1 0 3680 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_35
timestamp 1586364061
transform 1 0 4324 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_52
timestamp 1586364061
transform 1 0 5888 0 1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_57
timestamp 1586364061
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_71
timestamp 1586364061
transform 1 0 7636 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_75
timestamp 1586364061
transform 1 0 8004 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_82
timestamp 1586364061
transform 1 0 8648 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_86
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_90
timestamp 1586364061
transform 1 0 9384 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_101
timestamp 1586364061
transform 1 0 10396 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_105
timestamp 1586364061
transform 1 0 10764 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_112
timestamp 1586364061
transform 1 0 11408 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_116
timestamp 1586364061
transform 1 0 11776 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_120
timestamp 1586364061
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_126
timestamp 1586364061
transform 1 0 12696 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_130
timestamp 1586364061
transform 1 0 13064 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_137
timestamp 1586364061
transform 1 0 13708 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_141
timestamp 1586364061
transform 1 0 14076 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_145
timestamp 1586364061
transform 1 0 14444 0 1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3956 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_34
timestamp 1586364061
transform 1 0 4232 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_38
timestamp 1586364061
transform 1 0 4600 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_37
timestamp 1586364061
transform 1 0 4508 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_41
timestamp 1586364061
transform 1 0 4876 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 6072 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_54
timestamp 1586364061
transform 1 0 6072 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_58
timestamp 1586364061
transform 1 0 6440 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_56
timestamp 1586364061
transform 1 0 6256 0 1 27744
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 8740 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_71
timestamp 1586364061
transform 1 0 7636 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_6  FILLER_46_82
timestamp 1586364061
transform 1 0 8648 0 -1 27744
box -38 -48 590 592
use scs8hd_fill_2  FILLER_47_73
timestamp 1586364061
transform 1 0 7820 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_77
timestamp 1586364061
transform 1 0 8188 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_81
timestamp 1586364061
transform 1 0 8556 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 9292 0 1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 9108 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 9292 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_88
timestamp 1586364061
transform 1 0 9200 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_1  FILLER_46_91
timestamp 1586364061
transform 1 0 9476 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_85
timestamp 1586364061
transform 1 0 8924 0 1 27744
box -38 -48 222 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 10856 0 1 27744
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 10304 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_102
timestamp 1586364061
transform 1 0 10488 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_98
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_47_102
timestamp 1586364061
transform 1 0 10488 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_109
timestamp 1586364061
transform 1 0 11132 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 11316 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 11684 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_119
timestamp 1586364061
transform 1 0 12052 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_113
timestamp 1586364061
transform 1 0 11500 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_47_117
timestamp 1586364061
transform 1 0 11868 0 1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_47_121
timestamp 1586364061
transform 1 0 12236 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_130
timestamp 1586364061
transform 1 0 13064 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_decap_4  FILLER_46_142
timestamp 1586364061
transform 1 0 14168 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_3  FILLER_47_143
timestamp 1586364061
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 774 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 6072 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_43
timestamp 1586364061
transform 1 0 5060 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_47
timestamp 1586364061
transform 1 0 5428 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_51
timestamp 1586364061
transform 1 0 5796 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 7084 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_63
timestamp 1586364061
transform 1 0 6900 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_67
timestamp 1586364061
transform 1 0 7268 0 -1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 28832
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_48_82
timestamp 1586364061
transform 1 0 8648 0 -1 28832
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 8832 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_48_86
timestamp 1586364061
transform 1 0 9016 0 -1 28832
box -38 -48 590 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 11224 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_48_102
timestamp 1586364061
transform 1 0 10488 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_12  FILLER_48_113
timestamp 1586364061
transform 1 0 11500 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_125
timestamp 1586364061
transform 1 0 12604 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_48_137
timestamp 1586364061
transform 1 0 13708 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_48_145
timestamp 1586364061
transform 1 0 14444 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_53
timestamp 1586364061
transform 1 0 5980 0 1 28832
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7360 0 1 28832
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 6440 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_57
timestamp 1586364061
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use scs8hd_fill_1  FILLER_49_60
timestamp 1586364061
transform 1 0 6624 0 1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 8556 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_79
timestamp 1586364061
transform 1 0 8372 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_83
timestamp 1586364061
transform 1 0 8740 0 1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9108 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 28832
box -38 -48 222 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 10856 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_98
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_102
timestamp 1586364061
transform 1 0 10488 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_109
timestamp 1586364061
transform 1 0 11132 0 1 28832
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_115
timestamp 1586364061
transform 1 0 11684 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_118
timestamp 1586364061
transform 1 0 11960 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_143
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_50_46
timestamp 1586364061
transform 1 0 5336 0 -1 29920
box -38 -48 1142 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 6440 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 7452 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_67
timestamp 1586364061
transform 1 0 7268 0 -1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 8004 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_71
timestamp 1586364061
transform 1 0 7636 0 -1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_50_84
timestamp 1586364061
transform 1 0 8832 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_50_89
timestamp 1586364061
transform 1 0 9292 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 29920
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_50_108
timestamp 1586364061
transform 1 0 11040 0 -1 29920
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 29920
box -38 -48 866 592
use scs8hd_decap_12  FILLER_50_125
timestamp 1586364061
transform 1 0 12604 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_137
timestamp 1586364061
transform 1 0 13708 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_50_145
timestamp 1586364061
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 7268 0 1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 7084 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_76
timestamp 1586364061
transform 1 0 8096 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_80
timestamp 1586364061
transform 1 0 8464 0 1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9844 0 1 29920
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8832 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_87
timestamp 1586364061
transform 1 0 9108 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_91
timestamp 1586364061
transform 1 0 9476 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_106
timestamp 1586364061
transform 1 0 10856 0 1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_112
timestamp 1586364061
transform 1 0 11408 0 1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_51_116
timestamp 1586364061
transform 1 0 11776 0 1 29920
box -38 -48 590 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6072 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 5704 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_53_47
timestamp 1586364061
transform 1 0 5428 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_52
timestamp 1586364061
transform 1 0 5888 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 866 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 6992 0 -1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6808 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 590 592
use scs8hd_decap_4  FILLER_52_67
timestamp 1586364061
transform 1 0 7268 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_53_56
timestamp 1586364061
transform 1 0 6256 0 1 31008
box -38 -48 314 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 8648 0 1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 8464 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 7820 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7636 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_73
timestamp 1586364061
transform 1 0 7820 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_71
timestamp 1586364061
transform 1 0 7636 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_75
timestamp 1586364061
transform 1 0 8004 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_79
timestamp 1586364061
transform 1 0 8372 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 9660 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_84
timestamp 1586364061
transform 1 0 8832 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_2  FILLER_53_91
timestamp 1586364061
transform 1 0 9476 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_95
timestamp 1586364061
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 10028 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_102
timestamp 1586364061
transform 1 0 10488 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_106
timestamp 1586364061
transform 1 0 10856 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_99
timestamp 1586364061
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_119
timestamp 1586364061
transform 1 0 12052 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_112
timestamp 1586364061
transform 1 0 11408 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_53_116
timestamp 1586364061
transform 1 0 11776 0 1 31008
box -38 -48 590 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_131
timestamp 1586364061
transform 1 0 13156 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_52_143
timestamp 1586364061
transform 1 0 14260 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_53_143
timestamp 1586364061
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 6072 0 -1 32096
box -38 -48 866 592
use scs8hd_decap_8  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_54_52
timestamp 1586364061
transform 1 0 5888 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_63
timestamp 1586364061
transform 1 0 6900 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_67
timestamp 1586364061
transform 1 0 7268 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 7636 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 8648 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_84
timestamp 1586364061
transform 1 0 8832 0 -1 32096
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_102
timestamp 1586364061
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_106
timestamp 1586364061
transform 1 0 10856 0 -1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_113
timestamp 1586364061
transform 1 0 11500 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_54_117
timestamp 1586364061
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_129
timestamp 1586364061
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_4  FILLER_54_141
timestamp 1586364061
transform 1 0 14076 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_47
timestamp 1586364061
transform 1 0 5428 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_52
timestamp 1586364061
transform 1 0 5888 0 1 32096
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_57
timestamp 1586364061
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8556 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_73
timestamp 1586364061
transform 1 0 7820 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_77
timestamp 1586364061
transform 1 0 8188 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_92
timestamp 1586364061
transform 1 0 9568 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_96
timestamp 1586364061
transform 1 0 9936 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 10304 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 10120 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_109
timestamp 1586364061
transform 1 0 11132 0 1 32096
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_113
timestamp 1586364061
transform 1 0 11500 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_117
timestamp 1586364061
transform 1 0 11868 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_126
timestamp 1586364061
transform 1 0 12696 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_131
timestamp 1586364061
transform 1 0 13156 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_143
timestamp 1586364061
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 590 592
use scs8hd_fill_2  FILLER_56_53
timestamp 1586364061
transform 1 0 5980 0 -1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 33184
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_56_57
timestamp 1586364061
transform 1 0 6348 0 -1 33184
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_72
timestamp 1586364061
transform 1 0 7728 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_76
timestamp 1586364061
transform 1 0 8096 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_83
timestamp 1586364061
transform 1 0 8740 0 -1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_87
timestamp 1586364061
transform 1 0 9108 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_91
timestamp 1586364061
transform 1 0 9476 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_104
timestamp 1586364061
transform 1 0 10672 0 -1 33184
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_121
timestamp 1586364061
transform 1 0 12236 0 -1 33184
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_4  FILLER_56_125
timestamp 1586364061
transform 1 0 12604 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_132
timestamp 1586364061
transform 1 0 13248 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_56_144
timestamp 1586364061
transform 1 0 14352 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_42
timestamp 1586364061
transform 1 0 4968 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_46
timestamp 1586364061
transform 1 0 5336 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_53
timestamp 1586364061
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_57
timestamp 1586364061
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_57_66
timestamp 1586364061
transform 1 0 7176 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_78
timestamp 1586364061
transform 1 0 8280 0 1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_57_82
timestamp 1586364061
transform 1 0 8648 0 1 33184
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9292 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_85
timestamp 1586364061
transform 1 0 8924 0 1 33184
box -38 -48 222 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 11040 0 1 33184
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_100
timestamp 1586364061
transform 1 0 10304 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_104
timestamp 1586364061
transform 1 0 10672 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 11592 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_112
timestamp 1586364061
transform 1 0 11408 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_116
timestamp 1586364061
transform 1 0 11776 0 1 33184
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 13432 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_132
timestamp 1586364061
transform 1 0 13248 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_136
timestamp 1586364061
transform 1 0 13616 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_144
timestamp 1586364061
transform 1 0 14352 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 34272
box -38 -48 866 592
use scs8hd_decap_8  FILLER_58_47
timestamp 1586364061
transform 1 0 5428 0 -1 34272
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_64
timestamp 1586364061
transform 1 0 6992 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 34272
box -38 -48 866 592
use scs8hd_fill_1  FILLER_58_71
timestamp 1586364061
transform 1 0 7636 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_58_81
timestamp 1586364061
transform 1 0 8556 0 -1 34272
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  FILLER_58_89
timestamp 1586364061
transform 1 0 9292 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_104
timestamp 1586364061
transform 1 0 10672 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_108
timestamp 1586364061
transform 1 0 11040 0 -1 34272
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 34272
box -38 -48 866 592
use scs8hd_decap_8  FILLER_58_121
timestamp 1586364061
transform 1 0 12236 0 -1 34272
box -38 -48 774 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 12972 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_133
timestamp 1586364061
transform 1 0 13340 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 5612 0 1 34272
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 6164 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_47
timestamp 1586364061
transform 1 0 5428 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_53
timestamp 1586364061
transform 1 0 5980 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_8  FILLER_60_55
timestamp 1586364061
transform 1 0 6164 0 -1 35360
box -38 -48 774 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 6900 0 -1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 6992 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_57
timestamp 1586364061
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_66
timestamp 1586364061
transform 1 0 7176 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_60_67
timestamp 1586364061
transform 1 0 7268 0 -1 35360
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 34272
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_79
timestamp 1586364061
transform 1 0 8372 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_83
timestamp 1586364061
transform 1 0 8740 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_60_72
timestamp 1586364061
transform 1 0 7728 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_4  FILLER_60_88
timestamp 1586364061
transform 1 0 9200 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_84
timestamp 1586364061
transform 1 0 8832 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 34272
box -38 -48 222 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 9108 0 1 34272
box -38 -48 406 592
use scs8hd_decap_6  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_95
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_91
timestamp 1586364061
transform 1 0 9476 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 34272
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_108
timestamp 1586364061
transform 1 0 11040 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_110
timestamp 1586364061
transform 1 0 11224 0 -1 35360
box -38 -48 774 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 35360
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_59_112
timestamp 1586364061
transform 1 0 11408 0 1 34272
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_120
timestamp 1586364061
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_121
timestamp 1586364061
transform 1 0 12236 0 -1 35360
box -38 -48 774 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 12972 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 13340 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_127
timestamp 1586364061
transform 1 0 12788 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_131
timestamp 1586364061
transform 1 0 13156 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_59_135
timestamp 1586364061
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_133
timestamp 1586364061
transform 1 0 13340 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_59_143
timestamp 1586364061
transform 1 0 14260 0 1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 7360 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_66
timestamp 1586364061
transform 1 0 7176 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_70
timestamp 1586364061
transform 1 0 7544 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 9200 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_90
timestamp 1586364061
transform 1 0 9384 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_95
timestamp 1586364061
transform 1 0 9844 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_108
timestamp 1586364061
transform 1 0 11040 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_120
timestamp 1586364061
transform 1 0 12144 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7452 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 130 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_72
timestamp 1586364061
transform 1 0 7728 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_76
timestamp 1586364061
transform 1 0 8096 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_1  FILLER_62_79
timestamp 1586364061
transform 1 0 8372 0 -1 36448
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_84
timestamp 1586364061
transform 1 0 8832 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  FILLER_62_96
timestamp 1586364061
transform 1 0 9936 0 -1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_62_101
timestamp 1586364061
transform 1 0 10396 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_113
timestamp 1586364061
transform 1 0 11500 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_125
timestamp 1586364061
transform 1 0 12604 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_62_137
timestamp 1586364061
transform 1 0 13708 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 36448
box -38 -48 314 592
use scs8hd_decap_6  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 590 592
use scs8hd_fill_2  FILLER_63_95
timestamp 1586364061
transform 1 0 9844 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_99
timestamp 1586364061
transform 1 0 10212 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_63_111
timestamp 1586364061
transform 1 0 11316 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  FILLER_63_119
timestamp 1586364061
transform 1 0 12052 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal3 s 15520 5312 16000 5432 6 address[0]
port 0 nsew default input
rlabel metal3 s 15520 8984 16000 9104 6 address[1]
port 1 nsew default input
rlabel metal3 s 15520 12656 16000 12776 6 address[2]
port 2 nsew default input
rlabel metal3 s 15520 16192 16000 16312 6 address[3]
port 3 nsew default input
rlabel metal3 s 15520 19864 16000 19984 6 address[4]
port 4 nsew default input
rlabel metal3 s 15520 23536 16000 23656 6 address[5]
port 5 nsew default input
rlabel metal3 s 15520 27208 16000 27328 6 address[6]
port 6 nsew default input
rlabel metal2 s 386 0 442 480 6 chany_bottom_in[0]
port 7 nsew default input
rlabel metal2 s 1214 0 1270 480 6 chany_bottom_in[1]
port 8 nsew default input
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_in[2]
port 9 nsew default input
rlabel metal2 s 3054 0 3110 480 6 chany_bottom_in[3]
port 10 nsew default input
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[4]
port 11 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[5]
port 12 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[6]
port 13 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[7]
port 14 nsew default input
rlabel metal2 s 7470 0 7526 480 6 chany_bottom_in[8]
port 15 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_out[0]
port 16 nsew default tristate
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_out[1]
port 17 nsew default tristate
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_out[2]
port 18 nsew default tristate
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_out[3]
port 19 nsew default tristate
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_out[4]
port 20 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_out[5]
port 21 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[6]
port 22 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[7]
port 23 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[8]
port 24 nsew default tristate
rlabel metal2 s 386 39520 442 40000 6 chany_top_in[0]
port 25 nsew default input
rlabel metal2 s 1214 39520 1270 40000 6 chany_top_in[1]
port 26 nsew default input
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_in[2]
port 27 nsew default input
rlabel metal2 s 3054 39520 3110 40000 6 chany_top_in[3]
port 28 nsew default input
rlabel metal2 s 3882 39520 3938 40000 6 chany_top_in[4]
port 29 nsew default input
rlabel metal2 s 4802 39520 4858 40000 6 chany_top_in[5]
port 30 nsew default input
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_in[6]
port 31 nsew default input
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_in[7]
port 32 nsew default input
rlabel metal2 s 7470 39520 7526 40000 6 chany_top_in[8]
port 33 nsew default input
rlabel metal2 s 8390 39520 8446 40000 6 chany_top_out[0]
port 34 nsew default tristate
rlabel metal2 s 9218 39520 9274 40000 6 chany_top_out[1]
port 35 nsew default tristate
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_out[2]
port 36 nsew default tristate
rlabel metal2 s 11058 39520 11114 40000 6 chany_top_out[3]
port 37 nsew default tristate
rlabel metal2 s 11886 39520 11942 40000 6 chany_top_out[4]
port 38 nsew default tristate
rlabel metal2 s 12806 39520 12862 40000 6 chany_top_out[5]
port 39 nsew default tristate
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_out[6]
port 40 nsew default tristate
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_out[7]
port 41 nsew default tristate
rlabel metal2 s 15474 39520 15530 40000 6 chany_top_out[8]
port 42 nsew default tristate
rlabel metal3 s 15520 30744 16000 30864 6 data_in
port 43 nsew default input
rlabel metal3 s 15520 1776 16000 1896 6 enable
port 44 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_grid_pin_0_
port 45 nsew default tristate
rlabel metal3 s 0 27344 480 27464 6 left_grid_pin_10_
port 46 nsew default tristate
rlabel metal3 s 0 32376 480 32496 6 left_grid_pin_12_
port 47 nsew default tristate
rlabel metal3 s 0 37408 480 37528 6 left_grid_pin_14_
port 48 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 left_grid_pin_2_
port 49 nsew default tristate
rlabel metal3 s 0 12384 480 12504 6 left_grid_pin_4_
port 50 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 left_grid_pin_6_
port 51 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 left_grid_pin_8_
port 52 nsew default tristate
rlabel metal3 s 15520 34416 16000 34536 6 right_grid_pin_3_
port 53 nsew default tristate
rlabel metal3 s 15520 38088 16000 38208 6 right_grid_pin_7_
port 54 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 55 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 56 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
