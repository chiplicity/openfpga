* NGSPICE file created from grid_io_bottom_bottom.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A Y VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B Z VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

.subckt grid_io_bottom_bottom IO_ISOL_N ccff_head ccff_tail gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] prog_clk
+ top_width_0_height_0__pin_0_ top_width_0_height_0__pin_10_ top_width_0_height_0__pin_11_lower
+ top_width_0_height_0__pin_11_upper top_width_0_height_0__pin_12_ top_width_0_height_0__pin_13_lower
+ top_width_0_height_0__pin_13_upper top_width_0_height_0__pin_14_ top_width_0_height_0__pin_15_lower
+ top_width_0_height_0__pin_15_upper top_width_0_height_0__pin_16_ top_width_0_height_0__pin_17_lower
+ top_width_0_height_0__pin_17_upper top_width_0_height_0__pin_1_lower top_width_0_height_0__pin_1_upper
+ top_width_0_height_0__pin_2_ top_width_0_height_0__pin_3_lower top_width_0_height_0__pin_3_upper
+ top_width_0_height_0__pin_4_ top_width_0_height_0__pin_5_lower top_width_0_height_0__pin_5_upper
+ top_width_0_height_0__pin_6_ top_width_0_height_0__pin_7_lower top_width_0_height_0__pin_7_upper
+ top_width_0_height_0__pin_8_ top_width_0_height_0__pin_9_lower top_width_0_height_0__pin_9_upper
+ VPWR VGND
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _04_/A
+ logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N _04_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
XFILLER_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A ccff_tail
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26_ top_width_0_height_0__pin_7_lower top_width_0_height_0__pin_7_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
X_09_ _09_/A gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _09_/A
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08_ _08_/A gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_25_ top_width_0_height_0__pin_5_lower top_width_0_height_0__pin_5_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N _06_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24_ top_width_0_height_0__pin_3_lower top_width_0_height_0__pin_3_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07_ _07_/A gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
+ logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y top_width_0_height_0__pin_13_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23_ top_width_0_height_0__pin_1_lower top_width_0_height_0__pin_1_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
+ logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y top_width_0_height_0__pin_7_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
X_06_ _06_/A gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_22_ top_width_0_height_0__pin_17_lower top_width_0_height_0__pin_17_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _05_/A
+ logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
X_05_ _05_/A gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y top_width_0_height_0__pin_1_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21_ top_width_0_height_0__pin_15_lower top_width_0_height_0__pin_15_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
X_04_ _04_/A gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N _08_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_03_ _03_/A gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_20_ top_width_0_height_0__pin_13_lower top_width_0_height_0__pin_13_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _01_/A
+ logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_02_ _02_/A gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_01_ _01_/A gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE ccff_tail
+ IO_ISOL_N _01_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
X_00_ top_width_0_height_0__pin_9_lower top_width_0_height_0__pin_9_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _06_/A
+ logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
XFILLER_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_0_
+ _09_/A _18_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N _03_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
+ logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y top_width_0_height_0__pin_17_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_2_
+ _08_/A _17_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
+ logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y top_width_0_height_0__pin_11_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _02_/A
+ logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
+ logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y top_width_0_height_0__pin_5_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_4_
+ _07_/A _16_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19_ top_width_0_height_0__pin_11_lower top_width_0_height_0__pin_11_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N _05_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
X_18_ _18_/A gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ccff_head logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_6_
+ _06_/A _15_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XPHY_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17_ _17_/A gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16_ _16_/A gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_8_
+ _05_/A _14_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _07_/A
+ logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
X_15_ _15_/A gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N _07_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14_ _14_/A gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_10_
+ _04_/A _13_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13_ _13_/A gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _03_/A
+ logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12_ _12_/A gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_12_
+ _03_/A _12_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11_ _11_/A gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_14_
+ _02_/A _11_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
X_10_ _10_/A gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N _09_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
XPHY_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
+ logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y top_width_0_height_0__pin_15_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XPHY_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
+ logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y top_width_0_height_0__pin_9_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_16_
+ _01_/A _10_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
+ logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y top_width_0_height_0__pin_3_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XPHY_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _08_/A
+ logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N _02_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
.ends

