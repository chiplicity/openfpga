VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__0_
  CLASS BLOCK ;
  FOREIGN sb_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 137.600 3.130 140.000 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 137.600 9.110 140.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 137.600 15.550 140.000 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 137.600 21.990 140.000 ;
    END
  END address[6]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 2.760 140.000 3.360 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 137.600 28.430 140.000 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.400 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 8.880 140.000 9.480 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 2.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 2.400 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 2.400 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 15.680 140.000 16.280 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 137.600 34.870 140.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 22.480 140.000 23.080 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 29.280 140.000 29.880 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 36.080 140.000 36.680 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 137.600 40.850 140.000 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 137.600 47.290 140.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 137.600 53.730 140.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 42.200 140.000 42.800 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 137.600 60.170 140.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 137.600 66.610 140.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 49.000 140.000 49.600 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 55.800 140.000 56.400 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 2.400 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 137.600 73.050 140.000 ;
    END
  END chanx_right_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.400 90.400 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 62.600 140.000 63.200 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 137.600 79.030 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.190 137.600 85.470 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 137.600 91.910 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 2.400 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 2.400 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 75.520 140.000 76.120 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 82.320 140.000 82.920 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 137.600 98.350 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 137.600 104.790 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.120 140.000 89.720 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 2.400 111.480 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 137.600 117.210 140.000 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 115.640 140.000 116.240 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.920 140.000 96.520 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 102.720 140.000 103.320 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 137.600 110.770 140.000 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 2.400 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 108.840 140.000 109.440 ;
    END
  END left_bottom_grid_pin_9_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 2.400 121.680 ;
    END
  END left_top_grid_pin_10_
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 2.400 131.880 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.240 140.000 129.840 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.040 140.000 136.640 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.370 137.600 123.650 140.000 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 2.400 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 2.400 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 122.440 140.000 123.040 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END right_bottom_grid_pin_9_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 137.600 130.090 140.000 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.250 137.600 136.530 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 2.400 137.320 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.070 0.380 138.850 137.660 ;
      LAYER met2 ;
        RECT 0.090 137.320 2.570 137.770 ;
        RECT 3.410 137.320 8.550 137.770 ;
        RECT 9.390 137.320 14.990 137.770 ;
        RECT 15.830 137.320 21.430 137.770 ;
        RECT 22.270 137.320 27.870 137.770 ;
        RECT 28.710 137.320 34.310 137.770 ;
        RECT 35.150 137.320 40.290 137.770 ;
        RECT 41.130 137.320 46.730 137.770 ;
        RECT 47.570 137.320 53.170 137.770 ;
        RECT 54.010 137.320 59.610 137.770 ;
        RECT 60.450 137.320 66.050 137.770 ;
        RECT 66.890 137.320 72.490 137.770 ;
        RECT 73.330 137.320 78.470 137.770 ;
        RECT 79.310 137.320 84.910 137.770 ;
        RECT 85.750 137.320 91.350 137.770 ;
        RECT 92.190 137.320 97.790 137.770 ;
        RECT 98.630 137.320 104.230 137.770 ;
        RECT 105.070 137.320 110.210 137.770 ;
        RECT 111.050 137.320 116.650 137.770 ;
        RECT 117.490 137.320 123.090 137.770 ;
        RECT 123.930 137.320 129.530 137.770 ;
        RECT 130.370 137.320 135.970 137.770 ;
        RECT 136.810 137.320 138.830 137.770 ;
        RECT 0.090 2.680 138.830 137.320 ;
        RECT 0.090 0.270 4.870 2.680 ;
        RECT 5.710 0.270 15.450 2.680 ;
        RECT 16.290 0.270 26.030 2.680 ;
        RECT 26.870 0.270 37.070 2.680 ;
        RECT 37.910 0.270 47.650 2.680 ;
        RECT 48.490 0.270 58.230 2.680 ;
        RECT 59.070 0.270 69.270 2.680 ;
        RECT 70.110 0.270 79.850 2.680 ;
        RECT 80.690 0.270 90.890 2.680 ;
        RECT 91.730 0.270 101.470 2.680 ;
        RECT 102.310 0.270 112.050 2.680 ;
        RECT 112.890 0.270 123.090 2.680 ;
        RECT 123.930 0.270 133.670 2.680 ;
        RECT 134.510 0.270 138.830 2.680 ;
      LAYER met3 ;
        RECT 2.800 136.320 137.200 136.720 ;
        RECT 0.270 135.640 137.200 136.320 ;
        RECT 0.270 132.280 138.650 135.640 ;
        RECT 2.800 130.880 138.650 132.280 ;
        RECT 0.270 130.240 138.650 130.880 ;
        RECT 0.270 128.840 137.200 130.240 ;
        RECT 0.270 127.520 138.650 128.840 ;
        RECT 2.800 126.120 138.650 127.520 ;
        RECT 0.270 123.440 138.650 126.120 ;
        RECT 0.270 122.080 137.200 123.440 ;
        RECT 2.800 122.040 137.200 122.080 ;
        RECT 2.800 120.680 138.650 122.040 ;
        RECT 0.270 116.640 138.650 120.680 ;
        RECT 2.800 115.240 137.200 116.640 ;
        RECT 0.270 111.880 138.650 115.240 ;
        RECT 2.800 110.480 138.650 111.880 ;
        RECT 0.270 109.840 138.650 110.480 ;
        RECT 0.270 108.440 137.200 109.840 ;
        RECT 0.270 106.440 138.650 108.440 ;
        RECT 2.800 105.040 138.650 106.440 ;
        RECT 0.270 103.720 138.650 105.040 ;
        RECT 0.270 102.320 137.200 103.720 ;
        RECT 0.270 101.000 138.650 102.320 ;
        RECT 2.800 99.600 138.650 101.000 ;
        RECT 0.270 96.920 138.650 99.600 ;
        RECT 0.270 96.240 137.200 96.920 ;
        RECT 2.800 95.520 137.200 96.240 ;
        RECT 2.800 94.840 138.650 95.520 ;
        RECT 0.270 90.800 138.650 94.840 ;
        RECT 2.800 90.120 138.650 90.800 ;
        RECT 2.800 89.400 137.200 90.120 ;
        RECT 0.270 88.720 137.200 89.400 ;
        RECT 0.270 86.040 138.650 88.720 ;
        RECT 2.800 84.640 138.650 86.040 ;
        RECT 0.270 83.320 138.650 84.640 ;
        RECT 0.270 81.920 137.200 83.320 ;
        RECT 0.270 80.600 138.650 81.920 ;
        RECT 2.800 79.200 138.650 80.600 ;
        RECT 0.270 76.520 138.650 79.200 ;
        RECT 0.270 75.160 137.200 76.520 ;
        RECT 2.800 75.120 137.200 75.160 ;
        RECT 2.800 73.760 138.650 75.120 ;
        RECT 0.270 70.400 138.650 73.760 ;
        RECT 2.800 69.000 137.200 70.400 ;
        RECT 0.270 64.960 138.650 69.000 ;
        RECT 2.800 63.600 138.650 64.960 ;
        RECT 2.800 63.560 137.200 63.600 ;
        RECT 0.270 62.200 137.200 63.560 ;
        RECT 0.270 59.520 138.650 62.200 ;
        RECT 2.800 58.120 138.650 59.520 ;
        RECT 0.270 56.800 138.650 58.120 ;
        RECT 0.270 55.400 137.200 56.800 ;
        RECT 0.270 54.760 138.650 55.400 ;
        RECT 2.800 53.360 138.650 54.760 ;
        RECT 0.270 50.000 138.650 53.360 ;
        RECT 0.270 49.320 137.200 50.000 ;
        RECT 2.800 48.600 137.200 49.320 ;
        RECT 2.800 47.920 138.650 48.600 ;
        RECT 0.270 44.560 138.650 47.920 ;
        RECT 2.800 43.200 138.650 44.560 ;
        RECT 2.800 43.160 137.200 43.200 ;
        RECT 0.270 41.800 137.200 43.160 ;
        RECT 0.270 39.120 138.650 41.800 ;
        RECT 2.800 37.720 138.650 39.120 ;
        RECT 0.270 37.080 138.650 37.720 ;
        RECT 0.270 35.680 137.200 37.080 ;
        RECT 0.270 33.680 138.650 35.680 ;
        RECT 2.800 32.280 138.650 33.680 ;
        RECT 0.270 30.280 138.650 32.280 ;
        RECT 0.270 28.920 137.200 30.280 ;
        RECT 2.800 28.880 137.200 28.920 ;
        RECT 2.800 27.520 138.650 28.880 ;
        RECT 0.270 23.480 138.650 27.520 ;
        RECT 2.800 22.080 137.200 23.480 ;
        RECT 0.270 18.040 138.650 22.080 ;
        RECT 2.800 16.680 138.650 18.040 ;
        RECT 2.800 16.640 137.200 16.680 ;
        RECT 0.270 15.280 137.200 16.640 ;
        RECT 0.270 13.280 138.650 15.280 ;
        RECT 2.800 11.880 138.650 13.280 ;
        RECT 0.270 9.880 138.650 11.880 ;
        RECT 0.270 8.480 137.200 9.880 ;
        RECT 0.270 7.840 138.650 8.480 ;
        RECT 2.800 6.440 138.650 7.840 ;
        RECT 0.270 3.760 138.650 6.440 ;
        RECT 0.270 3.080 137.200 3.760 ;
        RECT 2.800 2.680 137.200 3.080 ;
      LAYER met4 ;
        RECT 0.295 10.240 27.655 128.080 ;
        RECT 30.055 10.240 50.985 128.080 ;
        RECT 53.385 10.240 138.625 128.080 ;
        RECT 0.295 9.015 138.625 10.240 ;
      LAYER met5 ;
        RECT 92.580 62.100 118.100 63.700 ;
  END
END sb_1__0_
END LIBRARY

