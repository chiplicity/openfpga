magic
tech EFS8A
magscale 1 2
timestamp 1604399100
<< viali >>
rect 23489 24829 23523 24863
rect 23949 24489 23983 24523
rect 23765 24421 23799 24455
rect 24961 24421 24995 24455
rect 25513 24421 25547 24455
rect 23213 24353 23247 24387
rect 23857 24353 23891 24387
rect 23397 24285 23431 24319
rect 25145 24285 25179 24319
rect 16865 24081 16899 24115
rect 23489 24081 23523 24115
rect 10977 23945 11011 23979
rect 13993 23945 14027 23979
rect 16681 23945 16715 23979
rect 19892 23945 19926 23979
rect 24501 23945 24535 23979
rect 13737 23877 13771 23911
rect 19625 23877 19659 23911
rect 24593 23877 24627 23911
rect 24685 23877 24719 23911
rect 24133 23809 24167 23843
rect 11161 23741 11195 23775
rect 15117 23741 15151 23775
rect 16589 23741 16623 23775
rect 17233 23741 17267 23775
rect 19349 23741 19383 23775
rect 21005 23741 21039 23775
rect 23949 23741 23983 23775
rect 11713 23537 11747 23571
rect 12909 23537 12943 23571
rect 13921 23537 13955 23571
rect 14289 23537 14323 23571
rect 15485 23537 15519 23571
rect 16313 23537 16347 23571
rect 17877 23537 17911 23571
rect 18797 23537 18831 23571
rect 21465 23537 21499 23571
rect 23305 23537 23339 23571
rect 25145 23537 25179 23571
rect 25697 23537 25731 23571
rect 20269 23469 20303 23503
rect 16497 23401 16531 23435
rect 19901 23401 19935 23435
rect 22753 23401 22787 23435
rect 9689 23333 9723 23367
rect 10241 23333 10275 23367
rect 10793 23333 10827 23367
rect 11345 23333 11379 23367
rect 11897 23333 11931 23367
rect 12449 23333 12483 23367
rect 13001 23333 13035 23367
rect 13553 23333 13587 23367
rect 14105 23333 14139 23367
rect 14657 23333 14691 23367
rect 15301 23333 15335 23367
rect 15853 23333 15887 23367
rect 16764 23333 16798 23367
rect 19625 23333 19659 23367
rect 21281 23333 21315 23367
rect 23765 23333 23799 23367
rect 19073 23265 19107 23299
rect 19717 23265 19751 23299
rect 24032 23265 24066 23299
rect 9873 23197 9907 23231
rect 10977 23197 11011 23231
rect 12081 23197 12115 23231
rect 13185 23197 13219 23231
rect 19257 23197 19291 23231
rect 21833 23197 21867 23231
rect 23673 23197 23707 23231
rect 16405 22993 16439 23027
rect 18521 22993 18555 23027
rect 19349 22993 19383 23027
rect 23489 22993 23523 23027
rect 25053 22993 25087 23027
rect 19892 22925 19926 22959
rect 14197 22857 14231 22891
rect 14289 22857 14323 22891
rect 16773 22857 16807 22891
rect 18429 22857 18463 22891
rect 19625 22857 19659 22891
rect 22569 22857 22603 22891
rect 23940 22857 23974 22891
rect 14473 22789 14507 22823
rect 16865 22789 16899 22823
rect 16957 22789 16991 22823
rect 18613 22789 18647 22823
rect 23673 22789 23707 22823
rect 10885 22653 10919 22687
rect 13645 22653 13679 22687
rect 13829 22653 13863 22687
rect 16313 22653 16347 22687
rect 18061 22653 18095 22687
rect 21005 22653 21039 22687
rect 22017 22653 22051 22687
rect 22753 22653 22787 22687
rect 13553 22449 13587 22483
rect 14657 22449 14691 22483
rect 15853 22449 15887 22483
rect 17693 22449 17727 22483
rect 18613 22449 18647 22483
rect 18981 22449 19015 22483
rect 19717 22449 19751 22483
rect 20269 22449 20303 22483
rect 21097 22449 21131 22483
rect 16129 22381 16163 22415
rect 21741 22381 21775 22415
rect 12817 22313 12851 22347
rect 14105 22313 14139 22347
rect 14197 22313 14231 22347
rect 16313 22313 16347 22347
rect 21925 22313 21959 22347
rect 10701 22245 10735 22279
rect 10793 22245 10827 22279
rect 16580 22245 16614 22279
rect 20913 22245 20947 22279
rect 21373 22245 21407 22279
rect 22181 22245 22215 22279
rect 23857 22245 23891 22279
rect 24593 22245 24627 22279
rect 25145 22245 25179 22279
rect 11060 22177 11094 22211
rect 13185 22177 13219 22211
rect 14013 22177 14047 22211
rect 15025 22177 15059 22211
rect 12173 22109 12207 22143
rect 13645 22109 13679 22143
rect 18245 22109 18279 22143
rect 19809 22109 19843 22143
rect 23305 22109 23339 22143
rect 24225 22109 24259 22143
rect 24777 22109 24811 22143
rect 15025 21905 15059 21939
rect 16313 21905 16347 21939
rect 16773 21905 16807 21939
rect 20177 21905 20211 21939
rect 21741 21905 21775 21939
rect 22661 21905 22695 21939
rect 11161 21837 11195 21871
rect 13912 21837 13946 21871
rect 17325 21837 17359 21871
rect 18061 21769 18095 21803
rect 19717 21769 19751 21803
rect 24041 21769 24075 21803
rect 25237 21769 25271 21803
rect 11253 21701 11287 21735
rect 11345 21701 11379 21735
rect 13645 21701 13679 21735
rect 20269 21701 20303 21735
rect 20453 21701 20487 21735
rect 21833 21701 21867 21735
rect 22017 21701 22051 21735
rect 24133 21701 24167 21735
rect 24225 21701 24259 21735
rect 18245 21633 18279 21667
rect 19809 21633 19843 21667
rect 10609 21565 10643 21599
rect 10793 21565 10827 21599
rect 21373 21565 21407 21599
rect 23673 21565 23707 21599
rect 25421 21565 25455 21599
rect 10517 21361 10551 21395
rect 12081 21361 12115 21395
rect 13645 21361 13679 21395
rect 14105 21361 14139 21395
rect 17509 21361 17543 21395
rect 18153 21361 18187 21395
rect 20269 21361 20303 21395
rect 20729 21361 20763 21395
rect 22293 21361 22327 21395
rect 23305 21361 23339 21395
rect 23949 21361 23983 21395
rect 24225 21361 24259 21395
rect 25237 21361 25271 21395
rect 18337 21225 18371 21259
rect 20913 21225 20947 21259
rect 23397 21225 23431 21259
rect 10241 21157 10275 21191
rect 10701 21157 10735 21191
rect 24409 21157 24443 21191
rect 24869 21157 24903 21191
rect 10946 21089 10980 21123
rect 18582 21089 18616 21123
rect 21158 21089 21192 21123
rect 9689 21021 9723 21055
rect 14197 21021 14231 21055
rect 17785 21021 17819 21055
rect 19717 21021 19751 21055
rect 24593 21021 24627 21055
rect 10333 20817 10367 20851
rect 14197 20817 14231 20851
rect 18521 20817 18555 20851
rect 19533 20817 19567 20851
rect 21373 20817 21407 20851
rect 21741 20817 21775 20851
rect 22109 20817 22143 20851
rect 24685 20817 24719 20851
rect 11161 20681 11195 20715
rect 12449 20681 12483 20715
rect 14565 20681 14599 20715
rect 16773 20681 16807 20715
rect 18429 20681 18463 20715
rect 19993 20681 20027 20715
rect 25329 20681 25363 20715
rect 11253 20613 11287 20647
rect 11345 20613 11379 20647
rect 14657 20613 14691 20647
rect 14749 20613 14783 20647
rect 16865 20613 16899 20647
rect 17049 20613 17083 20647
rect 18613 20613 18647 20647
rect 20085 20613 20119 20647
rect 20177 20613 20211 20647
rect 20913 20613 20947 20647
rect 24777 20613 24811 20647
rect 24869 20613 24903 20647
rect 10793 20545 10827 20579
rect 12633 20545 12667 20579
rect 18061 20545 18095 20579
rect 10701 20477 10735 20511
rect 16221 20477 16255 20511
rect 16405 20477 16439 20511
rect 19165 20477 19199 20511
rect 19625 20477 19659 20511
rect 24317 20477 24351 20511
rect 10425 20273 10459 20307
rect 13369 20273 13403 20307
rect 14105 20273 14139 20307
rect 15025 20273 15059 20307
rect 16037 20273 16071 20307
rect 18245 20273 18279 20307
rect 19809 20273 19843 20307
rect 20085 20273 20119 20307
rect 20453 20273 20487 20307
rect 24685 20273 24719 20307
rect 25145 20273 25179 20307
rect 10149 20205 10183 20239
rect 14657 20205 14691 20239
rect 10793 20137 10827 20171
rect 18613 20137 18647 20171
rect 19165 20137 19199 20171
rect 19257 20137 19291 20171
rect 23213 20137 23247 20171
rect 24317 20137 24351 20171
rect 11345 20069 11379 20103
rect 11437 20069 11471 20103
rect 16221 20069 16255 20103
rect 19073 20069 19107 20103
rect 20913 20069 20947 20103
rect 21373 20069 21407 20103
rect 25237 20069 25271 20103
rect 11704 20001 11738 20035
rect 15761 20001 15795 20035
rect 16466 20001 16500 20035
rect 23489 20001 23523 20035
rect 24133 20001 24167 20035
rect 12817 19933 12851 19967
rect 14197 19933 14231 19967
rect 17601 19933 17635 19967
rect 18705 19933 18739 19967
rect 21097 19933 21131 19967
rect 22661 19933 22695 19967
rect 23673 19933 23707 19967
rect 24041 19933 24075 19967
rect 25421 19933 25455 19967
rect 25789 19933 25823 19967
rect 11253 19729 11287 19763
rect 13645 19729 13679 19763
rect 13921 19729 13955 19763
rect 15853 19729 15887 19763
rect 16405 19729 16439 19763
rect 16865 19729 16899 19763
rect 17785 19729 17819 19763
rect 18429 19729 18463 19763
rect 19441 19729 19475 19763
rect 19625 19729 19659 19763
rect 20177 19729 20211 19763
rect 11161 19661 11195 19695
rect 19073 19661 19107 19695
rect 13461 19593 13495 19627
rect 14729 19593 14763 19627
rect 21364 19593 21398 19627
rect 24041 19593 24075 19627
rect 24308 19593 24342 19627
rect 11437 19525 11471 19559
rect 12449 19525 12483 19559
rect 14473 19525 14507 19559
rect 18521 19525 18555 19559
rect 18613 19525 18647 19559
rect 21097 19525 21131 19559
rect 23949 19525 23983 19559
rect 10793 19389 10827 19423
rect 11805 19389 11839 19423
rect 17417 19389 17451 19423
rect 18061 19389 18095 19423
rect 21005 19389 21039 19423
rect 22477 19389 22511 19423
rect 25421 19389 25455 19423
rect 14657 19185 14691 19219
rect 23489 19185 23523 19219
rect 24593 19185 24627 19219
rect 11805 19049 11839 19083
rect 15945 19049 15979 19083
rect 18153 19049 18187 19083
rect 19809 19049 19843 19083
rect 24041 19049 24075 19083
rect 24225 19049 24259 19083
rect 10885 18981 10919 19015
rect 11621 18981 11655 19015
rect 12173 18981 12207 19015
rect 12725 18981 12759 19015
rect 12981 18981 13015 19015
rect 16681 18981 16715 19015
rect 18797 18981 18831 19015
rect 20913 18981 20947 19015
rect 21169 18981 21203 19015
rect 23949 18981 23983 19015
rect 24961 18981 24995 19015
rect 25145 18981 25179 19015
rect 25697 18981 25731 19015
rect 10517 18913 10551 18947
rect 11529 18913 11563 18947
rect 12633 18913 12667 18947
rect 15025 18913 15059 18947
rect 15761 18913 15795 18947
rect 17509 18913 17543 18947
rect 19717 18913 19751 18947
rect 20269 18913 20303 18947
rect 20637 18913 20671 18947
rect 23121 18913 23155 18947
rect 11161 18845 11195 18879
rect 14105 18845 14139 18879
rect 15301 18845 15335 18879
rect 15669 18845 15703 18879
rect 16405 18845 16439 18879
rect 17141 18845 17175 18879
rect 17601 18845 17635 18879
rect 17969 18845 18003 18879
rect 18061 18845 18095 18879
rect 19073 18845 19107 18879
rect 19257 18845 19291 18879
rect 19625 18845 19659 18879
rect 22293 18845 22327 18879
rect 23581 18845 23615 18879
rect 25329 18845 25363 18879
rect 11253 18641 11287 18675
rect 11621 18641 11655 18675
rect 12817 18641 12851 18675
rect 15301 18641 15335 18675
rect 15945 18641 15979 18675
rect 16957 18641 16991 18675
rect 17693 18641 17727 18675
rect 18521 18641 18555 18675
rect 19349 18641 19383 18675
rect 21465 18641 21499 18675
rect 21925 18641 21959 18675
rect 22477 18641 22511 18675
rect 24133 18641 24167 18675
rect 14565 18573 14599 18607
rect 18429 18573 18463 18607
rect 20821 18573 20855 18607
rect 23489 18573 23523 18607
rect 22385 18505 22419 18539
rect 23029 18505 23063 18539
rect 24041 18505 24075 18539
rect 25237 18505 25271 18539
rect 15393 18437 15427 18471
rect 15577 18437 15611 18471
rect 18613 18437 18647 18471
rect 20913 18437 20947 18471
rect 21097 18437 21131 18471
rect 22569 18437 22603 18471
rect 24317 18437 24351 18471
rect 23673 18369 23707 18403
rect 10885 18301 10919 18335
rect 13737 18301 13771 18335
rect 14933 18301 14967 18335
rect 18061 18301 18095 18335
rect 20453 18301 20487 18335
rect 22017 18301 22051 18335
rect 24685 18301 24719 18335
rect 25421 18301 25455 18335
rect 10977 18097 11011 18131
rect 12449 18097 12483 18131
rect 14933 18097 14967 18131
rect 16129 18097 16163 18131
rect 19073 18097 19107 18131
rect 20177 18097 20211 18131
rect 21465 18097 21499 18131
rect 24961 18097 24995 18131
rect 25697 18097 25731 18131
rect 15853 18029 15887 18063
rect 21189 18029 21223 18063
rect 23949 18029 23983 18063
rect 25421 18029 25455 18063
rect 11069 17961 11103 17995
rect 14197 17961 14231 17995
rect 21925 17961 21959 17995
rect 22937 17961 22971 17995
rect 24501 17961 24535 17995
rect 14013 17893 14047 17927
rect 15301 17893 15335 17927
rect 16497 17893 16531 17927
rect 17141 17893 17175 17927
rect 22753 17893 22787 17927
rect 23489 17893 23523 17927
rect 23857 17893 23891 17927
rect 24409 17893 24443 17927
rect 11314 17825 11348 17859
rect 13461 17825 13495 17859
rect 14105 17825 14139 17859
rect 17386 17825 17420 17859
rect 22201 17825 22235 17859
rect 22845 17825 22879 17859
rect 13645 17757 13679 17791
rect 15485 17757 15519 17791
rect 16957 17757 16991 17791
rect 18521 17757 18555 17791
rect 20545 17757 20579 17791
rect 22385 17757 22419 17791
rect 24317 17757 24351 17791
rect 13645 17553 13679 17587
rect 18613 17553 18647 17587
rect 21741 17553 21775 17587
rect 22477 17553 22511 17587
rect 22753 17553 22787 17587
rect 23213 17553 23247 17587
rect 23949 17553 23983 17587
rect 25513 17553 25547 17587
rect 14197 17485 14231 17519
rect 14534 17485 14568 17519
rect 18245 17485 18279 17519
rect 20913 17485 20947 17519
rect 21833 17485 21867 17519
rect 14289 17417 14323 17451
rect 20177 17417 20211 17451
rect 24400 17417 24434 17451
rect 20269 17349 20303 17383
rect 20361 17349 20395 17383
rect 21925 17349 21959 17383
rect 24133 17349 24167 17383
rect 19809 17281 19843 17315
rect 11161 17213 11195 17247
rect 15669 17213 15703 17247
rect 17233 17213 17267 17247
rect 21373 17213 21407 17247
rect 15025 17009 15059 17043
rect 18429 17009 18463 17043
rect 19165 17009 19199 17043
rect 19901 17009 19935 17043
rect 20913 17009 20947 17043
rect 24041 17009 24075 17043
rect 22661 16941 22695 16975
rect 25237 16941 25271 16975
rect 14105 16873 14139 16907
rect 14289 16873 14323 16907
rect 14657 16873 14691 16907
rect 15853 16873 15887 16907
rect 17049 16873 17083 16907
rect 20269 16873 20303 16907
rect 21465 16873 21499 16907
rect 23213 16873 23247 16907
rect 24685 16873 24719 16907
rect 24869 16873 24903 16907
rect 13553 16805 13587 16839
rect 15761 16805 15795 16839
rect 20729 16805 20763 16839
rect 21373 16805 21407 16839
rect 23029 16805 23063 16839
rect 23765 16805 23799 16839
rect 13185 16737 13219 16771
rect 14013 16737 14047 16771
rect 15669 16737 15703 16771
rect 16313 16737 16347 16771
rect 17294 16737 17328 16771
rect 21281 16737 21315 16771
rect 23121 16737 23155 16771
rect 13645 16669 13679 16703
rect 15301 16669 15335 16703
rect 16957 16669 16991 16703
rect 19441 16669 19475 16703
rect 21925 16669 21959 16703
rect 22569 16669 22603 16703
rect 24225 16669 24259 16703
rect 24593 16669 24627 16703
rect 13645 16465 13679 16499
rect 15485 16465 15519 16499
rect 16037 16465 16071 16499
rect 17141 16465 17175 16499
rect 21005 16465 21039 16499
rect 21925 16465 21959 16499
rect 24041 16465 24075 16499
rect 24777 16465 24811 16499
rect 25421 16465 25455 16499
rect 14372 16397 14406 16431
rect 19892 16397 19926 16431
rect 21649 16397 21683 16431
rect 25053 16397 25087 16431
rect 14105 16329 14139 16363
rect 22569 16329 22603 16363
rect 25237 16329 25271 16363
rect 19625 16261 19659 16295
rect 24133 16261 24167 16295
rect 24317 16261 24351 16295
rect 23213 16125 23247 16159
rect 23673 16125 23707 16159
rect 14105 15921 14139 15955
rect 14657 15921 14691 15955
rect 16865 15921 16899 15955
rect 18429 15921 18463 15955
rect 20269 15921 20303 15955
rect 23029 15921 23063 15955
rect 24501 15921 24535 15955
rect 25053 15921 25087 15955
rect 25789 15921 25823 15955
rect 25421 15853 25455 15887
rect 15301 15785 15335 15819
rect 17049 15785 17083 15819
rect 19809 15785 19843 15819
rect 21373 15785 21407 15819
rect 21465 15785 21499 15819
rect 23121 15785 23155 15819
rect 12081 15717 12115 15751
rect 12541 15717 12575 15751
rect 14197 15717 14231 15751
rect 15025 15717 15059 15751
rect 19625 15717 19659 15751
rect 17294 15649 17328 15683
rect 23388 15649 23422 15683
rect 12265 15581 12299 15615
rect 14381 15581 14415 15615
rect 20637 15581 20671 15615
rect 20913 15581 20947 15615
rect 21281 15581 21315 15615
rect 21925 15581 21959 15615
rect 12633 15377 12667 15411
rect 14841 15377 14875 15411
rect 17141 15377 17175 15411
rect 20545 15377 20579 15411
rect 21189 15377 21223 15411
rect 23397 15377 23431 15411
rect 24133 15377 24167 15411
rect 24685 15377 24719 15411
rect 25421 15377 25455 15411
rect 24041 15309 24075 15343
rect 12449 15241 12483 15275
rect 14657 15241 14691 15275
rect 19165 15241 19199 15275
rect 19432 15241 19466 15275
rect 25237 15241 25271 15275
rect 24317 15173 24351 15207
rect 23673 15105 23707 15139
rect 13001 15037 13035 15071
rect 15393 15037 15427 15071
rect 12081 14833 12115 14867
rect 12909 14833 12943 14867
rect 17233 14833 17267 14867
rect 19165 14833 19199 14867
rect 19533 14833 19567 14867
rect 21465 14833 21499 14867
rect 23397 14833 23431 14867
rect 23673 14833 23707 14867
rect 25237 14833 25271 14867
rect 14381 14765 14415 14799
rect 15301 14765 15335 14799
rect 24041 14765 24075 14799
rect 24777 14765 24811 14799
rect 13461 14697 13495 14731
rect 15853 14697 15887 14731
rect 17049 14629 17083 14663
rect 18061 14629 18095 14663
rect 18521 14629 18555 14663
rect 21281 14629 21315 14663
rect 21741 14629 21775 14663
rect 23489 14629 23523 14663
rect 24593 14629 24627 14663
rect 12817 14561 12851 14595
rect 13277 14561 13311 14595
rect 15117 14561 15151 14595
rect 15669 14561 15703 14595
rect 22937 14561 22971 14595
rect 12449 14493 12483 14527
rect 13369 14493 13403 14527
rect 14749 14493 14783 14527
rect 15761 14493 15795 14527
rect 17601 14493 17635 14527
rect 18245 14493 18279 14527
rect 24501 14493 24535 14527
rect 12725 14289 12759 14323
rect 16221 14289 16255 14323
rect 18061 14289 18095 14323
rect 21005 14289 21039 14323
rect 25053 14289 25087 14323
rect 13982 14221 14016 14255
rect 23918 14221 23952 14255
rect 13737 14153 13771 14187
rect 18429 14153 18463 14187
rect 21373 14153 21407 14187
rect 22569 14153 22603 14187
rect 23673 14153 23707 14187
rect 18521 14085 18555 14119
rect 18613 14085 18647 14119
rect 21465 14085 21499 14119
rect 21649 14085 21683 14119
rect 22293 14017 22327 14051
rect 15117 13949 15151 13983
rect 22753 13949 22787 13983
rect 13645 13745 13679 13779
rect 14565 13745 14599 13779
rect 16681 13745 16715 13779
rect 17325 13745 17359 13779
rect 21649 13745 21683 13779
rect 22109 13745 22143 13779
rect 24133 13745 24167 13779
rect 24869 13745 24903 13779
rect 14289 13677 14323 13711
rect 15025 13677 15059 13711
rect 17693 13677 17727 13711
rect 23581 13677 23615 13711
rect 24501 13677 24535 13711
rect 15301 13609 15335 13643
rect 21189 13609 21223 13643
rect 22201 13609 22235 13643
rect 11713 13541 11747 13575
rect 12081 13541 12115 13575
rect 12265 13541 12299 13575
rect 12532 13541 12566 13575
rect 15557 13541 15591 13575
rect 17785 13541 17819 13575
rect 18041 13541 18075 13575
rect 20361 13541 20395 13575
rect 24685 13541 24719 13575
rect 25237 13541 25271 13575
rect 20729 13473 20763 13507
rect 22446 13473 22480 13507
rect 19165 13405 19199 13439
rect 2789 13201 2823 13235
rect 12909 13201 12943 13235
rect 15485 13201 15519 13235
rect 17877 13201 17911 13235
rect 18061 13201 18095 13235
rect 18889 13201 18923 13235
rect 21925 13201 21959 13235
rect 22937 13201 22971 13235
rect 24777 13201 24811 13235
rect 15393 13133 15427 13167
rect 18613 13133 18647 13167
rect 19686 13133 19720 13167
rect 1409 13065 1443 13099
rect 1665 13065 1699 13099
rect 13277 13065 13311 13099
rect 15853 13065 15887 13099
rect 22293 13065 22327 13099
rect 24593 13065 24627 13099
rect 13369 12997 13403 13031
rect 13553 12997 13587 13031
rect 15945 12997 15979 13031
rect 16037 12997 16071 13031
rect 19441 12997 19475 13031
rect 22385 12997 22419 13031
rect 22477 12997 22511 13031
rect 20821 12861 20855 12895
rect 1593 12657 1627 12691
rect 2053 12657 2087 12691
rect 13001 12657 13035 12691
rect 13645 12657 13679 12691
rect 15577 12657 15611 12691
rect 16221 12657 16255 12691
rect 17969 12657 18003 12691
rect 19441 12657 19475 12691
rect 22293 12657 22327 12691
rect 23673 12657 23707 12691
rect 24501 12657 24535 12691
rect 19993 12589 20027 12623
rect 20637 12589 20671 12623
rect 24777 12589 24811 12623
rect 17601 12521 17635 12555
rect 20913 12521 20947 12555
rect 13369 12453 13403 12487
rect 15945 12453 15979 12487
rect 18061 12453 18095 12487
rect 18328 12453 18362 12487
rect 21169 12453 21203 12487
rect 22845 12453 22879 12487
rect 23489 12453 23523 12487
rect 24041 12453 24075 12487
rect 24593 12453 24627 12487
rect 25145 12385 25179 12419
rect 18245 12113 18279 12147
rect 19441 12113 19475 12147
rect 20913 12113 20947 12147
rect 22293 12113 22327 12147
rect 22753 12113 22787 12147
rect 24777 12113 24811 12147
rect 18613 11977 18647 12011
rect 22569 11977 22603 12011
rect 24593 11977 24627 12011
rect 18705 11909 18739 11943
rect 18889 11909 18923 11943
rect 22017 11909 22051 11943
rect 18613 11569 18647 11603
rect 19073 11569 19107 11603
rect 22569 11569 22603 11603
rect 23765 11569 23799 11603
rect 24501 11569 24535 11603
rect 24777 11569 24811 11603
rect 24041 11501 24075 11535
rect 25237 11433 25271 11467
rect 23581 11365 23615 11399
rect 24593 11365 24627 11399
rect 18337 11229 18371 11263
rect 24777 11025 24811 11059
rect 24593 10889 24627 10923
rect 24777 10481 24811 10515
rect 24501 10413 24535 10447
rect 24593 10277 24627 10311
rect 25237 10209 25271 10243
rect 24777 9937 24811 9971
rect 24593 9801 24627 9835
rect 24685 9393 24719 9427
rect 23949 9325 23983 9359
rect 23765 9189 23799 9223
rect 24409 9121 24443 9155
rect 24593 8849 24627 8883
rect 24409 8713 24443 8747
rect 24501 8305 24535 8339
rect 24777 7761 24811 7795
rect 24593 7625 24627 7659
rect 21189 7217 21223 7251
rect 24685 7217 24719 7251
rect 21005 7013 21039 7047
rect 21649 6877 21683 6911
rect 20361 6537 20395 6571
rect 20545 6401 20579 6435
rect 19809 6129 19843 6163
rect 20361 6129 20395 6163
rect 19625 5925 19659 5959
rect 19533 5789 19567 5823
rect 24777 5041 24811 5075
rect 25237 5041 25271 5075
rect 24593 4837 24627 4871
rect 24777 4497 24811 4531
rect 24593 4361 24627 4395
rect 24501 3953 24535 3987
rect 25237 3817 25271 3851
rect 24593 3749 24627 3783
rect 24777 3613 24811 3647
rect 16313 2865 16347 2899
rect 24777 2865 24811 2899
rect 16773 2729 16807 2763
rect 16129 2661 16163 2695
rect 24593 2661 24627 2695
rect 25145 2661 25179 2695
rect 24593 2185 24627 2219
rect 24777 2049 24811 2083
rect 25237 1981 25271 2015
<< metal1 >>
rect 19978 26248 19984 26300
rect 20036 26288 20042 26300
rect 24762 26288 24768 26300
rect 20036 26260 24768 26288
rect 20036 26248 20042 26260
rect 24762 26248 24768 26260
rect 24820 26248 24826 26300
rect 1104 25314 26864 25336
rect 1104 25262 10315 25314
rect 10367 25262 10379 25314
rect 10431 25262 10443 25314
rect 10495 25262 10507 25314
rect 10559 25262 19648 25314
rect 19700 25262 19712 25314
rect 19764 25262 19776 25314
rect 19828 25262 19840 25314
rect 19892 25262 26864 25314
rect 1104 25240 26864 25262
rect 23477 24863 23535 24869
rect 23477 24829 23489 24863
rect 23523 24860 23535 24863
rect 23934 24860 23940 24872
rect 23523 24832 23940 24860
rect 23523 24829 23535 24832
rect 23477 24823 23535 24829
rect 23934 24820 23940 24832
rect 23992 24820 23998 24872
rect 1104 24770 26864 24792
rect 1104 24718 5648 24770
rect 5700 24718 5712 24770
rect 5764 24718 5776 24770
rect 5828 24718 5840 24770
rect 5892 24718 14982 24770
rect 15034 24718 15046 24770
rect 15098 24718 15110 24770
rect 15162 24718 15174 24770
rect 15226 24718 24315 24770
rect 24367 24718 24379 24770
rect 24431 24718 24443 24770
rect 24495 24718 24507 24770
rect 24559 24718 26864 24770
rect 1104 24696 26864 24718
rect 21726 24548 21732 24600
rect 21784 24588 21790 24600
rect 24762 24588 24768 24600
rect 21784 24560 24768 24588
rect 21784 24548 21790 24560
rect 24762 24548 24768 24560
rect 24820 24548 24826 24600
rect 15286 24480 15292 24532
rect 15344 24520 15350 24532
rect 16482 24520 16488 24532
rect 15344 24492 16488 24520
rect 15344 24480 15350 24492
rect 16482 24480 16488 24492
rect 16540 24480 16546 24532
rect 17954 24480 17960 24532
rect 18012 24520 18018 24532
rect 18874 24520 18880 24532
rect 18012 24492 18880 24520
rect 18012 24480 18018 24492
rect 18874 24480 18880 24492
rect 18932 24480 18938 24532
rect 23934 24520 23940 24532
rect 23895 24492 23940 24520
rect 23934 24480 23940 24492
rect 23992 24480 23998 24532
rect 20714 24412 20720 24464
rect 20772 24452 20778 24464
rect 21266 24452 21272 24464
rect 20772 24424 21272 24452
rect 20772 24412 20778 24424
rect 21266 24412 21272 24424
rect 21324 24412 21330 24464
rect 23750 24452 23756 24464
rect 23711 24424 23756 24452
rect 23750 24412 23756 24424
rect 23808 24412 23814 24464
rect 24946 24452 24952 24464
rect 24907 24424 24952 24452
rect 24946 24412 24952 24424
rect 25004 24452 25010 24464
rect 25501 24455 25559 24461
rect 25501 24452 25513 24455
rect 25004 24424 25513 24452
rect 25004 24412 25010 24424
rect 25501 24421 25513 24424
rect 25547 24421 25559 24455
rect 25501 24415 25559 24421
rect 23198 24384 23204 24396
rect 23159 24356 23204 24384
rect 23198 24344 23204 24356
rect 23256 24384 23262 24396
rect 23845 24387 23903 24393
rect 23845 24384 23857 24387
rect 23256 24356 23857 24384
rect 23256 24344 23262 24356
rect 23845 24353 23857 24356
rect 23891 24353 23903 24387
rect 23845 24347 23903 24353
rect 23385 24319 23443 24325
rect 23385 24285 23397 24319
rect 23431 24316 23443 24319
rect 23566 24316 23572 24328
rect 23431 24288 23572 24316
rect 23431 24285 23443 24288
rect 23385 24279 23443 24285
rect 23566 24276 23572 24288
rect 23624 24276 23630 24328
rect 25130 24316 25136 24328
rect 25091 24288 25136 24316
rect 25130 24276 25136 24288
rect 25188 24276 25194 24328
rect 1104 24226 26864 24248
rect 1104 24174 10315 24226
rect 10367 24174 10379 24226
rect 10431 24174 10443 24226
rect 10495 24174 10507 24226
rect 10559 24174 19648 24226
rect 19700 24174 19712 24226
rect 19764 24174 19776 24226
rect 19828 24174 19840 24226
rect 19892 24174 26864 24226
rect 1104 24152 26864 24174
rect 16853 24115 16911 24121
rect 16853 24081 16865 24115
rect 16899 24112 16911 24115
rect 17310 24112 17316 24124
rect 16899 24084 17316 24112
rect 16899 24081 16911 24084
rect 16853 24075 16911 24081
rect 17310 24072 17316 24084
rect 17368 24072 17374 24124
rect 23477 24115 23535 24121
rect 23477 24081 23489 24115
rect 23523 24112 23535 24115
rect 23750 24112 23756 24124
rect 23523 24084 23756 24112
rect 23523 24081 23535 24084
rect 23477 24075 23535 24081
rect 23750 24072 23756 24084
rect 23808 24072 23814 24124
rect 23842 24072 23848 24124
rect 23900 24112 23906 24124
rect 24210 24112 24216 24124
rect 23900 24084 24216 24112
rect 23900 24072 23906 24084
rect 24210 24072 24216 24084
rect 24268 24072 24274 24124
rect 19334 24004 19340 24056
rect 19392 24044 19398 24056
rect 20438 24044 20444 24056
rect 19392 24016 20444 24044
rect 19392 24004 19398 24016
rect 20438 24004 20444 24016
rect 20496 24004 20502 24056
rect 10965 23979 11023 23985
rect 10965 23945 10977 23979
rect 11011 23976 11023 23979
rect 11146 23976 11152 23988
rect 11011 23948 11152 23976
rect 11011 23945 11023 23948
rect 10965 23939 11023 23945
rect 11146 23936 11152 23948
rect 11204 23936 11210 23988
rect 12894 23936 12900 23988
rect 12952 23976 12958 23988
rect 13981 23979 14039 23985
rect 13981 23976 13993 23979
rect 12952 23948 13993 23976
rect 12952 23936 12958 23948
rect 13981 23945 13993 23948
rect 14027 23976 14039 23979
rect 15102 23976 15108 23988
rect 14027 23948 15108 23976
rect 14027 23945 14039 23948
rect 13981 23939 14039 23945
rect 15102 23936 15108 23948
rect 15160 23936 15166 23988
rect 16669 23979 16727 23985
rect 16669 23945 16681 23979
rect 16715 23976 16727 23979
rect 17218 23976 17224 23988
rect 16715 23948 17224 23976
rect 16715 23945 16727 23948
rect 16669 23939 16727 23945
rect 17218 23936 17224 23948
rect 17276 23936 17282 23988
rect 19886 23985 19892 23988
rect 19880 23976 19892 23985
rect 19847 23948 19892 23976
rect 19880 23939 19892 23948
rect 19886 23936 19892 23939
rect 19944 23936 19950 23988
rect 23290 23936 23296 23988
rect 23348 23976 23354 23988
rect 24489 23979 24547 23985
rect 24489 23976 24501 23979
rect 23348 23948 24501 23976
rect 23348 23936 23354 23948
rect 24489 23945 24501 23948
rect 24535 23945 24547 23979
rect 24489 23939 24547 23945
rect 13722 23908 13728 23920
rect 13683 23880 13728 23908
rect 13722 23868 13728 23880
rect 13780 23868 13786 23920
rect 19610 23908 19616 23920
rect 19571 23880 19616 23908
rect 19610 23868 19616 23880
rect 19668 23868 19674 23920
rect 23566 23868 23572 23920
rect 23624 23908 23630 23920
rect 24581 23911 24639 23917
rect 24581 23908 24593 23911
rect 23624 23880 24593 23908
rect 23624 23868 23630 23880
rect 24581 23877 24593 23880
rect 24627 23877 24639 23911
rect 24581 23871 24639 23877
rect 24670 23868 24676 23920
rect 24728 23908 24734 23920
rect 24728 23880 24773 23908
rect 24728 23868 24734 23880
rect 23750 23800 23756 23852
rect 23808 23840 23814 23852
rect 24121 23843 24179 23849
rect 24121 23840 24133 23843
rect 23808 23812 24133 23840
rect 23808 23800 23814 23812
rect 24121 23809 24133 23812
rect 24167 23809 24179 23843
rect 24121 23803 24179 23809
rect 11149 23775 11207 23781
rect 11149 23741 11161 23775
rect 11195 23772 11207 23775
rect 12342 23772 12348 23784
rect 11195 23744 12348 23772
rect 11195 23741 11207 23744
rect 11149 23735 11207 23741
rect 12342 23732 12348 23744
rect 12400 23732 12406 23784
rect 14458 23732 14464 23784
rect 14516 23772 14522 23784
rect 15105 23775 15163 23781
rect 15105 23772 15117 23775
rect 14516 23744 15117 23772
rect 14516 23732 14522 23744
rect 15105 23741 15117 23744
rect 15151 23741 15163 23775
rect 15105 23735 15163 23741
rect 16577 23775 16635 23781
rect 16577 23741 16589 23775
rect 16623 23772 16635 23775
rect 16758 23772 16764 23784
rect 16623 23744 16764 23772
rect 16623 23741 16635 23744
rect 16577 23735 16635 23741
rect 16758 23732 16764 23744
rect 16816 23732 16822 23784
rect 17218 23772 17224 23784
rect 17179 23744 17224 23772
rect 17218 23732 17224 23744
rect 17276 23732 17282 23784
rect 19337 23775 19395 23781
rect 19337 23741 19349 23775
rect 19383 23772 19395 23775
rect 19886 23772 19892 23784
rect 19383 23744 19892 23772
rect 19383 23741 19395 23744
rect 19337 23735 19395 23741
rect 19886 23732 19892 23744
rect 19944 23772 19950 23784
rect 20993 23775 21051 23781
rect 20993 23772 21005 23775
rect 19944 23744 21005 23772
rect 19944 23732 19950 23744
rect 20993 23741 21005 23744
rect 21039 23741 21051 23775
rect 20993 23735 21051 23741
rect 23937 23775 23995 23781
rect 23937 23741 23949 23775
rect 23983 23772 23995 23775
rect 24026 23772 24032 23784
rect 23983 23744 24032 23772
rect 23983 23741 23995 23744
rect 23937 23735 23995 23741
rect 24026 23732 24032 23744
rect 24084 23732 24090 23784
rect 1104 23682 26864 23704
rect 1104 23630 5648 23682
rect 5700 23630 5712 23682
rect 5764 23630 5776 23682
rect 5828 23630 5840 23682
rect 5892 23630 14982 23682
rect 15034 23630 15046 23682
rect 15098 23630 15110 23682
rect 15162 23630 15174 23682
rect 15226 23630 24315 23682
rect 24367 23630 24379 23682
rect 24431 23630 24443 23682
rect 24495 23630 24507 23682
rect 24559 23630 26864 23682
rect 1104 23608 26864 23630
rect 11146 23528 11152 23580
rect 11204 23568 11210 23580
rect 11701 23571 11759 23577
rect 11701 23568 11713 23571
rect 11204 23540 11713 23568
rect 11204 23528 11210 23540
rect 11701 23537 11713 23540
rect 11747 23537 11759 23571
rect 12894 23568 12900 23580
rect 12855 23540 12900 23568
rect 11701 23531 11759 23537
rect 12894 23528 12900 23540
rect 12952 23528 12958 23580
rect 13722 23528 13728 23580
rect 13780 23568 13786 23580
rect 13909 23571 13967 23577
rect 13909 23568 13921 23571
rect 13780 23540 13921 23568
rect 13780 23528 13786 23540
rect 13909 23537 13921 23540
rect 13955 23537 13967 23571
rect 13909 23531 13967 23537
rect 14277 23571 14335 23577
rect 14277 23537 14289 23571
rect 14323 23568 14335 23571
rect 14550 23568 14556 23580
rect 14323 23540 14556 23568
rect 14323 23537 14335 23540
rect 14277 23531 14335 23537
rect 13924 23500 13952 23531
rect 14550 23528 14556 23540
rect 14608 23528 14614 23580
rect 15473 23571 15531 23577
rect 15473 23537 15485 23571
rect 15519 23568 15531 23571
rect 15930 23568 15936 23580
rect 15519 23540 15936 23568
rect 15519 23537 15531 23540
rect 15473 23531 15531 23537
rect 15930 23528 15936 23540
rect 15988 23528 15994 23580
rect 16298 23568 16304 23580
rect 16040 23540 16304 23568
rect 16040 23500 16068 23540
rect 16298 23528 16304 23540
rect 16356 23568 16362 23580
rect 17862 23568 17868 23580
rect 16356 23540 16528 23568
rect 17823 23540 17868 23568
rect 16356 23528 16362 23540
rect 13924 23472 16068 23500
rect 16500 23441 16528 23540
rect 17862 23528 17868 23540
rect 17920 23528 17926 23580
rect 18785 23571 18843 23577
rect 18785 23537 18797 23571
rect 18831 23568 18843 23571
rect 19794 23568 19800 23580
rect 18831 23540 19800 23568
rect 18831 23537 18843 23540
rect 18785 23531 18843 23537
rect 19794 23528 19800 23540
rect 19852 23528 19858 23580
rect 21453 23571 21511 23577
rect 21453 23537 21465 23571
rect 21499 23568 21511 23571
rect 22738 23568 22744 23580
rect 21499 23540 22744 23568
rect 21499 23537 21511 23540
rect 21453 23531 21511 23537
rect 22738 23528 22744 23540
rect 22796 23528 22802 23580
rect 23290 23568 23296 23580
rect 23251 23540 23296 23568
rect 23290 23528 23296 23540
rect 23348 23528 23354 23580
rect 23658 23528 23664 23580
rect 23716 23568 23722 23580
rect 23934 23568 23940 23580
rect 23716 23540 23940 23568
rect 23716 23528 23722 23540
rect 23934 23528 23940 23540
rect 23992 23528 23998 23580
rect 24670 23528 24676 23580
rect 24728 23568 24734 23580
rect 25133 23571 25191 23577
rect 25133 23568 25145 23571
rect 24728 23540 25145 23568
rect 24728 23528 24734 23540
rect 25133 23537 25145 23540
rect 25179 23568 25191 23571
rect 25685 23571 25743 23577
rect 25685 23568 25697 23571
rect 25179 23540 25697 23568
rect 25179 23537 25191 23540
rect 25133 23531 25191 23537
rect 25685 23537 25697 23540
rect 25731 23537 25743 23571
rect 25685 23531 25743 23537
rect 19610 23460 19616 23512
rect 19668 23500 19674 23512
rect 20162 23500 20168 23512
rect 19668 23472 20168 23500
rect 19668 23460 19674 23472
rect 20162 23460 20168 23472
rect 20220 23500 20226 23512
rect 20257 23503 20315 23509
rect 20257 23500 20269 23503
rect 20220 23472 20269 23500
rect 20220 23460 20226 23472
rect 20257 23469 20269 23472
rect 20303 23469 20315 23503
rect 20257 23463 20315 23469
rect 16485 23435 16543 23441
rect 16485 23401 16497 23435
rect 16531 23401 16543 23435
rect 19886 23432 19892 23444
rect 19847 23404 19892 23432
rect 16485 23395 16543 23401
rect 19886 23392 19892 23404
rect 19944 23392 19950 23444
rect 22741 23435 22799 23441
rect 22741 23401 22753 23435
rect 22787 23432 22799 23435
rect 23308 23432 23336 23528
rect 22787 23404 23336 23432
rect 22787 23401 22799 23404
rect 22741 23395 22799 23401
rect 9677 23367 9735 23373
rect 9677 23333 9689 23367
rect 9723 23364 9735 23367
rect 9766 23364 9772 23376
rect 9723 23336 9772 23364
rect 9723 23333 9735 23336
rect 9677 23327 9735 23333
rect 9766 23324 9772 23336
rect 9824 23364 9830 23376
rect 10229 23367 10287 23373
rect 10229 23364 10241 23367
rect 9824 23336 10241 23364
rect 9824 23324 9830 23336
rect 10229 23333 10241 23336
rect 10275 23333 10287 23367
rect 10778 23364 10784 23376
rect 10739 23336 10784 23364
rect 10229 23327 10287 23333
rect 10778 23324 10784 23336
rect 10836 23364 10842 23376
rect 11333 23367 11391 23373
rect 11333 23364 11345 23367
rect 10836 23336 11345 23364
rect 10836 23324 10842 23336
rect 11333 23333 11345 23336
rect 11379 23333 11391 23367
rect 11882 23364 11888 23376
rect 11843 23336 11888 23364
rect 11333 23327 11391 23333
rect 11882 23324 11888 23336
rect 11940 23364 11946 23376
rect 12437 23367 12495 23373
rect 12437 23364 12449 23367
rect 11940 23336 12449 23364
rect 11940 23324 11946 23336
rect 12437 23333 12449 23336
rect 12483 23333 12495 23367
rect 12437 23327 12495 23333
rect 12526 23324 12532 23376
rect 12584 23364 12590 23376
rect 12989 23367 13047 23373
rect 12989 23364 13001 23367
rect 12584 23336 13001 23364
rect 12584 23324 12590 23336
rect 12989 23333 13001 23336
rect 13035 23364 13047 23367
rect 13541 23367 13599 23373
rect 13541 23364 13553 23367
rect 13035 23336 13553 23364
rect 13035 23333 13047 23336
rect 12989 23327 13047 23333
rect 13541 23333 13553 23336
rect 13587 23333 13599 23367
rect 14090 23364 14096 23376
rect 14051 23336 14096 23364
rect 13541 23327 13599 23333
rect 14090 23324 14096 23336
rect 14148 23364 14154 23376
rect 14645 23367 14703 23373
rect 14645 23364 14657 23367
rect 14148 23336 14657 23364
rect 14148 23324 14154 23336
rect 14645 23333 14657 23336
rect 14691 23333 14703 23367
rect 15286 23364 15292 23376
rect 15247 23336 15292 23364
rect 14645 23327 14703 23333
rect 15286 23324 15292 23336
rect 15344 23364 15350 23376
rect 16758 23373 16764 23376
rect 15841 23367 15899 23373
rect 15841 23364 15853 23367
rect 15344 23336 15853 23364
rect 15344 23324 15350 23336
rect 15841 23333 15853 23336
rect 15887 23333 15899 23367
rect 16752 23364 16764 23373
rect 16719 23336 16764 23364
rect 15841 23327 15899 23333
rect 16752 23327 16764 23336
rect 16758 23324 16764 23327
rect 16816 23324 16822 23376
rect 19426 23324 19432 23376
rect 19484 23364 19490 23376
rect 19613 23367 19671 23373
rect 19613 23364 19625 23367
rect 19484 23336 19625 23364
rect 19484 23324 19490 23336
rect 19613 23333 19625 23336
rect 19659 23364 19671 23367
rect 19978 23364 19984 23376
rect 19659 23336 19984 23364
rect 19659 23333 19671 23336
rect 19613 23327 19671 23333
rect 19978 23324 19984 23336
rect 20036 23364 20042 23376
rect 20346 23364 20352 23376
rect 20036 23336 20352 23364
rect 20036 23324 20042 23336
rect 20346 23324 20352 23336
rect 20404 23324 20410 23376
rect 21269 23367 21327 23373
rect 21269 23333 21281 23367
rect 21315 23364 21327 23367
rect 23753 23367 23811 23373
rect 23753 23364 23765 23367
rect 21315 23336 21588 23364
rect 21315 23333 21327 23336
rect 21269 23327 21327 23333
rect 19058 23296 19064 23308
rect 19019 23268 19064 23296
rect 19058 23256 19064 23268
rect 19116 23296 19122 23308
rect 19705 23299 19763 23305
rect 19705 23296 19717 23299
rect 19116 23268 19717 23296
rect 19116 23256 19122 23268
rect 19705 23265 19717 23268
rect 19751 23265 19763 23299
rect 19705 23259 19763 23265
rect 21560 23240 21588 23336
rect 23676 23336 23765 23364
rect 23676 23240 23704 23336
rect 23753 23333 23765 23336
rect 23799 23333 23811 23367
rect 23753 23327 23811 23333
rect 24026 23305 24032 23308
rect 24020 23259 24032 23305
rect 24084 23296 24090 23308
rect 25038 23296 25044 23308
rect 24084 23268 25044 23296
rect 24026 23256 24032 23259
rect 24084 23256 24090 23268
rect 25038 23256 25044 23268
rect 25096 23256 25102 23308
rect 9858 23228 9864 23240
rect 9819 23200 9864 23228
rect 9858 23188 9864 23200
rect 9916 23188 9922 23240
rect 10962 23228 10968 23240
rect 10923 23200 10968 23228
rect 10962 23188 10968 23200
rect 11020 23188 11026 23240
rect 12066 23228 12072 23240
rect 12027 23200 12072 23228
rect 12066 23188 12072 23200
rect 12124 23188 12130 23240
rect 13173 23231 13231 23237
rect 13173 23197 13185 23231
rect 13219 23228 13231 23231
rect 14274 23228 14280 23240
rect 13219 23200 14280 23228
rect 13219 23197 13231 23200
rect 13173 23191 13231 23197
rect 14274 23188 14280 23200
rect 14332 23188 14338 23240
rect 19245 23231 19303 23237
rect 19245 23197 19257 23231
rect 19291 23228 19303 23231
rect 19334 23228 19340 23240
rect 19291 23200 19340 23228
rect 19291 23197 19303 23200
rect 19245 23191 19303 23197
rect 19334 23188 19340 23200
rect 19392 23188 19398 23240
rect 21542 23188 21548 23240
rect 21600 23228 21606 23240
rect 21821 23231 21879 23237
rect 21821 23228 21833 23231
rect 21600 23200 21833 23228
rect 21600 23188 21606 23200
rect 21821 23197 21833 23200
rect 21867 23197 21879 23231
rect 23658 23228 23664 23240
rect 23619 23200 23664 23228
rect 21821 23191 21879 23197
rect 23658 23188 23664 23200
rect 23716 23188 23722 23240
rect 1104 23138 26864 23160
rect 1104 23086 10315 23138
rect 10367 23086 10379 23138
rect 10431 23086 10443 23138
rect 10495 23086 10507 23138
rect 10559 23086 19648 23138
rect 19700 23086 19712 23138
rect 19764 23086 19776 23138
rect 19828 23086 19840 23138
rect 19892 23086 26864 23138
rect 1104 23064 26864 23086
rect 16393 23027 16451 23033
rect 16393 22993 16405 23027
rect 16439 23024 16451 23027
rect 18509 23027 18567 23033
rect 18509 23024 18521 23027
rect 16439 22996 18521 23024
rect 16439 22993 16451 22996
rect 16393 22987 16451 22993
rect 18509 22993 18521 22996
rect 18555 23024 18567 23027
rect 18966 23024 18972 23036
rect 18555 22996 18972 23024
rect 18555 22993 18567 22996
rect 18509 22987 18567 22993
rect 18966 22984 18972 22996
rect 19024 22984 19030 23036
rect 19337 23027 19395 23033
rect 19337 22993 19349 23027
rect 19383 23024 19395 23027
rect 19426 23024 19432 23036
rect 19383 22996 19432 23024
rect 19383 22993 19395 22996
rect 19337 22987 19395 22993
rect 19426 22984 19432 22996
rect 19484 22984 19490 23036
rect 23477 23027 23535 23033
rect 23477 22993 23489 23027
rect 23523 23024 23535 23027
rect 23566 23024 23572 23036
rect 23523 22996 23572 23024
rect 23523 22993 23535 22996
rect 23477 22987 23535 22993
rect 23566 22984 23572 22996
rect 23624 22984 23630 23036
rect 25038 23024 25044 23036
rect 24999 22996 25044 23024
rect 25038 22984 25044 22996
rect 25096 22984 25102 23036
rect 19880 22959 19938 22965
rect 19880 22925 19892 22959
rect 19926 22956 19938 22959
rect 19978 22956 19984 22968
rect 19926 22928 19984 22956
rect 19926 22925 19938 22928
rect 19880 22919 19938 22925
rect 19978 22916 19984 22928
rect 20036 22916 20042 22968
rect 14182 22888 14188 22900
rect 14143 22860 14188 22888
rect 14182 22848 14188 22860
rect 14240 22848 14246 22900
rect 14274 22848 14280 22900
rect 14332 22888 14338 22900
rect 16761 22891 16819 22897
rect 14332 22860 14377 22888
rect 14332 22848 14338 22860
rect 16761 22857 16773 22891
rect 16807 22888 16819 22891
rect 17494 22888 17500 22900
rect 16807 22860 17500 22888
rect 16807 22857 16819 22860
rect 16761 22851 16819 22857
rect 17494 22848 17500 22860
rect 17552 22848 17558 22900
rect 18230 22848 18236 22900
rect 18288 22888 18294 22900
rect 18417 22891 18475 22897
rect 18417 22888 18429 22891
rect 18288 22860 18429 22888
rect 18288 22848 18294 22860
rect 18417 22857 18429 22860
rect 18463 22857 18475 22891
rect 18417 22851 18475 22857
rect 19613 22891 19671 22897
rect 19613 22857 19625 22891
rect 19659 22888 19671 22891
rect 19702 22888 19708 22900
rect 19659 22860 19708 22888
rect 19659 22857 19671 22860
rect 19613 22851 19671 22857
rect 19702 22848 19708 22860
rect 19760 22888 19766 22900
rect 20162 22888 20168 22900
rect 19760 22860 20168 22888
rect 19760 22848 19766 22860
rect 20162 22848 20168 22860
rect 20220 22848 20226 22900
rect 22557 22891 22615 22897
rect 22557 22857 22569 22891
rect 22603 22888 22615 22891
rect 22646 22888 22652 22900
rect 22603 22860 22652 22888
rect 22603 22857 22615 22860
rect 22557 22851 22615 22857
rect 22646 22848 22652 22860
rect 22704 22888 22710 22900
rect 23750 22888 23756 22900
rect 22704 22860 23756 22888
rect 22704 22848 22710 22860
rect 23750 22848 23756 22860
rect 23808 22848 23814 22900
rect 23928 22891 23986 22897
rect 23928 22857 23940 22891
rect 23974 22888 23986 22891
rect 24210 22888 24216 22900
rect 23974 22860 24216 22888
rect 23974 22857 23986 22860
rect 23928 22851 23986 22857
rect 24210 22848 24216 22860
rect 24268 22848 24274 22900
rect 14090 22780 14096 22832
rect 14148 22820 14154 22832
rect 14458 22820 14464 22832
rect 14148 22792 14464 22820
rect 14148 22780 14154 22792
rect 14458 22780 14464 22792
rect 14516 22780 14522 22832
rect 16114 22780 16120 22832
rect 16172 22820 16178 22832
rect 16853 22823 16911 22829
rect 16853 22820 16865 22823
rect 16172 22792 16865 22820
rect 16172 22780 16178 22792
rect 16853 22789 16865 22792
rect 16899 22789 16911 22823
rect 16853 22783 16911 22789
rect 16945 22823 17003 22829
rect 16945 22789 16957 22823
rect 16991 22789 17003 22823
rect 16945 22783 17003 22789
rect 16758 22712 16764 22764
rect 16816 22752 16822 22764
rect 16960 22752 16988 22783
rect 17954 22780 17960 22832
rect 18012 22820 18018 22832
rect 18598 22820 18604 22832
rect 18012 22792 18604 22820
rect 18012 22780 18018 22792
rect 18598 22780 18604 22792
rect 18656 22780 18662 22832
rect 23658 22820 23664 22832
rect 23619 22792 23664 22820
rect 23658 22780 23664 22792
rect 23716 22780 23722 22832
rect 17678 22752 17684 22764
rect 16816 22724 17684 22752
rect 16816 22712 16822 22724
rect 17678 22712 17684 22724
rect 17736 22712 17742 22764
rect 10873 22687 10931 22693
rect 10873 22653 10885 22687
rect 10919 22684 10931 22687
rect 11330 22684 11336 22696
rect 10919 22656 11336 22684
rect 10919 22653 10931 22656
rect 10873 22647 10931 22653
rect 11330 22644 11336 22656
rect 11388 22644 11394 22696
rect 13630 22684 13636 22696
rect 13591 22656 13636 22684
rect 13630 22644 13636 22656
rect 13688 22644 13694 22696
rect 13814 22684 13820 22696
rect 13775 22656 13820 22684
rect 13814 22644 13820 22656
rect 13872 22644 13878 22696
rect 16301 22687 16359 22693
rect 16301 22653 16313 22687
rect 16347 22684 16359 22687
rect 16850 22684 16856 22696
rect 16347 22656 16856 22684
rect 16347 22653 16359 22656
rect 16301 22647 16359 22653
rect 16850 22644 16856 22656
rect 16908 22644 16914 22696
rect 18046 22684 18052 22696
rect 18007 22656 18052 22684
rect 18046 22644 18052 22656
rect 18104 22644 18110 22696
rect 20530 22644 20536 22696
rect 20588 22684 20594 22696
rect 20993 22687 21051 22693
rect 20993 22684 21005 22687
rect 20588 22656 21005 22684
rect 20588 22644 20594 22656
rect 20993 22653 21005 22656
rect 21039 22653 21051 22687
rect 22002 22684 22008 22696
rect 21963 22656 22008 22684
rect 20993 22647 21051 22653
rect 22002 22644 22008 22656
rect 22060 22644 22066 22696
rect 22738 22684 22744 22696
rect 22699 22656 22744 22684
rect 22738 22644 22744 22656
rect 22796 22644 22802 22696
rect 1104 22594 26864 22616
rect 1104 22542 5648 22594
rect 5700 22542 5712 22594
rect 5764 22542 5776 22594
rect 5828 22542 5840 22594
rect 5892 22542 14982 22594
rect 15034 22542 15046 22594
rect 15098 22542 15110 22594
rect 15162 22542 15174 22594
rect 15226 22542 24315 22594
rect 24367 22542 24379 22594
rect 24431 22542 24443 22594
rect 24495 22542 24507 22594
rect 24559 22542 26864 22594
rect 1104 22520 26864 22542
rect 13538 22480 13544 22492
rect 13451 22452 13544 22480
rect 13538 22440 13544 22452
rect 13596 22480 13602 22492
rect 14182 22480 14188 22492
rect 13596 22452 14188 22480
rect 13596 22440 13602 22452
rect 14182 22440 14188 22452
rect 14240 22440 14246 22492
rect 14274 22440 14280 22492
rect 14332 22480 14338 22492
rect 14645 22483 14703 22489
rect 14645 22480 14657 22483
rect 14332 22452 14657 22480
rect 14332 22440 14338 22452
rect 14645 22449 14657 22452
rect 14691 22449 14703 22483
rect 14645 22443 14703 22449
rect 15841 22483 15899 22489
rect 15841 22449 15853 22483
rect 15887 22480 15899 22483
rect 17494 22480 17500 22492
rect 15887 22452 17500 22480
rect 15887 22449 15899 22452
rect 15841 22443 15899 22449
rect 17494 22440 17500 22452
rect 17552 22440 17558 22492
rect 17678 22480 17684 22492
rect 17639 22452 17684 22480
rect 17678 22440 17684 22452
rect 17736 22440 17742 22492
rect 18598 22480 18604 22492
rect 18559 22452 18604 22480
rect 18598 22440 18604 22452
rect 18656 22440 18662 22492
rect 18966 22480 18972 22492
rect 18927 22452 18972 22480
rect 18966 22440 18972 22452
rect 19024 22440 19030 22492
rect 19426 22440 19432 22492
rect 19484 22480 19490 22492
rect 19702 22480 19708 22492
rect 19484 22452 19708 22480
rect 19484 22440 19490 22452
rect 19702 22440 19708 22452
rect 19760 22440 19766 22492
rect 19978 22440 19984 22492
rect 20036 22480 20042 22492
rect 20257 22483 20315 22489
rect 20257 22480 20269 22483
rect 20036 22452 20269 22480
rect 20036 22440 20042 22452
rect 20257 22449 20269 22452
rect 20303 22449 20315 22483
rect 20257 22443 20315 22449
rect 21085 22483 21143 22489
rect 21085 22449 21097 22483
rect 21131 22480 21143 22483
rect 25222 22480 25228 22492
rect 21131 22452 25228 22480
rect 21131 22449 21143 22452
rect 21085 22443 21143 22449
rect 25222 22440 25228 22452
rect 25280 22440 25286 22492
rect 16114 22412 16120 22424
rect 16075 22384 16120 22412
rect 16114 22372 16120 22384
rect 16172 22372 16178 22424
rect 19720 22412 19748 22440
rect 21729 22415 21787 22421
rect 21729 22412 21741 22415
rect 19720 22384 21741 22412
rect 21729 22381 21741 22384
rect 21775 22412 21787 22415
rect 21775 22384 21956 22412
rect 21775 22381 21787 22384
rect 21729 22375 21787 22381
rect 12805 22347 12863 22353
rect 12805 22313 12817 22347
rect 12851 22344 12863 22347
rect 13814 22344 13820 22356
rect 12851 22316 13820 22344
rect 12851 22313 12863 22316
rect 12805 22307 12863 22313
rect 13814 22304 13820 22316
rect 13872 22344 13878 22356
rect 14093 22347 14151 22353
rect 14093 22344 14105 22347
rect 13872 22316 14105 22344
rect 13872 22304 13878 22316
rect 14093 22313 14105 22316
rect 14139 22313 14151 22347
rect 14093 22307 14151 22313
rect 14185 22347 14243 22353
rect 14185 22313 14197 22347
rect 14231 22313 14243 22347
rect 16298 22344 16304 22356
rect 16259 22316 16304 22344
rect 14185 22307 14243 22313
rect 10689 22279 10747 22285
rect 10689 22245 10701 22279
rect 10735 22276 10747 22279
rect 10781 22279 10839 22285
rect 10781 22276 10793 22279
rect 10735 22248 10793 22276
rect 10735 22245 10747 22248
rect 10689 22239 10747 22245
rect 10781 22245 10793 22248
rect 10827 22276 10839 22279
rect 10870 22276 10876 22288
rect 10827 22248 10876 22276
rect 10827 22245 10839 22248
rect 10781 22239 10839 22245
rect 10870 22236 10876 22248
rect 10928 22236 10934 22288
rect 13630 22236 13636 22288
rect 13688 22276 13694 22288
rect 14200 22276 14228 22307
rect 16298 22304 16304 22316
rect 16356 22304 16362 22356
rect 21928 22353 21956 22384
rect 21913 22347 21971 22353
rect 21913 22313 21925 22347
rect 21959 22313 21971 22347
rect 21913 22307 21971 22313
rect 13688 22248 14228 22276
rect 16568 22279 16626 22285
rect 13688 22236 13694 22248
rect 16568 22245 16580 22279
rect 16614 22276 16626 22279
rect 16850 22276 16856 22288
rect 16614 22248 16856 22276
rect 16614 22245 16626 22248
rect 16568 22239 16626 22245
rect 16850 22236 16856 22248
rect 16908 22236 16914 22288
rect 20622 22236 20628 22288
rect 20680 22276 20686 22288
rect 20901 22279 20959 22285
rect 20901 22276 20913 22279
rect 20680 22248 20913 22276
rect 20680 22236 20686 22248
rect 20901 22245 20913 22248
rect 20947 22276 20959 22279
rect 21361 22279 21419 22285
rect 21361 22276 21373 22279
rect 20947 22248 21373 22276
rect 20947 22245 20959 22248
rect 20901 22239 20959 22245
rect 21361 22245 21373 22248
rect 21407 22245 21419 22279
rect 21361 22239 21419 22245
rect 11048 22211 11106 22217
rect 11048 22177 11060 22211
rect 11094 22208 11106 22211
rect 11330 22208 11336 22220
rect 11094 22180 11336 22208
rect 11094 22177 11106 22180
rect 11048 22171 11106 22177
rect 11330 22168 11336 22180
rect 11388 22168 11394 22220
rect 13173 22211 13231 22217
rect 13173 22177 13185 22211
rect 13219 22208 13231 22211
rect 14001 22211 14059 22217
rect 13219 22180 13952 22208
rect 13219 22177 13231 22180
rect 13173 22171 13231 22177
rect 12158 22140 12164 22152
rect 12119 22112 12164 22140
rect 12158 22100 12164 22112
rect 12216 22100 12222 22152
rect 13633 22143 13691 22149
rect 13633 22109 13645 22143
rect 13679 22140 13691 22143
rect 13722 22140 13728 22152
rect 13679 22112 13728 22140
rect 13679 22109 13691 22112
rect 13633 22103 13691 22109
rect 13722 22100 13728 22112
rect 13780 22100 13786 22152
rect 13924 22140 13952 22180
rect 14001 22177 14013 22211
rect 14047 22208 14059 22211
rect 14182 22208 14188 22220
rect 14047 22180 14188 22208
rect 14047 22177 14059 22180
rect 14001 22171 14059 22177
rect 14182 22168 14188 22180
rect 14240 22208 14246 22220
rect 15013 22211 15071 22217
rect 15013 22208 15025 22211
rect 14240 22180 15025 22208
rect 14240 22168 14246 22180
rect 15013 22177 15025 22180
rect 15059 22177 15071 22211
rect 21928 22208 21956 22307
rect 22002 22236 22008 22288
rect 22060 22276 22066 22288
rect 22169 22279 22227 22285
rect 22169 22276 22181 22279
rect 22060 22248 22181 22276
rect 22060 22236 22066 22248
rect 22169 22245 22181 22248
rect 22215 22245 22227 22279
rect 23658 22276 23664 22288
rect 22169 22239 22227 22245
rect 23216 22248 23664 22276
rect 23216 22208 23244 22248
rect 23658 22236 23664 22248
rect 23716 22276 23722 22288
rect 23845 22279 23903 22285
rect 23845 22276 23857 22279
rect 23716 22248 23857 22276
rect 23716 22236 23722 22248
rect 23845 22245 23857 22248
rect 23891 22245 23903 22279
rect 24578 22276 24584 22288
rect 24539 22248 24584 22276
rect 23845 22239 23903 22245
rect 24578 22236 24584 22248
rect 24636 22276 24642 22288
rect 25133 22279 25191 22285
rect 25133 22276 25145 22279
rect 24636 22248 25145 22276
rect 24636 22236 24642 22248
rect 25133 22245 25145 22248
rect 25179 22245 25191 22279
rect 25133 22239 25191 22245
rect 21928 22180 23244 22208
rect 23308 22180 24256 22208
rect 15013 22171 15071 22177
rect 14090 22140 14096 22152
rect 13924 22112 14096 22140
rect 14090 22100 14096 22112
rect 14148 22100 14154 22152
rect 18230 22140 18236 22152
rect 18191 22112 18236 22140
rect 18230 22100 18236 22112
rect 18288 22100 18294 22152
rect 19797 22143 19855 22149
rect 19797 22109 19809 22143
rect 19843 22140 19855 22143
rect 20162 22140 20168 22152
rect 19843 22112 20168 22140
rect 19843 22109 19855 22112
rect 19797 22103 19855 22109
rect 20162 22100 20168 22112
rect 20220 22100 20226 22152
rect 23308 22149 23336 22180
rect 24228 22152 24256 22180
rect 23293 22143 23351 22149
rect 23293 22109 23305 22143
rect 23339 22109 23351 22143
rect 24210 22140 24216 22152
rect 24171 22112 24216 22140
rect 23293 22103 23351 22109
rect 24210 22100 24216 22112
rect 24268 22100 24274 22152
rect 24670 22100 24676 22152
rect 24728 22140 24734 22152
rect 24765 22143 24823 22149
rect 24765 22140 24777 22143
rect 24728 22112 24777 22140
rect 24728 22100 24734 22112
rect 24765 22109 24777 22112
rect 24811 22109 24823 22143
rect 24765 22103 24823 22109
rect 1104 22050 26864 22072
rect 1104 21998 10315 22050
rect 10367 21998 10379 22050
rect 10431 21998 10443 22050
rect 10495 21998 10507 22050
rect 10559 21998 19648 22050
rect 19700 21998 19712 22050
rect 19764 21998 19776 22050
rect 19828 21998 19840 22050
rect 19892 21998 26864 22050
rect 1104 21976 26864 21998
rect 13630 21896 13636 21948
rect 13688 21936 13694 21948
rect 15013 21939 15071 21945
rect 15013 21936 15025 21939
rect 13688 21908 15025 21936
rect 13688 21896 13694 21908
rect 15013 21905 15025 21908
rect 15059 21905 15071 21939
rect 16298 21936 16304 21948
rect 16259 21908 16304 21936
rect 15013 21899 15071 21905
rect 16298 21896 16304 21908
rect 16356 21896 16362 21948
rect 16761 21939 16819 21945
rect 16761 21905 16773 21939
rect 16807 21936 16819 21939
rect 18230 21936 18236 21948
rect 16807 21908 18236 21936
rect 16807 21905 16819 21908
rect 16761 21899 16819 21905
rect 18230 21896 18236 21908
rect 18288 21896 18294 21948
rect 20162 21936 20168 21948
rect 20123 21908 20168 21936
rect 20162 21896 20168 21908
rect 20220 21896 20226 21948
rect 21726 21936 21732 21948
rect 21687 21908 21732 21936
rect 21726 21896 21732 21908
rect 21784 21896 21790 21948
rect 22646 21936 22652 21948
rect 22607 21908 22652 21936
rect 22646 21896 22652 21908
rect 22704 21896 22710 21948
rect 11146 21868 11152 21880
rect 11107 21840 11152 21868
rect 11146 21828 11152 21840
rect 11204 21828 11210 21880
rect 13900 21871 13958 21877
rect 13900 21837 13912 21871
rect 13946 21868 13958 21871
rect 14090 21868 14096 21880
rect 13946 21840 14096 21868
rect 13946 21837 13958 21840
rect 13900 21831 13958 21837
rect 14090 21828 14096 21840
rect 14148 21828 14154 21880
rect 17313 21871 17371 21877
rect 17313 21837 17325 21871
rect 17359 21868 17371 21871
rect 17678 21868 17684 21880
rect 17359 21840 17684 21868
rect 17359 21837 17371 21840
rect 17313 21831 17371 21837
rect 17678 21828 17684 21840
rect 17736 21828 17742 21880
rect 18046 21800 18052 21812
rect 18007 21772 18052 21800
rect 18046 21760 18052 21772
rect 18104 21760 18110 21812
rect 19705 21803 19763 21809
rect 19705 21769 19717 21803
rect 19751 21800 19763 21803
rect 24029 21803 24087 21809
rect 19751 21772 20484 21800
rect 19751 21769 19763 21772
rect 19705 21763 19763 21769
rect 10502 21692 10508 21744
rect 10560 21732 10566 21744
rect 11241 21735 11299 21741
rect 11241 21732 11253 21735
rect 10560 21704 11253 21732
rect 10560 21692 10566 21704
rect 11241 21701 11253 21704
rect 11287 21701 11299 21735
rect 11241 21695 11299 21701
rect 11330 21692 11336 21744
rect 11388 21732 11394 21744
rect 13630 21732 13636 21744
rect 11388 21704 11433 21732
rect 13591 21704 13636 21732
rect 11388 21692 11394 21704
rect 13630 21692 13636 21704
rect 13688 21692 13694 21744
rect 19334 21692 19340 21744
rect 19392 21732 19398 21744
rect 19518 21732 19524 21744
rect 19392 21704 19524 21732
rect 19392 21692 19398 21704
rect 19518 21692 19524 21704
rect 19576 21732 19582 21744
rect 20456 21741 20484 21772
rect 24029 21769 24041 21803
rect 24075 21800 24087 21803
rect 25222 21800 25228 21812
rect 24075 21772 24440 21800
rect 25183 21772 25228 21800
rect 24075 21769 24087 21772
rect 24029 21763 24087 21769
rect 20257 21735 20315 21741
rect 20257 21732 20269 21735
rect 19576 21704 20269 21732
rect 19576 21692 19582 21704
rect 20257 21701 20269 21704
rect 20303 21701 20315 21735
rect 20257 21695 20315 21701
rect 20441 21735 20499 21741
rect 20441 21701 20453 21735
rect 20487 21732 20499 21735
rect 20530 21732 20536 21744
rect 20487 21704 20536 21732
rect 20487 21701 20499 21704
rect 20441 21695 20499 21701
rect 20530 21692 20536 21704
rect 20588 21692 20594 21744
rect 21358 21692 21364 21744
rect 21416 21732 21422 21744
rect 21821 21735 21879 21741
rect 21821 21732 21833 21735
rect 21416 21704 21833 21732
rect 21416 21692 21422 21704
rect 21821 21701 21833 21704
rect 21867 21701 21879 21735
rect 22002 21732 22008 21744
rect 21963 21704 22008 21732
rect 21821 21695 21879 21701
rect 22002 21692 22008 21704
rect 22060 21692 22066 21744
rect 23474 21692 23480 21744
rect 23532 21732 23538 21744
rect 24121 21735 24179 21741
rect 24121 21732 24133 21735
rect 23532 21704 24133 21732
rect 23532 21692 23538 21704
rect 24121 21701 24133 21704
rect 24167 21701 24179 21735
rect 24121 21695 24179 21701
rect 24210 21692 24216 21744
rect 24268 21732 24274 21744
rect 24268 21704 24313 21732
rect 24268 21692 24274 21704
rect 18230 21664 18236 21676
rect 18191 21636 18236 21664
rect 18230 21624 18236 21636
rect 18288 21624 18294 21676
rect 19797 21667 19855 21673
rect 19797 21633 19809 21667
rect 19843 21664 19855 21667
rect 20622 21664 20628 21676
rect 19843 21636 20628 21664
rect 19843 21633 19855 21636
rect 19797 21627 19855 21633
rect 20622 21624 20628 21636
rect 20680 21624 20686 21676
rect 24026 21624 24032 21676
rect 24084 21664 24090 21676
rect 24412 21664 24440 21772
rect 25222 21760 25228 21772
rect 25280 21760 25286 21812
rect 24084 21636 24440 21664
rect 24084 21624 24090 21636
rect 10594 21596 10600 21608
rect 10555 21568 10600 21596
rect 10594 21556 10600 21568
rect 10652 21556 10658 21608
rect 10686 21556 10692 21608
rect 10744 21596 10750 21608
rect 10781 21599 10839 21605
rect 10781 21596 10793 21599
rect 10744 21568 10793 21596
rect 10744 21556 10750 21568
rect 10781 21565 10793 21568
rect 10827 21565 10839 21599
rect 10781 21559 10839 21565
rect 21361 21599 21419 21605
rect 21361 21565 21373 21599
rect 21407 21596 21419 21599
rect 23474 21596 23480 21608
rect 21407 21568 23480 21596
rect 21407 21565 21419 21568
rect 21361 21559 21419 21565
rect 23474 21556 23480 21568
rect 23532 21556 23538 21608
rect 23658 21596 23664 21608
rect 23619 21568 23664 21596
rect 23658 21556 23664 21568
rect 23716 21556 23722 21608
rect 24854 21556 24860 21608
rect 24912 21596 24918 21608
rect 25409 21599 25467 21605
rect 25409 21596 25421 21599
rect 24912 21568 25421 21596
rect 24912 21556 24918 21568
rect 25409 21565 25421 21568
rect 25455 21565 25467 21599
rect 25409 21559 25467 21565
rect 1104 21506 26864 21528
rect 1104 21454 5648 21506
rect 5700 21454 5712 21506
rect 5764 21454 5776 21506
rect 5828 21454 5840 21506
rect 5892 21454 14982 21506
rect 15034 21454 15046 21506
rect 15098 21454 15110 21506
rect 15162 21454 15174 21506
rect 15226 21454 24315 21506
rect 24367 21454 24379 21506
rect 24431 21454 24443 21506
rect 24495 21454 24507 21506
rect 24559 21454 26864 21506
rect 1104 21432 26864 21454
rect 9122 21352 9128 21404
rect 9180 21392 9186 21404
rect 10502 21392 10508 21404
rect 9180 21364 10508 21392
rect 9180 21352 9186 21364
rect 10502 21352 10508 21364
rect 10560 21352 10566 21404
rect 11330 21352 11336 21404
rect 11388 21392 11394 21404
rect 12069 21395 12127 21401
rect 12069 21392 12081 21395
rect 11388 21364 12081 21392
rect 11388 21352 11394 21364
rect 12069 21361 12081 21364
rect 12115 21361 12127 21395
rect 13630 21392 13636 21404
rect 13591 21364 13636 21392
rect 12069 21355 12127 21361
rect 13630 21352 13636 21364
rect 13688 21392 13694 21404
rect 13814 21392 13820 21404
rect 13688 21364 13820 21392
rect 13688 21352 13694 21364
rect 13814 21352 13820 21364
rect 13872 21352 13878 21404
rect 14090 21392 14096 21404
rect 14051 21364 14096 21392
rect 14090 21352 14096 21364
rect 14148 21352 14154 21404
rect 17497 21395 17555 21401
rect 17497 21361 17509 21395
rect 17543 21392 17555 21395
rect 18046 21392 18052 21404
rect 17543 21364 18052 21392
rect 17543 21361 17555 21364
rect 17497 21355 17555 21361
rect 18046 21352 18052 21364
rect 18104 21352 18110 21404
rect 18138 21352 18144 21404
rect 18196 21392 18202 21404
rect 18196 21364 18241 21392
rect 18196 21352 18202 21364
rect 20162 21352 20168 21404
rect 20220 21392 20226 21404
rect 20257 21395 20315 21401
rect 20257 21392 20269 21395
rect 20220 21364 20269 21392
rect 20220 21352 20226 21364
rect 20257 21361 20269 21364
rect 20303 21361 20315 21395
rect 20714 21392 20720 21404
rect 20675 21364 20720 21392
rect 20257 21355 20315 21361
rect 20714 21352 20720 21364
rect 20772 21352 20778 21404
rect 22002 21352 22008 21404
rect 22060 21392 22066 21404
rect 22281 21395 22339 21401
rect 22281 21392 22293 21395
rect 22060 21364 22293 21392
rect 22060 21352 22066 21364
rect 22281 21361 22293 21364
rect 22327 21361 22339 21395
rect 22281 21355 22339 21361
rect 23293 21395 23351 21401
rect 23293 21361 23305 21395
rect 23339 21392 23351 21395
rect 23474 21392 23480 21404
rect 23339 21364 23480 21392
rect 23339 21361 23351 21364
rect 23293 21355 23351 21361
rect 23474 21352 23480 21364
rect 23532 21352 23538 21404
rect 23937 21395 23995 21401
rect 23937 21361 23949 21395
rect 23983 21392 23995 21395
rect 24026 21392 24032 21404
rect 23983 21364 24032 21392
rect 23983 21361 23995 21364
rect 23937 21355 23995 21361
rect 18156 21256 18184 21352
rect 18325 21259 18383 21265
rect 18325 21256 18337 21259
rect 18156 21228 18337 21256
rect 18325 21225 18337 21228
rect 18371 21225 18383 21259
rect 20732 21256 20760 21352
rect 20901 21259 20959 21265
rect 20901 21256 20913 21259
rect 20732 21228 20913 21256
rect 18325 21219 18383 21225
rect 20901 21225 20913 21228
rect 20947 21225 20959 21259
rect 20901 21219 20959 21225
rect 23385 21259 23443 21265
rect 23385 21225 23397 21259
rect 23431 21256 23443 21259
rect 23952 21256 23980 21355
rect 24026 21352 24032 21364
rect 24084 21352 24090 21404
rect 24210 21392 24216 21404
rect 24171 21364 24216 21392
rect 24210 21352 24216 21364
rect 24268 21352 24274 21404
rect 25222 21392 25228 21404
rect 25183 21364 25228 21392
rect 25222 21352 25228 21364
rect 25280 21352 25286 21404
rect 23431 21228 23980 21256
rect 23431 21225 23443 21228
rect 23385 21219 23443 21225
rect 24210 21216 24216 21268
rect 24268 21256 24274 21268
rect 24670 21256 24676 21268
rect 24268 21228 24676 21256
rect 24268 21216 24274 21228
rect 24670 21216 24676 21228
rect 24728 21216 24734 21268
rect 10229 21191 10287 21197
rect 10229 21157 10241 21191
rect 10275 21188 10287 21191
rect 10689 21191 10747 21197
rect 10689 21188 10701 21191
rect 10275 21160 10701 21188
rect 10275 21157 10287 21160
rect 10229 21151 10287 21157
rect 10689 21157 10701 21160
rect 10735 21188 10747 21191
rect 10778 21188 10784 21200
rect 10735 21160 10784 21188
rect 10735 21157 10747 21160
rect 10689 21151 10747 21157
rect 10778 21148 10784 21160
rect 10836 21148 10842 21200
rect 23658 21148 23664 21200
rect 23716 21188 23722 21200
rect 24397 21191 24455 21197
rect 24397 21188 24409 21191
rect 23716 21160 24409 21188
rect 23716 21148 23722 21160
rect 24397 21157 24409 21160
rect 24443 21188 24455 21191
rect 24857 21191 24915 21197
rect 24857 21188 24869 21191
rect 24443 21160 24869 21188
rect 24443 21157 24455 21160
rect 24397 21151 24455 21157
rect 24857 21157 24869 21160
rect 24903 21157 24915 21191
rect 24857 21151 24915 21157
rect 10594 21080 10600 21132
rect 10652 21120 10658 21132
rect 10934 21123 10992 21129
rect 10934 21120 10946 21123
rect 10652 21092 10946 21120
rect 10652 21080 10658 21092
rect 10934 21089 10946 21092
rect 10980 21089 10992 21123
rect 18570 21123 18628 21129
rect 18570 21120 18582 21123
rect 10934 21083 10992 21089
rect 17788 21092 18582 21120
rect 17788 21064 17816 21092
rect 18570 21089 18582 21092
rect 18616 21089 18628 21123
rect 21146 21123 21204 21129
rect 21146 21120 21158 21123
rect 18570 21083 18628 21089
rect 20180 21092 21158 21120
rect 20180 21064 20208 21092
rect 21146 21089 21158 21092
rect 21192 21089 21204 21123
rect 21146 21083 21204 21089
rect 9674 21052 9680 21064
rect 9635 21024 9680 21052
rect 9674 21012 9680 21024
rect 9732 21012 9738 21064
rect 14185 21055 14243 21061
rect 14185 21021 14197 21055
rect 14231 21052 14243 21055
rect 14550 21052 14556 21064
rect 14231 21024 14556 21052
rect 14231 21021 14243 21024
rect 14185 21015 14243 21021
rect 14550 21012 14556 21024
rect 14608 21012 14614 21064
rect 17770 21052 17776 21064
rect 17731 21024 17776 21052
rect 17770 21012 17776 21024
rect 17828 21012 17834 21064
rect 19705 21055 19763 21061
rect 19705 21021 19717 21055
rect 19751 21052 19763 21055
rect 20162 21052 20168 21064
rect 19751 21024 20168 21052
rect 19751 21021 19763 21024
rect 19705 21015 19763 21021
rect 20162 21012 20168 21024
rect 20220 21012 20226 21064
rect 24581 21055 24639 21061
rect 24581 21021 24593 21055
rect 24627 21052 24639 21055
rect 24670 21052 24676 21064
rect 24627 21024 24676 21052
rect 24627 21021 24639 21024
rect 24581 21015 24639 21021
rect 24670 21012 24676 21024
rect 24728 21012 24734 21064
rect 1104 20962 26864 20984
rect 1104 20910 10315 20962
rect 10367 20910 10379 20962
rect 10431 20910 10443 20962
rect 10495 20910 10507 20962
rect 10559 20910 19648 20962
rect 19700 20910 19712 20962
rect 19764 20910 19776 20962
rect 19828 20910 19840 20962
rect 19892 20910 26864 20962
rect 1104 20888 26864 20910
rect 10321 20851 10379 20857
rect 10321 20817 10333 20851
rect 10367 20848 10379 20851
rect 11330 20848 11336 20860
rect 10367 20820 11336 20848
rect 10367 20817 10379 20820
rect 10321 20811 10379 20817
rect 11330 20808 11336 20820
rect 11388 20808 11394 20860
rect 14182 20848 14188 20860
rect 14143 20820 14188 20848
rect 14182 20808 14188 20820
rect 14240 20808 14246 20860
rect 18506 20848 18512 20860
rect 18467 20820 18512 20848
rect 18506 20808 18512 20820
rect 18564 20808 18570 20860
rect 19518 20848 19524 20860
rect 19479 20820 19524 20848
rect 19518 20808 19524 20820
rect 19576 20808 19582 20860
rect 21358 20848 21364 20860
rect 21319 20820 21364 20848
rect 21358 20808 21364 20820
rect 21416 20808 21422 20860
rect 21726 20848 21732 20860
rect 21687 20820 21732 20848
rect 21726 20808 21732 20820
rect 21784 20808 21790 20860
rect 22002 20808 22008 20860
rect 22060 20848 22066 20860
rect 22097 20851 22155 20857
rect 22097 20848 22109 20851
rect 22060 20820 22109 20848
rect 22060 20808 22066 20820
rect 22097 20817 22109 20820
rect 22143 20817 22155 20851
rect 22097 20811 22155 20817
rect 23934 20808 23940 20860
rect 23992 20848 23998 20860
rect 24673 20851 24731 20857
rect 24673 20848 24685 20851
rect 23992 20820 24685 20848
rect 23992 20808 23998 20820
rect 24673 20817 24685 20820
rect 24719 20848 24731 20851
rect 25130 20848 25136 20860
rect 24719 20820 25136 20848
rect 24719 20817 24731 20820
rect 24673 20811 24731 20817
rect 25130 20808 25136 20820
rect 25188 20808 25194 20860
rect 11054 20740 11060 20792
rect 11112 20780 11118 20792
rect 12158 20780 12164 20792
rect 11112 20752 12164 20780
rect 11112 20740 11118 20752
rect 9674 20672 9680 20724
rect 9732 20712 9738 20724
rect 11149 20715 11207 20721
rect 11149 20712 11161 20715
rect 9732 20684 11161 20712
rect 9732 20672 9738 20684
rect 11149 20681 11161 20684
rect 11195 20681 11207 20715
rect 11149 20675 11207 20681
rect 10134 20604 10140 20656
rect 10192 20644 10198 20656
rect 10686 20644 10692 20656
rect 10192 20616 10692 20644
rect 10192 20604 10198 20616
rect 10686 20604 10692 20616
rect 10744 20644 10750 20656
rect 11348 20653 11376 20752
rect 12158 20740 12164 20752
rect 12216 20740 12222 20792
rect 12434 20672 12440 20724
rect 12492 20712 12498 20724
rect 14550 20712 14556 20724
rect 12492 20684 12537 20712
rect 14511 20684 14556 20712
rect 12492 20672 12498 20684
rect 14550 20672 14556 20684
rect 14608 20672 14614 20724
rect 16758 20712 16764 20724
rect 16719 20684 16764 20712
rect 16758 20672 16764 20684
rect 16816 20672 16822 20724
rect 18414 20712 18420 20724
rect 18375 20684 18420 20712
rect 18414 20672 18420 20684
rect 18472 20672 18478 20724
rect 19978 20712 19984 20724
rect 19939 20684 19984 20712
rect 19978 20672 19984 20684
rect 20036 20672 20042 20724
rect 24946 20712 24952 20724
rect 24780 20684 24952 20712
rect 11241 20647 11299 20653
rect 11241 20644 11253 20647
rect 10744 20616 11253 20644
rect 10744 20604 10750 20616
rect 11241 20613 11253 20616
rect 11287 20613 11299 20647
rect 11241 20607 11299 20613
rect 11333 20647 11391 20653
rect 11333 20613 11345 20647
rect 11379 20613 11391 20647
rect 14642 20644 14648 20656
rect 14603 20616 14648 20644
rect 11333 20607 11391 20613
rect 14642 20604 14648 20616
rect 14700 20604 14706 20656
rect 14737 20647 14795 20653
rect 14737 20613 14749 20647
rect 14783 20613 14795 20647
rect 14737 20607 14795 20613
rect 10781 20579 10839 20585
rect 10781 20545 10793 20579
rect 10827 20576 10839 20579
rect 12434 20576 12440 20588
rect 10827 20548 12440 20576
rect 10827 20545 10839 20548
rect 10781 20539 10839 20545
rect 12434 20536 12440 20548
rect 12492 20536 12498 20588
rect 12618 20576 12624 20588
rect 12579 20548 12624 20576
rect 12618 20536 12624 20548
rect 12676 20536 12682 20588
rect 14090 20536 14096 20588
rect 14148 20576 14154 20588
rect 14752 20576 14780 20607
rect 16022 20604 16028 20656
rect 16080 20644 16086 20656
rect 16853 20647 16911 20653
rect 16853 20644 16865 20647
rect 16080 20616 16865 20644
rect 16080 20604 16086 20616
rect 16853 20613 16865 20616
rect 16899 20613 16911 20647
rect 16853 20607 16911 20613
rect 17037 20647 17095 20653
rect 17037 20613 17049 20647
rect 17083 20613 17095 20647
rect 17037 20607 17095 20613
rect 14148 20548 14780 20576
rect 14148 20536 14154 20548
rect 10689 20511 10747 20517
rect 10689 20477 10701 20511
rect 10735 20508 10747 20511
rect 11146 20508 11152 20520
rect 10735 20480 11152 20508
rect 10735 20477 10747 20480
rect 10689 20471 10747 20477
rect 11146 20468 11152 20480
rect 11204 20468 11210 20520
rect 16206 20508 16212 20520
rect 16167 20480 16212 20508
rect 16206 20468 16212 20480
rect 16264 20468 16270 20520
rect 16393 20511 16451 20517
rect 16393 20477 16405 20511
rect 16439 20508 16451 20511
rect 16666 20508 16672 20520
rect 16439 20480 16672 20508
rect 16439 20477 16451 20480
rect 16393 20471 16451 20477
rect 16666 20468 16672 20480
rect 16724 20468 16730 20520
rect 16850 20468 16856 20520
rect 16908 20508 16914 20520
rect 17052 20508 17080 20607
rect 17770 20604 17776 20656
rect 17828 20644 17834 20656
rect 18601 20647 18659 20653
rect 18601 20644 18613 20647
rect 17828 20616 18613 20644
rect 17828 20604 17834 20616
rect 18601 20613 18613 20616
rect 18647 20613 18659 20647
rect 18601 20607 18659 20613
rect 20073 20647 20131 20653
rect 20073 20613 20085 20647
rect 20119 20613 20131 20647
rect 20073 20607 20131 20613
rect 18049 20579 18107 20585
rect 18049 20545 18061 20579
rect 18095 20576 18107 20579
rect 20088 20576 20116 20607
rect 20162 20604 20168 20656
rect 20220 20644 20226 20656
rect 20901 20647 20959 20653
rect 20901 20644 20913 20647
rect 20220 20616 20913 20644
rect 20220 20604 20226 20616
rect 20901 20613 20913 20616
rect 20947 20613 20959 20647
rect 20901 20607 20959 20613
rect 24026 20604 24032 20656
rect 24084 20644 24090 20656
rect 24780 20653 24808 20684
rect 24946 20672 24952 20684
rect 25004 20672 25010 20724
rect 25314 20712 25320 20724
rect 25275 20684 25320 20712
rect 25314 20672 25320 20684
rect 25372 20672 25378 20724
rect 24765 20647 24823 20653
rect 24765 20644 24777 20647
rect 24084 20616 24777 20644
rect 24084 20604 24090 20616
rect 24765 20613 24777 20616
rect 24811 20613 24823 20647
rect 24765 20607 24823 20613
rect 24854 20604 24860 20656
rect 24912 20644 24918 20656
rect 24912 20616 24957 20644
rect 24912 20604 24918 20616
rect 20254 20576 20260 20588
rect 18095 20548 20260 20576
rect 18095 20545 18107 20548
rect 18049 20539 18107 20545
rect 20254 20536 20260 20548
rect 20312 20536 20318 20588
rect 19153 20511 19211 20517
rect 19153 20508 19165 20511
rect 16908 20480 19165 20508
rect 16908 20468 16914 20480
rect 19153 20477 19165 20480
rect 19199 20508 19211 20511
rect 19242 20508 19248 20520
rect 19199 20480 19248 20508
rect 19199 20477 19211 20480
rect 19153 20471 19211 20477
rect 19242 20468 19248 20480
rect 19300 20468 19306 20520
rect 19613 20511 19671 20517
rect 19613 20477 19625 20511
rect 19659 20508 19671 20511
rect 20714 20508 20720 20520
rect 19659 20480 20720 20508
rect 19659 20477 19671 20480
rect 19613 20471 19671 20477
rect 20714 20468 20720 20480
rect 20772 20468 20778 20520
rect 23934 20468 23940 20520
rect 23992 20508 23998 20520
rect 24305 20511 24363 20517
rect 24305 20508 24317 20511
rect 23992 20480 24317 20508
rect 23992 20468 23998 20480
rect 24305 20477 24317 20480
rect 24351 20477 24363 20511
rect 24305 20471 24363 20477
rect 1104 20418 26864 20440
rect 1104 20366 5648 20418
rect 5700 20366 5712 20418
rect 5764 20366 5776 20418
rect 5828 20366 5840 20418
rect 5892 20366 14982 20418
rect 15034 20366 15046 20418
rect 15098 20366 15110 20418
rect 15162 20366 15174 20418
rect 15226 20366 24315 20418
rect 24367 20366 24379 20418
rect 24431 20366 24443 20418
rect 24495 20366 24507 20418
rect 24559 20366 26864 20418
rect 1104 20344 26864 20366
rect 9674 20264 9680 20316
rect 9732 20304 9738 20316
rect 10413 20307 10471 20313
rect 10413 20304 10425 20307
rect 9732 20276 10425 20304
rect 9732 20264 9738 20276
rect 10413 20273 10425 20276
rect 10459 20273 10471 20307
rect 10413 20267 10471 20273
rect 12434 20264 12440 20316
rect 12492 20304 12498 20316
rect 13357 20307 13415 20313
rect 13357 20304 13369 20307
rect 12492 20276 13369 20304
rect 12492 20264 12498 20276
rect 13357 20273 13369 20276
rect 13403 20273 13415 20307
rect 14090 20304 14096 20316
rect 14051 20276 14096 20304
rect 13357 20267 13415 20273
rect 14090 20264 14096 20276
rect 14148 20264 14154 20316
rect 14550 20264 14556 20316
rect 14608 20304 14614 20316
rect 15013 20307 15071 20313
rect 15013 20304 15025 20307
rect 14608 20276 15025 20304
rect 14608 20264 14614 20276
rect 15013 20273 15025 20276
rect 15059 20273 15071 20307
rect 16022 20304 16028 20316
rect 15983 20276 16028 20304
rect 15013 20267 15071 20273
rect 16022 20264 16028 20276
rect 16080 20264 16086 20316
rect 18233 20307 18291 20313
rect 18233 20273 18245 20307
rect 18279 20304 18291 20307
rect 18506 20304 18512 20316
rect 18279 20276 18512 20304
rect 18279 20273 18291 20276
rect 18233 20267 18291 20273
rect 18506 20264 18512 20276
rect 18564 20264 18570 20316
rect 19794 20304 19800 20316
rect 19168 20276 19800 20304
rect 10134 20236 10140 20248
rect 10095 20208 10140 20236
rect 10134 20196 10140 20208
rect 10192 20196 10198 20248
rect 14642 20236 14648 20248
rect 14603 20208 14648 20236
rect 14642 20196 14648 20208
rect 14700 20196 14706 20248
rect 10042 20128 10048 20180
rect 10100 20168 10106 20180
rect 10781 20171 10839 20177
rect 10781 20168 10793 20171
rect 10100 20140 10793 20168
rect 10100 20128 10106 20140
rect 10781 20137 10793 20140
rect 10827 20168 10839 20171
rect 10962 20168 10968 20180
rect 10827 20140 10968 20168
rect 10827 20137 10839 20140
rect 10781 20131 10839 20137
rect 10962 20128 10968 20140
rect 11020 20128 11026 20180
rect 18414 20128 18420 20180
rect 18472 20168 18478 20180
rect 19168 20177 19196 20276
rect 19794 20264 19800 20276
rect 19852 20264 19858 20316
rect 19978 20264 19984 20316
rect 20036 20304 20042 20316
rect 20073 20307 20131 20313
rect 20073 20304 20085 20307
rect 20036 20276 20085 20304
rect 20036 20264 20042 20276
rect 20073 20273 20085 20276
rect 20119 20273 20131 20307
rect 20073 20267 20131 20273
rect 20162 20264 20168 20316
rect 20220 20304 20226 20316
rect 20441 20307 20499 20313
rect 20441 20304 20453 20307
rect 20220 20276 20453 20304
rect 20220 20264 20226 20276
rect 20441 20273 20453 20276
rect 20487 20273 20499 20307
rect 20441 20267 20499 20273
rect 24026 20264 24032 20316
rect 24084 20304 24090 20316
rect 24673 20307 24731 20313
rect 24673 20304 24685 20307
rect 24084 20276 24685 20304
rect 24084 20264 24090 20276
rect 24673 20273 24685 20276
rect 24719 20273 24731 20307
rect 25130 20304 25136 20316
rect 25091 20276 25136 20304
rect 24673 20267 24731 20273
rect 25130 20264 25136 20276
rect 25188 20264 25194 20316
rect 18601 20171 18659 20177
rect 18601 20168 18613 20171
rect 18472 20140 18613 20168
rect 18472 20128 18478 20140
rect 18601 20137 18613 20140
rect 18647 20168 18659 20171
rect 19153 20171 19211 20177
rect 19153 20168 19165 20171
rect 18647 20140 19165 20168
rect 18647 20137 18659 20140
rect 18601 20131 18659 20137
rect 19153 20137 19165 20140
rect 19199 20137 19211 20171
rect 19153 20131 19211 20137
rect 19242 20128 19248 20180
rect 19300 20168 19306 20180
rect 19300 20140 19345 20168
rect 19300 20128 19306 20140
rect 22646 20128 22652 20180
rect 22704 20168 22710 20180
rect 23201 20171 23259 20177
rect 23201 20168 23213 20171
rect 22704 20140 23213 20168
rect 22704 20128 22710 20140
rect 23201 20137 23213 20140
rect 23247 20168 23259 20171
rect 24302 20168 24308 20180
rect 23247 20140 24164 20168
rect 24263 20140 24308 20168
rect 23247 20137 23259 20140
rect 23201 20131 23259 20137
rect 10870 20060 10876 20112
rect 10928 20100 10934 20112
rect 11333 20103 11391 20109
rect 11333 20100 11345 20103
rect 10928 20072 11345 20100
rect 10928 20060 10934 20072
rect 11333 20069 11345 20072
rect 11379 20100 11391 20103
rect 11425 20103 11483 20109
rect 11425 20100 11437 20103
rect 11379 20072 11437 20100
rect 11379 20069 11391 20072
rect 11333 20063 11391 20069
rect 11425 20069 11437 20072
rect 11471 20100 11483 20103
rect 12250 20100 12256 20112
rect 11471 20072 12256 20100
rect 11471 20069 11483 20072
rect 11425 20063 11483 20069
rect 12250 20060 12256 20072
rect 12308 20060 12314 20112
rect 14458 20060 14464 20112
rect 14516 20100 14522 20112
rect 16206 20100 16212 20112
rect 14516 20072 16212 20100
rect 14516 20060 14522 20072
rect 16206 20060 16212 20072
rect 16264 20060 16270 20112
rect 19058 20100 19064 20112
rect 19019 20072 19064 20100
rect 19058 20060 19064 20072
rect 19116 20060 19122 20112
rect 20714 20060 20720 20112
rect 20772 20100 20778 20112
rect 20901 20103 20959 20109
rect 20901 20100 20913 20103
rect 20772 20072 20913 20100
rect 20772 20060 20778 20072
rect 20901 20069 20913 20072
rect 20947 20100 20959 20103
rect 21361 20103 21419 20109
rect 21361 20100 21373 20103
rect 20947 20072 21373 20100
rect 20947 20069 20959 20072
rect 20901 20063 20959 20069
rect 21361 20069 21373 20072
rect 21407 20069 21419 20103
rect 24136 20100 24164 20140
rect 24302 20128 24308 20140
rect 24360 20128 24366 20180
rect 25225 20103 25283 20109
rect 24136 20072 24256 20100
rect 21361 20063 21419 20069
rect 11692 20035 11750 20041
rect 11692 20001 11704 20035
rect 11738 20032 11750 20035
rect 11790 20032 11796 20044
rect 11738 20004 11796 20032
rect 11738 20001 11750 20004
rect 11692 19995 11750 20001
rect 11790 19992 11796 20004
rect 11848 19992 11854 20044
rect 15749 20035 15807 20041
rect 15749 20001 15761 20035
rect 15795 20032 15807 20035
rect 15838 20032 15844 20044
rect 15795 20004 15844 20032
rect 15795 20001 15807 20004
rect 15749 19995 15807 20001
rect 15838 19992 15844 20004
rect 15896 20032 15902 20044
rect 16454 20035 16512 20041
rect 16454 20032 16466 20035
rect 15896 20004 16466 20032
rect 15896 19992 15902 20004
rect 16454 20001 16466 20004
rect 16500 20001 16512 20035
rect 23474 20032 23480 20044
rect 23435 20004 23480 20032
rect 16454 19995 16512 20001
rect 23474 19992 23480 20004
rect 23532 20032 23538 20044
rect 24121 20035 24179 20041
rect 24121 20032 24133 20035
rect 23532 20004 24133 20032
rect 23532 19992 23538 20004
rect 24121 20001 24133 20004
rect 24167 20001 24179 20035
rect 24121 19995 24179 20001
rect 24228 20032 24256 20072
rect 25225 20069 25237 20103
rect 25271 20100 25283 20103
rect 25314 20100 25320 20112
rect 25271 20072 25320 20100
rect 25271 20069 25283 20072
rect 25225 20063 25283 20069
rect 25314 20060 25320 20072
rect 25372 20060 25378 20112
rect 25498 20032 25504 20044
rect 24228 20004 25504 20032
rect 12802 19964 12808 19976
rect 12763 19936 12808 19964
rect 12802 19924 12808 19936
rect 12860 19924 12866 19976
rect 14182 19964 14188 19976
rect 14143 19936 14188 19964
rect 14182 19924 14188 19936
rect 14240 19924 14246 19976
rect 17589 19967 17647 19973
rect 17589 19933 17601 19967
rect 17635 19964 17647 19967
rect 17770 19964 17776 19976
rect 17635 19936 17776 19964
rect 17635 19933 17647 19936
rect 17589 19927 17647 19933
rect 17770 19924 17776 19936
rect 17828 19924 17834 19976
rect 18690 19964 18696 19976
rect 18651 19936 18696 19964
rect 18690 19924 18696 19936
rect 18748 19924 18754 19976
rect 21082 19964 21088 19976
rect 21043 19936 21088 19964
rect 21082 19924 21088 19936
rect 21140 19924 21146 19976
rect 22649 19967 22707 19973
rect 22649 19933 22661 19967
rect 22695 19964 22707 19967
rect 23382 19964 23388 19976
rect 22695 19936 23388 19964
rect 22695 19933 22707 19936
rect 22649 19927 22707 19933
rect 23382 19924 23388 19936
rect 23440 19924 23446 19976
rect 23658 19964 23664 19976
rect 23619 19936 23664 19964
rect 23658 19924 23664 19936
rect 23716 19924 23722 19976
rect 24029 19967 24087 19973
rect 24029 19933 24041 19967
rect 24075 19964 24087 19967
rect 24228 19964 24256 20004
rect 25498 19992 25504 20004
rect 25556 19992 25562 20044
rect 25406 19964 25412 19976
rect 24075 19936 24256 19964
rect 25367 19936 25412 19964
rect 24075 19933 24087 19936
rect 24029 19927 24087 19933
rect 25406 19924 25412 19936
rect 25464 19924 25470 19976
rect 25774 19964 25780 19976
rect 25735 19936 25780 19964
rect 25774 19924 25780 19936
rect 25832 19924 25838 19976
rect 1104 19874 26864 19896
rect 1104 19822 10315 19874
rect 10367 19822 10379 19874
rect 10431 19822 10443 19874
rect 10495 19822 10507 19874
rect 10559 19822 19648 19874
rect 19700 19822 19712 19874
rect 19764 19822 19776 19874
rect 19828 19822 19840 19874
rect 19892 19822 26864 19874
rect 1104 19800 26864 19822
rect 11238 19760 11244 19772
rect 11199 19732 11244 19760
rect 11238 19720 11244 19732
rect 11296 19720 11302 19772
rect 13630 19760 13636 19772
rect 13591 19732 13636 19760
rect 13630 19720 13636 19732
rect 13688 19720 13694 19772
rect 13722 19720 13728 19772
rect 13780 19760 13786 19772
rect 13909 19763 13967 19769
rect 13909 19760 13921 19763
rect 13780 19732 13921 19760
rect 13780 19720 13786 19732
rect 13909 19729 13921 19732
rect 13955 19729 13967 19763
rect 15838 19760 15844 19772
rect 15799 19732 15844 19760
rect 13909 19723 13967 19729
rect 15838 19720 15844 19732
rect 15896 19720 15902 19772
rect 16390 19760 16396 19772
rect 16351 19732 16396 19760
rect 16390 19720 16396 19732
rect 16448 19720 16454 19772
rect 16850 19760 16856 19772
rect 16811 19732 16856 19760
rect 16850 19720 16856 19732
rect 16908 19720 16914 19772
rect 17770 19760 17776 19772
rect 17731 19732 17776 19760
rect 17770 19720 17776 19732
rect 17828 19720 17834 19772
rect 18417 19763 18475 19769
rect 18417 19729 18429 19763
rect 18463 19760 18475 19763
rect 18690 19760 18696 19772
rect 18463 19732 18696 19760
rect 18463 19729 18475 19732
rect 18417 19723 18475 19729
rect 18690 19720 18696 19732
rect 18748 19760 18754 19772
rect 19429 19763 19487 19769
rect 19429 19760 19441 19763
rect 18748 19732 19441 19760
rect 18748 19720 18754 19732
rect 19429 19729 19441 19732
rect 19475 19729 19487 19763
rect 19429 19723 19487 19729
rect 19613 19763 19671 19769
rect 19613 19729 19625 19763
rect 19659 19760 19671 19763
rect 19978 19760 19984 19772
rect 19659 19732 19984 19760
rect 19659 19729 19671 19732
rect 19613 19723 19671 19729
rect 19978 19720 19984 19732
rect 20036 19720 20042 19772
rect 20165 19763 20223 19769
rect 20165 19729 20177 19763
rect 20211 19760 20223 19763
rect 20254 19760 20260 19772
rect 20211 19732 20260 19760
rect 20211 19729 20223 19732
rect 20165 19723 20223 19729
rect 20254 19720 20260 19732
rect 20312 19720 20318 19772
rect 11146 19692 11152 19704
rect 11107 19664 11152 19692
rect 11146 19652 11152 19664
rect 11204 19652 11210 19704
rect 13449 19627 13507 19633
rect 13449 19593 13461 19627
rect 13495 19624 13507 19627
rect 13740 19624 13768 19720
rect 19058 19692 19064 19704
rect 19019 19664 19064 19692
rect 19058 19652 19064 19664
rect 19116 19652 19122 19704
rect 21100 19664 21588 19692
rect 13495 19596 13768 19624
rect 13495 19593 13507 19596
rect 13449 19587 13507 19593
rect 14090 19584 14096 19636
rect 14148 19624 14154 19636
rect 14717 19627 14775 19633
rect 14717 19624 14729 19627
rect 14148 19596 14729 19624
rect 14148 19584 14154 19596
rect 14717 19593 14729 19596
rect 14763 19593 14775 19627
rect 14717 19587 14775 19593
rect 11425 19559 11483 19565
rect 11425 19525 11437 19559
rect 11471 19556 11483 19559
rect 11471 19528 11836 19556
rect 11471 19525 11483 19528
rect 11425 19519 11483 19525
rect 11808 19432 11836 19528
rect 12342 19516 12348 19568
rect 12400 19556 12406 19568
rect 12437 19559 12495 19565
rect 12437 19556 12449 19559
rect 12400 19528 12449 19556
rect 12400 19516 12406 19528
rect 12437 19525 12449 19528
rect 12483 19525 12495 19559
rect 12437 19519 12495 19525
rect 13814 19516 13820 19568
rect 13872 19556 13878 19568
rect 14458 19556 14464 19568
rect 13872 19528 14464 19556
rect 13872 19516 13878 19528
rect 14458 19516 14464 19528
rect 14516 19516 14522 19568
rect 17954 19516 17960 19568
rect 18012 19556 18018 19568
rect 18509 19559 18567 19565
rect 18509 19556 18521 19559
rect 18012 19528 18521 19556
rect 18012 19516 18018 19528
rect 18509 19525 18521 19528
rect 18555 19525 18567 19559
rect 18509 19519 18567 19525
rect 18601 19559 18659 19565
rect 18601 19525 18613 19559
rect 18647 19525 18659 19559
rect 18601 19519 18659 19525
rect 18616 19488 18644 19519
rect 20898 19516 20904 19568
rect 20956 19556 20962 19568
rect 21100 19565 21128 19664
rect 21358 19633 21364 19636
rect 21352 19587 21364 19633
rect 21416 19624 21422 19636
rect 21560 19624 21588 19664
rect 24026 19624 24032 19636
rect 21416 19596 21452 19624
rect 21560 19596 24032 19624
rect 21358 19584 21364 19587
rect 21416 19584 21422 19596
rect 24026 19584 24032 19596
rect 24084 19584 24090 19636
rect 24302 19633 24308 19636
rect 24296 19624 24308 19633
rect 24136 19596 24308 19624
rect 21085 19559 21143 19565
rect 21085 19556 21097 19559
rect 20956 19528 21097 19556
rect 20956 19516 20962 19528
rect 21085 19525 21097 19528
rect 21131 19525 21143 19559
rect 21085 19519 21143 19525
rect 23566 19516 23572 19568
rect 23624 19556 23630 19568
rect 23937 19559 23995 19565
rect 23937 19556 23949 19559
rect 23624 19528 23949 19556
rect 23624 19516 23630 19528
rect 23937 19525 23949 19528
rect 23983 19556 23995 19559
rect 24136 19556 24164 19596
rect 24296 19587 24308 19596
rect 24360 19624 24366 19636
rect 24854 19624 24860 19636
rect 24360 19596 24860 19624
rect 24302 19584 24308 19587
rect 24360 19584 24366 19596
rect 24854 19584 24860 19596
rect 24912 19624 24918 19636
rect 25774 19624 25780 19636
rect 24912 19596 25780 19624
rect 24912 19584 24918 19596
rect 25774 19584 25780 19596
rect 25832 19584 25838 19636
rect 23983 19528 24164 19556
rect 23983 19525 23995 19528
rect 23937 19519 23995 19525
rect 17420 19460 18644 19488
rect 10781 19423 10839 19429
rect 10781 19389 10793 19423
rect 10827 19420 10839 19423
rect 11054 19420 11060 19432
rect 10827 19392 11060 19420
rect 10827 19389 10839 19392
rect 10781 19383 10839 19389
rect 11054 19380 11060 19392
rect 11112 19380 11118 19432
rect 11790 19420 11796 19432
rect 11751 19392 11796 19420
rect 11790 19380 11796 19392
rect 11848 19380 11854 19432
rect 17310 19380 17316 19432
rect 17368 19420 17374 19432
rect 17420 19429 17448 19460
rect 17405 19423 17463 19429
rect 17405 19420 17417 19423
rect 17368 19392 17417 19420
rect 17368 19380 17374 19392
rect 17405 19389 17417 19392
rect 17451 19389 17463 19423
rect 18046 19420 18052 19432
rect 18007 19392 18052 19420
rect 17405 19383 17463 19389
rect 18046 19380 18052 19392
rect 18104 19380 18110 19432
rect 20990 19420 20996 19432
rect 20951 19392 20996 19420
rect 20990 19380 20996 19392
rect 21048 19420 21054 19432
rect 22465 19423 22523 19429
rect 22465 19420 22477 19423
rect 21048 19392 22477 19420
rect 21048 19380 21054 19392
rect 22465 19389 22477 19392
rect 22511 19420 22523 19423
rect 22554 19420 22560 19432
rect 22511 19392 22560 19420
rect 22511 19389 22523 19392
rect 22465 19383 22523 19389
rect 22554 19380 22560 19392
rect 22612 19380 22618 19432
rect 25409 19423 25467 19429
rect 25409 19389 25421 19423
rect 25455 19420 25467 19423
rect 25498 19420 25504 19432
rect 25455 19392 25504 19420
rect 25455 19389 25467 19392
rect 25409 19383 25467 19389
rect 25498 19380 25504 19392
rect 25556 19380 25562 19432
rect 1104 19330 26864 19352
rect 1104 19278 5648 19330
rect 5700 19278 5712 19330
rect 5764 19278 5776 19330
rect 5828 19278 5840 19330
rect 5892 19278 14982 19330
rect 15034 19278 15046 19330
rect 15098 19278 15110 19330
rect 15162 19278 15174 19330
rect 15226 19278 24315 19330
rect 24367 19278 24379 19330
rect 24431 19278 24443 19330
rect 24495 19278 24507 19330
rect 24559 19278 26864 19330
rect 1104 19256 26864 19278
rect 14458 19176 14464 19228
rect 14516 19216 14522 19228
rect 14645 19219 14703 19225
rect 14645 19216 14657 19219
rect 14516 19188 14657 19216
rect 14516 19176 14522 19188
rect 14645 19185 14657 19188
rect 14691 19185 14703 19219
rect 14645 19179 14703 19185
rect 22094 19176 22100 19228
rect 22152 19216 22158 19228
rect 23290 19216 23296 19228
rect 22152 19188 23296 19216
rect 22152 19176 22158 19188
rect 23290 19176 23296 19188
rect 23348 19176 23354 19228
rect 23477 19219 23535 19225
rect 23477 19185 23489 19219
rect 23523 19216 23535 19219
rect 23566 19216 23572 19228
rect 23523 19188 23572 19216
rect 23523 19185 23535 19188
rect 23477 19179 23535 19185
rect 23566 19176 23572 19188
rect 23624 19176 23630 19228
rect 24026 19176 24032 19228
rect 24084 19216 24090 19228
rect 24581 19219 24639 19225
rect 24581 19216 24593 19219
rect 24084 19188 24593 19216
rect 24084 19176 24090 19188
rect 24581 19185 24593 19188
rect 24627 19185 24639 19219
rect 24581 19179 24639 19185
rect 24486 19108 24492 19160
rect 24544 19148 24550 19160
rect 25866 19148 25872 19160
rect 24544 19120 25872 19148
rect 24544 19108 24550 19120
rect 25866 19108 25872 19120
rect 25924 19108 25930 19160
rect 11238 19080 11244 19092
rect 10980 19052 11244 19080
rect 10873 19015 10931 19021
rect 10873 18981 10885 19015
rect 10919 19012 10931 19015
rect 10980 19012 11008 19052
rect 11238 19040 11244 19052
rect 11296 19040 11302 19092
rect 11793 19083 11851 19089
rect 11793 19049 11805 19083
rect 11839 19080 11851 19083
rect 15930 19080 15936 19092
rect 11839 19052 12848 19080
rect 15891 19052 15936 19080
rect 11839 19049 11851 19052
rect 11793 19043 11851 19049
rect 12820 19024 12848 19052
rect 15930 19040 15936 19052
rect 15988 19040 15994 19092
rect 17310 19040 17316 19092
rect 17368 19080 17374 19092
rect 18141 19083 18199 19089
rect 18141 19080 18153 19083
rect 17368 19052 18153 19080
rect 17368 19040 17374 19052
rect 18141 19049 18153 19052
rect 18187 19049 18199 19083
rect 18141 19043 18199 19049
rect 19797 19083 19855 19089
rect 19797 19049 19809 19083
rect 19843 19049 19855 19083
rect 19797 19043 19855 19049
rect 10919 18984 11008 19012
rect 10919 18981 10931 18984
rect 10873 18975 10931 18981
rect 11054 18972 11060 19024
rect 11112 19012 11118 19024
rect 11609 19015 11667 19021
rect 11609 19012 11621 19015
rect 11112 18984 11621 19012
rect 11112 18972 11118 18984
rect 11609 18981 11621 18984
rect 11655 19012 11667 19015
rect 12161 19015 12219 19021
rect 12161 19012 12173 19015
rect 11655 18984 12173 19012
rect 11655 18981 11667 18984
rect 11609 18975 11667 18981
rect 12161 18981 12173 18984
rect 12207 18981 12219 19015
rect 12161 18975 12219 18981
rect 12250 18972 12256 19024
rect 12308 19012 12314 19024
rect 12713 19015 12771 19021
rect 12713 19012 12725 19015
rect 12308 18984 12725 19012
rect 12308 18972 12314 18984
rect 12713 18981 12725 18984
rect 12759 18981 12771 19015
rect 12713 18975 12771 18981
rect 10505 18947 10563 18953
rect 10505 18913 10517 18947
rect 10551 18944 10563 18947
rect 10962 18944 10968 18956
rect 10551 18916 10968 18944
rect 10551 18913 10563 18916
rect 10505 18907 10563 18913
rect 10962 18904 10968 18916
rect 11020 18904 11026 18956
rect 11238 18904 11244 18956
rect 11296 18944 11302 18956
rect 11517 18947 11575 18953
rect 11517 18944 11529 18947
rect 11296 18916 11529 18944
rect 11296 18904 11302 18916
rect 11517 18913 11529 18916
rect 11563 18944 11575 18947
rect 12342 18944 12348 18956
rect 11563 18916 12348 18944
rect 11563 18913 11575 18916
rect 11517 18907 11575 18913
rect 12342 18904 12348 18916
rect 12400 18904 12406 18956
rect 12621 18947 12679 18953
rect 12621 18913 12633 18947
rect 12667 18944 12679 18947
rect 12728 18944 12756 18975
rect 12802 18972 12808 19024
rect 12860 19012 12866 19024
rect 12969 19015 13027 19021
rect 12969 19012 12981 19015
rect 12860 18984 12981 19012
rect 12860 18972 12866 18984
rect 12969 18981 12981 18984
rect 13015 18981 13027 19015
rect 16666 19012 16672 19024
rect 16627 18984 16672 19012
rect 12969 18975 13027 18981
rect 16666 18972 16672 18984
rect 16724 19012 16730 19024
rect 17862 19012 17868 19024
rect 16724 18984 17868 19012
rect 16724 18972 16730 18984
rect 17862 18972 17868 18984
rect 17920 18972 17926 19024
rect 18785 19015 18843 19021
rect 18785 18981 18797 19015
rect 18831 19012 18843 19015
rect 19518 19012 19524 19024
rect 18831 18984 19524 19012
rect 18831 18981 18843 18984
rect 18785 18975 18843 18981
rect 19518 18972 19524 18984
rect 19576 19012 19582 19024
rect 19812 19012 19840 19043
rect 23658 19040 23664 19092
rect 23716 19080 23722 19092
rect 24029 19083 24087 19089
rect 24029 19080 24041 19083
rect 23716 19052 24041 19080
rect 23716 19040 23722 19052
rect 24029 19049 24041 19052
rect 24075 19049 24087 19083
rect 24029 19043 24087 19049
rect 24213 19083 24271 19089
rect 24213 19049 24225 19083
rect 24259 19080 24271 19083
rect 24302 19080 24308 19092
rect 24259 19052 24308 19080
rect 24259 19049 24271 19052
rect 24213 19043 24271 19049
rect 20898 19012 20904 19024
rect 19576 18984 19840 19012
rect 20811 18984 20904 19012
rect 19576 18972 19582 18984
rect 20898 18972 20904 18984
rect 20956 18972 20962 19024
rect 20990 18972 20996 19024
rect 21048 19012 21054 19024
rect 21157 19015 21215 19021
rect 21157 19012 21169 19015
rect 21048 18984 21169 19012
rect 21048 18972 21054 18984
rect 21157 18981 21169 18984
rect 21203 18981 21215 19015
rect 23934 19012 23940 19024
rect 23895 18984 23940 19012
rect 21157 18975 21215 18981
rect 23934 18972 23940 18984
rect 23992 18972 23998 19024
rect 24044 19012 24072 19043
rect 24302 19040 24308 19052
rect 24360 19040 24366 19092
rect 24949 19015 25007 19021
rect 24949 19012 24961 19015
rect 24044 18984 24961 19012
rect 24949 18981 24961 18984
rect 24995 18981 25007 19015
rect 25130 19012 25136 19024
rect 25091 18984 25136 19012
rect 24949 18975 25007 18981
rect 25130 18972 25136 18984
rect 25188 19012 25194 19024
rect 25685 19015 25743 19021
rect 25685 19012 25697 19015
rect 25188 18984 25697 19012
rect 25188 18972 25194 18984
rect 25685 18981 25697 18984
rect 25731 18981 25743 19015
rect 25685 18975 25743 18981
rect 13814 18944 13820 18956
rect 12667 18916 13820 18944
rect 12667 18913 12679 18916
rect 12621 18907 12679 18913
rect 13814 18904 13820 18916
rect 13872 18904 13878 18956
rect 15010 18944 15016 18956
rect 14971 18916 15016 18944
rect 15010 18904 15016 18916
rect 15068 18944 15074 18956
rect 15749 18947 15807 18953
rect 15749 18944 15761 18947
rect 15068 18916 15761 18944
rect 15068 18904 15074 18916
rect 15749 18913 15761 18916
rect 15795 18913 15807 18947
rect 17494 18944 17500 18956
rect 17407 18916 17500 18944
rect 15749 18907 15807 18913
rect 17494 18904 17500 18916
rect 17552 18944 17558 18956
rect 19705 18947 19763 18953
rect 19705 18944 19717 18947
rect 17552 18916 18092 18944
rect 17552 18904 17558 18916
rect 11054 18836 11060 18888
rect 11112 18876 11118 18888
rect 11149 18879 11207 18885
rect 11149 18876 11161 18879
rect 11112 18848 11161 18876
rect 11112 18836 11118 18848
rect 11149 18845 11161 18848
rect 11195 18845 11207 18879
rect 14090 18876 14096 18888
rect 14051 18848 14096 18876
rect 11149 18839 11207 18845
rect 14090 18836 14096 18848
rect 14148 18836 14154 18888
rect 15289 18879 15347 18885
rect 15289 18845 15301 18879
rect 15335 18876 15347 18879
rect 15378 18876 15384 18888
rect 15335 18848 15384 18876
rect 15335 18845 15347 18848
rect 15289 18839 15347 18845
rect 15378 18836 15384 18848
rect 15436 18836 15442 18888
rect 15657 18879 15715 18885
rect 15657 18845 15669 18879
rect 15703 18876 15715 18879
rect 16390 18876 16396 18888
rect 15703 18848 16396 18876
rect 15703 18845 15715 18848
rect 15657 18839 15715 18845
rect 16390 18836 16396 18848
rect 16448 18836 16454 18888
rect 17129 18879 17187 18885
rect 17129 18845 17141 18879
rect 17175 18876 17187 18879
rect 17310 18876 17316 18888
rect 17175 18848 17316 18876
rect 17175 18845 17187 18848
rect 17129 18839 17187 18845
rect 17310 18836 17316 18848
rect 17368 18836 17374 18888
rect 17586 18876 17592 18888
rect 17547 18848 17592 18876
rect 17586 18836 17592 18848
rect 17644 18836 17650 18888
rect 17678 18836 17684 18888
rect 17736 18876 17742 18888
rect 18064 18885 18092 18916
rect 19076 18916 19717 18944
rect 17957 18879 18015 18885
rect 17957 18876 17969 18879
rect 17736 18848 17969 18876
rect 17736 18836 17742 18848
rect 17957 18845 17969 18848
rect 18003 18845 18015 18879
rect 17957 18839 18015 18845
rect 18049 18879 18107 18885
rect 18049 18845 18061 18879
rect 18095 18876 18107 18879
rect 18138 18876 18144 18888
rect 18095 18848 18144 18876
rect 18095 18845 18107 18848
rect 18049 18839 18107 18845
rect 18138 18836 18144 18848
rect 18196 18836 18202 18888
rect 18966 18836 18972 18888
rect 19024 18876 19030 18888
rect 19076 18885 19104 18916
rect 19705 18913 19717 18916
rect 19751 18913 19763 18947
rect 19705 18907 19763 18913
rect 19794 18904 19800 18956
rect 19852 18944 19858 18956
rect 20257 18947 20315 18953
rect 20257 18944 20269 18947
rect 19852 18916 20269 18944
rect 19852 18904 19858 18916
rect 20257 18913 20269 18916
rect 20303 18944 20315 18947
rect 20625 18947 20683 18953
rect 20625 18944 20637 18947
rect 20303 18916 20637 18944
rect 20303 18913 20315 18916
rect 20257 18907 20315 18913
rect 20625 18913 20637 18916
rect 20671 18944 20683 18947
rect 20916 18944 20944 18972
rect 20671 18916 20944 18944
rect 20671 18913 20683 18916
rect 20625 18907 20683 18913
rect 21358 18904 21364 18956
rect 21416 18944 21422 18956
rect 23109 18947 23167 18953
rect 23109 18944 23121 18947
rect 21416 18916 23121 18944
rect 21416 18904 21422 18916
rect 23109 18913 23121 18916
rect 23155 18944 23167 18947
rect 24302 18944 24308 18956
rect 23155 18916 24308 18944
rect 23155 18913 23167 18916
rect 23109 18907 23167 18913
rect 24302 18904 24308 18916
rect 24360 18904 24366 18956
rect 19061 18879 19119 18885
rect 19061 18876 19073 18879
rect 19024 18848 19073 18876
rect 19024 18836 19030 18848
rect 19061 18845 19073 18848
rect 19107 18845 19119 18879
rect 19242 18876 19248 18888
rect 19203 18848 19248 18876
rect 19061 18839 19119 18845
rect 19242 18836 19248 18848
rect 19300 18836 19306 18888
rect 19334 18836 19340 18888
rect 19392 18876 19398 18888
rect 19613 18879 19671 18885
rect 19613 18876 19625 18879
rect 19392 18848 19625 18876
rect 19392 18836 19398 18848
rect 19613 18845 19625 18848
rect 19659 18876 19671 18879
rect 20162 18876 20168 18888
rect 19659 18848 20168 18876
rect 19659 18845 19671 18848
rect 19613 18839 19671 18845
rect 20162 18836 20168 18848
rect 20220 18836 20226 18888
rect 22278 18876 22284 18888
rect 22239 18848 22284 18876
rect 22278 18836 22284 18848
rect 22336 18836 22342 18888
rect 23566 18876 23572 18888
rect 23527 18848 23572 18876
rect 23566 18836 23572 18848
rect 23624 18836 23630 18888
rect 25314 18876 25320 18888
rect 25275 18848 25320 18876
rect 25314 18836 25320 18848
rect 25372 18836 25378 18888
rect 1104 18786 26864 18808
rect 1104 18734 10315 18786
rect 10367 18734 10379 18786
rect 10431 18734 10443 18786
rect 10495 18734 10507 18786
rect 10559 18734 19648 18786
rect 19700 18734 19712 18786
rect 19764 18734 19776 18786
rect 19828 18734 19840 18786
rect 19892 18734 26864 18786
rect 1104 18712 26864 18734
rect 11238 18672 11244 18684
rect 11199 18644 11244 18672
rect 11238 18632 11244 18644
rect 11296 18632 11302 18684
rect 11609 18675 11667 18681
rect 11609 18641 11621 18675
rect 11655 18672 11667 18675
rect 12802 18672 12808 18684
rect 11655 18644 12808 18672
rect 11655 18641 11667 18644
rect 11609 18635 11667 18641
rect 12802 18632 12808 18644
rect 12860 18632 12866 18684
rect 14182 18632 14188 18684
rect 14240 18672 14246 18684
rect 14826 18672 14832 18684
rect 14240 18644 14832 18672
rect 14240 18632 14246 18644
rect 14826 18632 14832 18644
rect 14884 18672 14890 18684
rect 15289 18675 15347 18681
rect 15289 18672 15301 18675
rect 14884 18644 15301 18672
rect 14884 18632 14890 18644
rect 15289 18641 15301 18644
rect 15335 18641 15347 18675
rect 15930 18672 15936 18684
rect 15891 18644 15936 18672
rect 15289 18635 15347 18641
rect 15930 18632 15936 18644
rect 15988 18632 15994 18684
rect 16945 18675 17003 18681
rect 16945 18641 16957 18675
rect 16991 18672 17003 18675
rect 17678 18672 17684 18684
rect 16991 18644 17684 18672
rect 16991 18641 17003 18644
rect 16945 18635 17003 18641
rect 17678 18632 17684 18644
rect 17736 18632 17742 18684
rect 18046 18632 18052 18684
rect 18104 18672 18110 18684
rect 18509 18675 18567 18681
rect 18509 18672 18521 18675
rect 18104 18644 18521 18672
rect 18104 18632 18110 18644
rect 18509 18641 18521 18644
rect 18555 18672 18567 18675
rect 19058 18672 19064 18684
rect 18555 18644 19064 18672
rect 18555 18641 18567 18644
rect 18509 18635 18567 18641
rect 19058 18632 19064 18644
rect 19116 18632 19122 18684
rect 19334 18672 19340 18684
rect 19295 18644 19340 18672
rect 19334 18632 19340 18644
rect 19392 18632 19398 18684
rect 21358 18632 21364 18684
rect 21416 18672 21422 18684
rect 21453 18675 21511 18681
rect 21453 18672 21465 18675
rect 21416 18644 21465 18672
rect 21416 18632 21422 18644
rect 21453 18641 21465 18644
rect 21499 18641 21511 18675
rect 21453 18635 21511 18641
rect 21913 18675 21971 18681
rect 21913 18641 21925 18675
rect 21959 18672 21971 18675
rect 22465 18675 22523 18681
rect 22465 18672 22477 18675
rect 21959 18644 22477 18672
rect 21959 18641 21971 18644
rect 21913 18635 21971 18641
rect 22465 18641 22477 18644
rect 22511 18672 22523 18675
rect 23566 18672 23572 18684
rect 22511 18644 23572 18672
rect 22511 18641 22523 18644
rect 22465 18635 22523 18641
rect 23566 18632 23572 18644
rect 23624 18632 23630 18684
rect 23658 18632 23664 18684
rect 23716 18672 23722 18684
rect 24121 18675 24179 18681
rect 24121 18672 24133 18675
rect 23716 18644 24133 18672
rect 23716 18632 23722 18644
rect 24121 18641 24133 18644
rect 24167 18672 24179 18675
rect 24486 18672 24492 18684
rect 24167 18644 24492 18672
rect 24167 18641 24179 18644
rect 24121 18635 24179 18641
rect 24486 18632 24492 18644
rect 24544 18632 24550 18684
rect 14090 18564 14096 18616
rect 14148 18604 14154 18616
rect 14553 18607 14611 18613
rect 14553 18604 14565 18607
rect 14148 18576 14565 18604
rect 14148 18564 14154 18576
rect 14553 18573 14565 18576
rect 14599 18604 14611 18607
rect 15948 18604 15976 18632
rect 14599 18576 15976 18604
rect 14599 18573 14611 18576
rect 14553 18567 14611 18573
rect 17586 18564 17592 18616
rect 17644 18604 17650 18616
rect 18417 18607 18475 18613
rect 18417 18604 18429 18607
rect 17644 18576 18429 18604
rect 17644 18564 17650 18576
rect 18417 18573 18429 18576
rect 18463 18604 18475 18607
rect 18598 18604 18604 18616
rect 18463 18576 18604 18604
rect 18463 18573 18475 18576
rect 18417 18567 18475 18573
rect 18598 18564 18604 18576
rect 18656 18564 18662 18616
rect 20809 18607 20867 18613
rect 20809 18573 20821 18607
rect 20855 18604 20867 18607
rect 21726 18604 21732 18616
rect 20855 18576 21732 18604
rect 20855 18573 20867 18576
rect 20809 18567 20867 18573
rect 21726 18564 21732 18576
rect 21784 18564 21790 18616
rect 23477 18607 23535 18613
rect 23477 18573 23489 18607
rect 23523 18604 23535 18607
rect 23934 18604 23940 18616
rect 23523 18576 23940 18604
rect 23523 18573 23535 18576
rect 23477 18567 23535 18573
rect 23934 18564 23940 18576
rect 23992 18564 23998 18616
rect 22373 18539 22431 18545
rect 22373 18505 22385 18539
rect 22419 18536 22431 18539
rect 23017 18539 23075 18545
rect 23017 18536 23029 18539
rect 22419 18508 23029 18536
rect 22419 18505 22431 18508
rect 22373 18499 22431 18505
rect 23017 18505 23029 18508
rect 23063 18505 23075 18539
rect 23017 18499 23075 18505
rect 15378 18468 15384 18480
rect 15339 18440 15384 18468
rect 15378 18428 15384 18440
rect 15436 18428 15442 18480
rect 15565 18471 15623 18477
rect 15565 18437 15577 18471
rect 15611 18468 15623 18471
rect 15838 18468 15844 18480
rect 15611 18440 15844 18468
rect 15611 18437 15623 18440
rect 15565 18431 15623 18437
rect 15838 18428 15844 18440
rect 15896 18428 15902 18480
rect 18230 18428 18236 18480
rect 18288 18468 18294 18480
rect 18601 18471 18659 18477
rect 18601 18468 18613 18471
rect 18288 18440 18613 18468
rect 18288 18428 18294 18440
rect 18601 18437 18613 18440
rect 18647 18437 18659 18471
rect 18601 18431 18659 18437
rect 20530 18428 20536 18480
rect 20588 18468 20594 18480
rect 20901 18471 20959 18477
rect 20901 18468 20913 18471
rect 20588 18440 20913 18468
rect 20588 18428 20594 18440
rect 20901 18437 20913 18440
rect 20947 18437 20959 18471
rect 20901 18431 20959 18437
rect 21085 18471 21143 18477
rect 21085 18437 21097 18471
rect 21131 18468 21143 18471
rect 22278 18468 22284 18480
rect 21131 18440 22284 18468
rect 21131 18437 21143 18440
rect 21085 18431 21143 18437
rect 19518 18360 19524 18412
rect 19576 18400 19582 18412
rect 20162 18400 20168 18412
rect 19576 18372 20168 18400
rect 19576 18360 19582 18372
rect 20162 18360 20168 18372
rect 20220 18400 20226 18412
rect 21100 18400 21128 18431
rect 22278 18428 22284 18440
rect 22336 18428 22342 18480
rect 22554 18428 22560 18480
rect 22612 18468 22618 18480
rect 22612 18440 22657 18468
rect 22612 18428 22618 18440
rect 20220 18372 21128 18400
rect 23032 18400 23060 18499
rect 23382 18496 23388 18548
rect 23440 18536 23446 18548
rect 24029 18539 24087 18545
rect 24029 18536 24041 18539
rect 23440 18508 24041 18536
rect 23440 18496 23446 18508
rect 24029 18505 24041 18508
rect 24075 18536 24087 18539
rect 24946 18536 24952 18548
rect 24075 18508 24952 18536
rect 24075 18505 24087 18508
rect 24029 18499 24087 18505
rect 24946 18496 24952 18508
rect 25004 18496 25010 18548
rect 25038 18496 25044 18548
rect 25096 18536 25102 18548
rect 25225 18539 25283 18545
rect 25225 18536 25237 18539
rect 25096 18508 25237 18536
rect 25096 18496 25102 18508
rect 25225 18505 25237 18508
rect 25271 18505 25283 18539
rect 25225 18499 25283 18505
rect 24302 18468 24308 18480
rect 24215 18440 24308 18468
rect 24302 18428 24308 18440
rect 24360 18468 24366 18480
rect 25498 18468 25504 18480
rect 24360 18440 25504 18468
rect 24360 18428 24366 18440
rect 25498 18428 25504 18440
rect 25556 18428 25562 18480
rect 23661 18403 23719 18409
rect 23661 18400 23673 18403
rect 23032 18372 23673 18400
rect 20220 18360 20226 18372
rect 23661 18369 23673 18372
rect 23707 18369 23719 18403
rect 23661 18363 23719 18369
rect 10870 18332 10876 18344
rect 10831 18304 10876 18332
rect 10870 18292 10876 18304
rect 10928 18292 10934 18344
rect 13725 18335 13783 18341
rect 13725 18301 13737 18335
rect 13771 18332 13783 18335
rect 14182 18332 14188 18344
rect 13771 18304 14188 18332
rect 13771 18301 13783 18304
rect 13725 18295 13783 18301
rect 14182 18292 14188 18304
rect 14240 18292 14246 18344
rect 14921 18335 14979 18341
rect 14921 18301 14933 18335
rect 14967 18332 14979 18335
rect 15286 18332 15292 18344
rect 14967 18304 15292 18332
rect 14967 18301 14979 18304
rect 14921 18295 14979 18301
rect 15286 18292 15292 18304
rect 15344 18292 15350 18344
rect 18046 18332 18052 18344
rect 18007 18304 18052 18332
rect 18046 18292 18052 18304
rect 18104 18292 18110 18344
rect 20441 18335 20499 18341
rect 20441 18301 20453 18335
rect 20487 18332 20499 18335
rect 20714 18332 20720 18344
rect 20487 18304 20720 18332
rect 20487 18301 20499 18304
rect 20441 18295 20499 18301
rect 20714 18292 20720 18304
rect 20772 18292 20778 18344
rect 22002 18332 22008 18344
rect 21963 18304 22008 18332
rect 22002 18292 22008 18304
rect 22060 18292 22066 18344
rect 24210 18292 24216 18344
rect 24268 18332 24274 18344
rect 24673 18335 24731 18341
rect 24673 18332 24685 18335
rect 24268 18304 24685 18332
rect 24268 18292 24274 18304
rect 24673 18301 24685 18304
rect 24719 18301 24731 18335
rect 25406 18332 25412 18344
rect 25367 18304 25412 18332
rect 24673 18295 24731 18301
rect 25406 18292 25412 18304
rect 25464 18292 25470 18344
rect 1104 18242 26864 18264
rect 1104 18190 5648 18242
rect 5700 18190 5712 18242
rect 5764 18190 5776 18242
rect 5828 18190 5840 18242
rect 5892 18190 14982 18242
rect 15034 18190 15046 18242
rect 15098 18190 15110 18242
rect 15162 18190 15174 18242
rect 15226 18190 24315 18242
rect 24367 18190 24379 18242
rect 24431 18190 24443 18242
rect 24495 18190 24507 18242
rect 24559 18190 26864 18242
rect 1104 18168 26864 18190
rect 10965 18131 11023 18137
rect 10965 18097 10977 18131
rect 11011 18128 11023 18131
rect 12250 18128 12256 18140
rect 11011 18100 12256 18128
rect 11011 18097 11023 18100
rect 10965 18091 11023 18097
rect 11072 18001 11100 18100
rect 12250 18088 12256 18100
rect 12308 18088 12314 18140
rect 12434 18088 12440 18140
rect 12492 18128 12498 18140
rect 12492 18100 12537 18128
rect 12492 18088 12498 18100
rect 14826 18088 14832 18140
rect 14884 18128 14890 18140
rect 14921 18131 14979 18137
rect 14921 18128 14933 18131
rect 14884 18100 14933 18128
rect 14884 18088 14890 18100
rect 14921 18097 14933 18100
rect 14967 18097 14979 18131
rect 14921 18091 14979 18097
rect 15378 18088 15384 18140
rect 15436 18128 15442 18140
rect 16117 18131 16175 18137
rect 16117 18128 16129 18131
rect 15436 18100 16129 18128
rect 15436 18088 15442 18100
rect 16117 18097 16129 18100
rect 16163 18097 16175 18131
rect 19058 18128 19064 18140
rect 19019 18100 19064 18128
rect 16117 18091 16175 18097
rect 19058 18088 19064 18100
rect 19116 18088 19122 18140
rect 20162 18128 20168 18140
rect 20123 18100 20168 18128
rect 20162 18088 20168 18100
rect 20220 18088 20226 18140
rect 20990 18088 20996 18140
rect 21048 18128 21054 18140
rect 21453 18131 21511 18137
rect 21453 18128 21465 18131
rect 21048 18100 21465 18128
rect 21048 18088 21054 18100
rect 21453 18097 21465 18100
rect 21499 18097 21511 18131
rect 24946 18128 24952 18140
rect 24907 18100 24952 18128
rect 21453 18091 21511 18097
rect 24946 18088 24952 18100
rect 25004 18088 25010 18140
rect 25038 18088 25044 18140
rect 25096 18128 25102 18140
rect 25685 18131 25743 18137
rect 25685 18128 25697 18131
rect 25096 18100 25697 18128
rect 25096 18088 25102 18100
rect 25685 18097 25697 18100
rect 25731 18097 25743 18131
rect 25685 18091 25743 18097
rect 15838 18060 15844 18072
rect 15799 18032 15844 18060
rect 15838 18020 15844 18032
rect 15896 18020 15902 18072
rect 21177 18063 21235 18069
rect 21177 18029 21189 18063
rect 21223 18060 21235 18063
rect 21726 18060 21732 18072
rect 21223 18032 21732 18060
rect 21223 18029 21235 18032
rect 21177 18023 21235 18029
rect 21726 18020 21732 18032
rect 21784 18020 21790 18072
rect 23474 18020 23480 18072
rect 23532 18060 23538 18072
rect 23937 18063 23995 18069
rect 23937 18060 23949 18063
rect 23532 18032 23949 18060
rect 23532 18020 23538 18032
rect 23937 18029 23949 18032
rect 23983 18029 23995 18063
rect 23937 18023 23995 18029
rect 25409 18063 25467 18069
rect 25409 18029 25421 18063
rect 25455 18060 25467 18063
rect 25498 18060 25504 18072
rect 25455 18032 25504 18060
rect 25455 18029 25467 18032
rect 25409 18023 25467 18029
rect 25498 18020 25504 18032
rect 25556 18020 25562 18072
rect 11057 17995 11115 18001
rect 11057 17961 11069 17995
rect 11103 17961 11115 17995
rect 14182 17992 14188 18004
rect 14143 17964 14188 17992
rect 11057 17955 11115 17961
rect 14182 17952 14188 17964
rect 14240 17952 14246 18004
rect 21913 17995 21971 18001
rect 21913 17961 21925 17995
rect 21959 17992 21971 17995
rect 22925 17995 22983 18001
rect 22925 17992 22937 17995
rect 21959 17964 22937 17992
rect 21959 17961 21971 17964
rect 21913 17955 21971 17961
rect 22925 17961 22937 17964
rect 22971 17992 22983 17995
rect 24210 17992 24216 18004
rect 22971 17964 24216 17992
rect 22971 17961 22983 17964
rect 22925 17955 22983 17961
rect 24210 17952 24216 17964
rect 24268 17992 24274 18004
rect 24489 17995 24547 18001
rect 24489 17992 24501 17995
rect 24268 17964 24501 17992
rect 24268 17952 24274 17964
rect 24489 17961 24501 17964
rect 24535 17961 24547 17995
rect 24489 17955 24547 17961
rect 13538 17884 13544 17936
rect 13596 17924 13602 17936
rect 14001 17927 14059 17933
rect 14001 17924 14013 17927
rect 13596 17896 14013 17924
rect 13596 17884 13602 17896
rect 14001 17893 14013 17896
rect 14047 17893 14059 17927
rect 15286 17924 15292 17936
rect 15247 17896 15292 17924
rect 14001 17887 14059 17893
rect 15286 17884 15292 17896
rect 15344 17924 15350 17936
rect 16485 17927 16543 17933
rect 16485 17924 16497 17927
rect 15344 17896 16497 17924
rect 15344 17884 15350 17896
rect 16485 17893 16497 17896
rect 16531 17893 16543 17927
rect 17129 17927 17187 17933
rect 17129 17924 17141 17927
rect 16485 17887 16543 17893
rect 16960 17896 17141 17924
rect 11146 17816 11152 17868
rect 11204 17856 11210 17868
rect 11302 17859 11360 17865
rect 11302 17856 11314 17859
rect 11204 17828 11314 17856
rect 11204 17816 11210 17828
rect 11302 17825 11314 17828
rect 11348 17825 11360 17859
rect 13446 17856 13452 17868
rect 13407 17828 13452 17856
rect 11302 17819 11360 17825
rect 13446 17816 13452 17828
rect 13504 17856 13510 17868
rect 14093 17859 14151 17865
rect 14093 17856 14105 17859
rect 13504 17828 14105 17856
rect 13504 17816 13510 17828
rect 14093 17825 14105 17828
rect 14139 17825 14151 17859
rect 14093 17819 14151 17825
rect 16960 17800 16988 17896
rect 17129 17893 17141 17896
rect 17175 17893 17187 17927
rect 17129 17887 17187 17893
rect 22462 17884 22468 17936
rect 22520 17924 22526 17936
rect 22741 17927 22799 17933
rect 22741 17924 22753 17927
rect 22520 17896 22753 17924
rect 22520 17884 22526 17896
rect 22741 17893 22753 17896
rect 22787 17924 22799 17927
rect 23198 17924 23204 17936
rect 22787 17896 23204 17924
rect 22787 17893 22799 17896
rect 22741 17887 22799 17893
rect 23198 17884 23204 17896
rect 23256 17884 23262 17936
rect 23477 17927 23535 17933
rect 23477 17893 23489 17927
rect 23523 17924 23535 17927
rect 23658 17924 23664 17936
rect 23523 17896 23664 17924
rect 23523 17893 23535 17896
rect 23477 17887 23535 17893
rect 23658 17884 23664 17896
rect 23716 17884 23722 17936
rect 23842 17924 23848 17936
rect 23755 17896 23848 17924
rect 23842 17884 23848 17896
rect 23900 17924 23906 17936
rect 24397 17927 24455 17933
rect 24397 17924 24409 17927
rect 23900 17896 24409 17924
rect 23900 17884 23906 17896
rect 24397 17893 24409 17896
rect 24443 17924 24455 17927
rect 25682 17924 25688 17936
rect 24443 17896 25688 17924
rect 24443 17893 24455 17896
rect 24397 17887 24455 17893
rect 25682 17884 25688 17896
rect 25740 17884 25746 17936
rect 17310 17816 17316 17868
rect 17368 17865 17374 17868
rect 17368 17859 17432 17865
rect 17368 17825 17386 17859
rect 17420 17825 17432 17859
rect 22186 17856 22192 17868
rect 22147 17828 22192 17856
rect 17368 17819 17432 17825
rect 17368 17816 17374 17819
rect 22186 17816 22192 17828
rect 22244 17856 22250 17868
rect 22833 17859 22891 17865
rect 22833 17856 22845 17859
rect 22244 17828 22845 17856
rect 22244 17816 22250 17828
rect 22833 17825 22845 17828
rect 22879 17825 22891 17859
rect 22833 17819 22891 17825
rect 13630 17788 13636 17800
rect 13591 17760 13636 17788
rect 13630 17748 13636 17760
rect 13688 17748 13694 17800
rect 15470 17788 15476 17800
rect 15431 17760 15476 17788
rect 15470 17748 15476 17760
rect 15528 17748 15534 17800
rect 16942 17788 16948 17800
rect 16903 17760 16948 17788
rect 16942 17748 16948 17760
rect 17000 17748 17006 17800
rect 18230 17748 18236 17800
rect 18288 17788 18294 17800
rect 18509 17791 18567 17797
rect 18509 17788 18521 17791
rect 18288 17760 18521 17788
rect 18288 17748 18294 17760
rect 18509 17757 18521 17760
rect 18555 17757 18567 17791
rect 20530 17788 20536 17800
rect 20491 17760 20536 17788
rect 18509 17751 18567 17757
rect 20530 17748 20536 17760
rect 20588 17748 20594 17800
rect 22373 17791 22431 17797
rect 22373 17757 22385 17791
rect 22419 17788 22431 17791
rect 22738 17788 22744 17800
rect 22419 17760 22744 17788
rect 22419 17757 22431 17760
rect 22373 17751 22431 17757
rect 22738 17748 22744 17760
rect 22796 17748 22802 17800
rect 23934 17748 23940 17800
rect 23992 17788 23998 17800
rect 24305 17791 24363 17797
rect 24305 17788 24317 17791
rect 23992 17760 24317 17788
rect 23992 17748 23998 17760
rect 24305 17757 24317 17760
rect 24351 17757 24363 17791
rect 24305 17751 24363 17757
rect 1104 17698 26864 17720
rect 1104 17646 10315 17698
rect 10367 17646 10379 17698
rect 10431 17646 10443 17698
rect 10495 17646 10507 17698
rect 10559 17646 19648 17698
rect 19700 17646 19712 17698
rect 19764 17646 19776 17698
rect 19828 17646 19840 17698
rect 19892 17646 26864 17698
rect 1104 17624 26864 17646
rect 13538 17544 13544 17596
rect 13596 17584 13602 17596
rect 13633 17587 13691 17593
rect 13633 17584 13645 17587
rect 13596 17556 13645 17584
rect 13596 17544 13602 17556
rect 13633 17553 13645 17556
rect 13679 17553 13691 17587
rect 18598 17584 18604 17596
rect 18559 17556 18604 17584
rect 13633 17547 13691 17553
rect 18598 17544 18604 17556
rect 18656 17544 18662 17596
rect 20714 17544 20720 17596
rect 20772 17584 20778 17596
rect 21729 17587 21787 17593
rect 21729 17584 21741 17587
rect 20772 17556 21741 17584
rect 20772 17544 20778 17556
rect 21729 17553 21741 17556
rect 21775 17584 21787 17587
rect 21910 17584 21916 17596
rect 21775 17556 21916 17584
rect 21775 17553 21787 17556
rect 21729 17547 21787 17553
rect 21910 17544 21916 17556
rect 21968 17544 21974 17596
rect 22462 17584 22468 17596
rect 22423 17556 22468 17584
rect 22462 17544 22468 17556
rect 22520 17544 22526 17596
rect 22738 17584 22744 17596
rect 22699 17556 22744 17584
rect 22738 17544 22744 17556
rect 22796 17544 22802 17596
rect 23201 17587 23259 17593
rect 23201 17553 23213 17587
rect 23247 17584 23259 17587
rect 23382 17584 23388 17596
rect 23247 17556 23388 17584
rect 23247 17553 23259 17556
rect 23201 17547 23259 17553
rect 23382 17544 23388 17556
rect 23440 17544 23446 17596
rect 23934 17584 23940 17596
rect 23895 17556 23940 17584
rect 23934 17544 23940 17556
rect 23992 17544 23998 17596
rect 25501 17587 25559 17593
rect 25501 17553 25513 17587
rect 25547 17584 25559 17587
rect 25774 17584 25780 17596
rect 25547 17556 25780 17584
rect 25547 17553 25559 17556
rect 25501 17547 25559 17553
rect 25774 17544 25780 17556
rect 25832 17544 25838 17596
rect 14185 17519 14243 17525
rect 14185 17485 14197 17519
rect 14231 17516 14243 17519
rect 14522 17519 14580 17525
rect 14522 17516 14534 17519
rect 14231 17488 14534 17516
rect 14231 17485 14243 17488
rect 14185 17479 14243 17485
rect 14522 17485 14534 17488
rect 14568 17516 14580 17519
rect 15102 17516 15108 17528
rect 14568 17488 15108 17516
rect 14568 17485 14580 17488
rect 14522 17479 14580 17485
rect 15102 17476 15108 17488
rect 15160 17476 15166 17528
rect 18230 17516 18236 17528
rect 18191 17488 18236 17516
rect 18230 17476 18236 17488
rect 18288 17476 18294 17528
rect 20346 17476 20352 17528
rect 20404 17516 20410 17528
rect 20898 17516 20904 17528
rect 20404 17488 20904 17516
rect 20404 17476 20410 17488
rect 20898 17476 20904 17488
rect 20956 17476 20962 17528
rect 21818 17516 21824 17528
rect 21779 17488 21824 17516
rect 21818 17476 21824 17488
rect 21876 17476 21882 17528
rect 13814 17408 13820 17460
rect 13872 17448 13878 17460
rect 14277 17451 14335 17457
rect 14277 17448 14289 17451
rect 13872 17420 14289 17448
rect 13872 17408 13878 17420
rect 14277 17417 14289 17420
rect 14323 17448 14335 17451
rect 14366 17448 14372 17460
rect 14323 17420 14372 17448
rect 14323 17417 14335 17420
rect 14277 17411 14335 17417
rect 14366 17408 14372 17420
rect 14424 17408 14430 17460
rect 20162 17448 20168 17460
rect 20123 17420 20168 17448
rect 20162 17408 20168 17420
rect 20220 17408 20226 17460
rect 24388 17451 24446 17457
rect 24388 17417 24400 17451
rect 24434 17448 24446 17451
rect 24762 17448 24768 17460
rect 24434 17420 24768 17448
rect 24434 17417 24446 17420
rect 24388 17411 24446 17417
rect 24762 17408 24768 17420
rect 24820 17408 24826 17460
rect 19150 17340 19156 17392
rect 19208 17380 19214 17392
rect 20254 17380 20260 17392
rect 19208 17352 20260 17380
rect 19208 17340 19214 17352
rect 20254 17340 20260 17352
rect 20312 17340 20318 17392
rect 20346 17340 20352 17392
rect 20404 17380 20410 17392
rect 20404 17352 20449 17380
rect 20404 17340 20410 17352
rect 21726 17340 21732 17392
rect 21784 17380 21790 17392
rect 21913 17383 21971 17389
rect 21913 17380 21925 17383
rect 21784 17352 21925 17380
rect 21784 17340 21790 17352
rect 21913 17349 21925 17352
rect 21959 17349 21971 17383
rect 21913 17343 21971 17349
rect 24026 17340 24032 17392
rect 24084 17380 24090 17392
rect 24121 17383 24179 17389
rect 24121 17380 24133 17383
rect 24084 17352 24133 17380
rect 24084 17340 24090 17352
rect 24121 17349 24133 17352
rect 24167 17349 24179 17383
rect 24121 17343 24179 17349
rect 19797 17315 19855 17321
rect 19797 17281 19809 17315
rect 19843 17312 19855 17315
rect 20990 17312 20996 17324
rect 19843 17284 20996 17312
rect 19843 17281 19855 17284
rect 19797 17275 19855 17281
rect 20990 17272 20996 17284
rect 21048 17272 21054 17324
rect 11146 17244 11152 17256
rect 11107 17216 11152 17244
rect 11146 17204 11152 17216
rect 11204 17204 11210 17256
rect 14182 17204 14188 17256
rect 14240 17244 14246 17256
rect 15657 17247 15715 17253
rect 15657 17244 15669 17247
rect 14240 17216 15669 17244
rect 14240 17204 14246 17216
rect 15657 17213 15669 17216
rect 15703 17244 15715 17247
rect 15838 17244 15844 17256
rect 15703 17216 15844 17244
rect 15703 17213 15715 17216
rect 15657 17207 15715 17213
rect 15838 17204 15844 17216
rect 15896 17204 15902 17256
rect 17221 17247 17279 17253
rect 17221 17213 17233 17247
rect 17267 17244 17279 17247
rect 17310 17244 17316 17256
rect 17267 17216 17316 17244
rect 17267 17213 17279 17216
rect 17221 17207 17279 17213
rect 17310 17204 17316 17216
rect 17368 17204 17374 17256
rect 21358 17244 21364 17256
rect 21319 17216 21364 17244
rect 21358 17204 21364 17216
rect 21416 17204 21422 17256
rect 1104 17154 26864 17176
rect 1104 17102 5648 17154
rect 5700 17102 5712 17154
rect 5764 17102 5776 17154
rect 5828 17102 5840 17154
rect 5892 17102 14982 17154
rect 15034 17102 15046 17154
rect 15098 17102 15110 17154
rect 15162 17102 15174 17154
rect 15226 17102 24315 17154
rect 24367 17102 24379 17154
rect 24431 17102 24443 17154
rect 24495 17102 24507 17154
rect 24559 17102 26864 17154
rect 1104 17080 26864 17102
rect 14642 17000 14648 17052
rect 14700 17040 14706 17052
rect 15013 17043 15071 17049
rect 15013 17040 15025 17043
rect 14700 17012 15025 17040
rect 14700 17000 14706 17012
rect 15013 17009 15025 17012
rect 15059 17009 15071 17043
rect 15013 17003 15071 17009
rect 11146 16932 11152 16984
rect 11204 16972 11210 16984
rect 11204 16944 13584 16972
rect 11204 16932 11210 16944
rect 13556 16845 13584 16944
rect 13630 16864 13636 16916
rect 13688 16904 13694 16916
rect 14093 16907 14151 16913
rect 14093 16904 14105 16907
rect 13688 16876 14105 16904
rect 13688 16864 13694 16876
rect 14093 16873 14105 16876
rect 14139 16873 14151 16907
rect 14274 16904 14280 16916
rect 14235 16876 14280 16904
rect 14093 16867 14151 16873
rect 14274 16864 14280 16876
rect 14332 16864 14338 16916
rect 14366 16864 14372 16916
rect 14424 16904 14430 16916
rect 14645 16907 14703 16913
rect 14645 16904 14657 16907
rect 14424 16876 14657 16904
rect 14424 16864 14430 16876
rect 14645 16873 14657 16876
rect 14691 16873 14703 16907
rect 14645 16867 14703 16873
rect 13541 16839 13599 16845
rect 13541 16805 13553 16839
rect 13587 16836 13599 16839
rect 14292 16836 14320 16864
rect 13587 16808 14320 16836
rect 15028 16836 15056 17003
rect 17310 17000 17316 17052
rect 17368 17040 17374 17052
rect 18417 17043 18475 17049
rect 18417 17040 18429 17043
rect 17368 17012 18429 17040
rect 17368 17000 17374 17012
rect 18417 17009 18429 17012
rect 18463 17009 18475 17043
rect 19150 17040 19156 17052
rect 19111 17012 19156 17040
rect 18417 17003 18475 17009
rect 19150 17000 19156 17012
rect 19208 17000 19214 17052
rect 19889 17043 19947 17049
rect 19889 17009 19901 17043
rect 19935 17040 19947 17043
rect 20162 17040 20168 17052
rect 19935 17012 20168 17040
rect 19935 17009 19947 17012
rect 19889 17003 19947 17009
rect 20162 17000 20168 17012
rect 20220 17000 20226 17052
rect 20254 17000 20260 17052
rect 20312 17040 20318 17052
rect 20901 17043 20959 17049
rect 20901 17040 20913 17043
rect 20312 17012 20913 17040
rect 20312 17000 20318 17012
rect 20901 17009 20913 17012
rect 20947 17009 20959 17043
rect 20901 17003 20959 17009
rect 23474 17000 23480 17052
rect 23532 17040 23538 17052
rect 24026 17040 24032 17052
rect 23532 17012 24032 17040
rect 23532 17000 23538 17012
rect 24026 17000 24032 17012
rect 24084 17000 24090 17052
rect 22649 16975 22707 16981
rect 22649 16941 22661 16975
rect 22695 16972 22707 16975
rect 25225 16975 25283 16981
rect 25225 16972 25237 16975
rect 22695 16944 25237 16972
rect 22695 16941 22707 16944
rect 22649 16935 22707 16941
rect 15838 16904 15844 16916
rect 15799 16876 15844 16904
rect 15838 16864 15844 16876
rect 15896 16864 15902 16916
rect 16942 16864 16948 16916
rect 17000 16904 17006 16916
rect 17037 16907 17095 16913
rect 17037 16904 17049 16907
rect 17000 16876 17049 16904
rect 17000 16864 17006 16876
rect 17037 16873 17049 16876
rect 17083 16873 17095 16907
rect 17037 16867 17095 16873
rect 20070 16864 20076 16916
rect 20128 16904 20134 16916
rect 20257 16907 20315 16913
rect 20257 16904 20269 16907
rect 20128 16876 20269 16904
rect 20128 16864 20134 16876
rect 20257 16873 20269 16876
rect 20303 16904 20315 16907
rect 21453 16907 21511 16913
rect 21453 16904 21465 16907
rect 20303 16876 21465 16904
rect 20303 16873 20315 16876
rect 20257 16867 20315 16873
rect 21453 16873 21465 16876
rect 21499 16873 21511 16907
rect 23198 16904 23204 16916
rect 23159 16876 23204 16904
rect 21453 16867 21511 16873
rect 23198 16864 23204 16876
rect 23256 16864 23262 16916
rect 24688 16913 24716 16944
rect 25225 16941 25237 16944
rect 25271 16941 25283 16975
rect 25225 16935 25283 16941
rect 26234 16932 26240 16984
rect 26292 16972 26298 16984
rect 27522 16972 27528 16984
rect 26292 16944 27528 16972
rect 26292 16932 26298 16944
rect 27522 16932 27528 16944
rect 27580 16932 27586 16984
rect 24673 16907 24731 16913
rect 24673 16873 24685 16907
rect 24719 16873 24731 16907
rect 24673 16867 24731 16873
rect 24857 16907 24915 16913
rect 24857 16873 24869 16907
rect 24903 16873 24915 16907
rect 24857 16867 24915 16873
rect 15746 16836 15752 16848
rect 15028 16808 15752 16836
rect 13587 16805 13599 16808
rect 13541 16799 13599 16805
rect 15746 16796 15752 16808
rect 15804 16796 15810 16848
rect 16850 16796 16856 16848
rect 16908 16796 16914 16848
rect 20714 16836 20720 16848
rect 20675 16808 20720 16836
rect 20714 16796 20720 16808
rect 20772 16796 20778 16848
rect 20898 16796 20904 16848
rect 20956 16836 20962 16848
rect 21361 16839 21419 16845
rect 21361 16836 21373 16839
rect 20956 16808 21373 16836
rect 20956 16796 20962 16808
rect 21361 16805 21373 16808
rect 21407 16836 21419 16839
rect 21634 16836 21640 16848
rect 21407 16808 21640 16836
rect 21407 16805 21419 16808
rect 21361 16799 21419 16805
rect 21634 16796 21640 16808
rect 21692 16796 21698 16848
rect 23017 16839 23075 16845
rect 23017 16805 23029 16839
rect 23063 16836 23075 16839
rect 23382 16836 23388 16848
rect 23063 16808 23388 16836
rect 23063 16805 23075 16808
rect 23017 16799 23075 16805
rect 23382 16796 23388 16808
rect 23440 16796 23446 16848
rect 23753 16839 23811 16845
rect 23753 16805 23765 16839
rect 23799 16836 23811 16839
rect 23799 16808 24716 16836
rect 23799 16805 23811 16808
rect 23753 16799 23811 16805
rect 13173 16771 13231 16777
rect 13173 16737 13185 16771
rect 13219 16768 13231 16771
rect 14001 16771 14059 16777
rect 14001 16768 14013 16771
rect 13219 16740 14013 16768
rect 13219 16737 13231 16740
rect 13173 16731 13231 16737
rect 14001 16737 14013 16740
rect 14047 16768 14059 16771
rect 15654 16768 15660 16780
rect 14047 16740 15332 16768
rect 15567 16740 15660 16768
rect 14047 16737 14059 16740
rect 14001 16731 14059 16737
rect 13633 16703 13691 16709
rect 13633 16669 13645 16703
rect 13679 16700 13691 16703
rect 13814 16700 13820 16712
rect 13679 16672 13820 16700
rect 13679 16669 13691 16672
rect 13633 16663 13691 16669
rect 13814 16660 13820 16672
rect 13872 16660 13878 16712
rect 15304 16709 15332 16740
rect 15654 16728 15660 16740
rect 15712 16768 15718 16780
rect 16301 16771 16359 16777
rect 16301 16768 16313 16771
rect 15712 16740 16313 16768
rect 15712 16728 15718 16740
rect 16301 16737 16313 16740
rect 16347 16737 16359 16771
rect 16868 16768 16896 16796
rect 17282 16771 17340 16777
rect 17282 16768 17294 16771
rect 16868 16740 17294 16768
rect 16301 16731 16359 16737
rect 17282 16737 17294 16740
rect 17328 16737 17340 16771
rect 20732 16768 20760 16796
rect 21269 16771 21327 16777
rect 21269 16768 21281 16771
rect 20732 16740 21281 16768
rect 17282 16731 17340 16737
rect 21269 16737 21281 16740
rect 21315 16737 21327 16771
rect 21269 16731 21327 16737
rect 22738 16728 22744 16780
rect 22796 16768 22802 16780
rect 23109 16771 23167 16777
rect 23109 16768 23121 16771
rect 22796 16740 23121 16768
rect 22796 16728 22802 16740
rect 23109 16737 23121 16740
rect 23155 16737 23167 16771
rect 23109 16731 23167 16737
rect 23842 16728 23848 16780
rect 23900 16768 23906 16780
rect 24688 16768 24716 16808
rect 24762 16768 24768 16780
rect 23900 16740 24256 16768
rect 24675 16740 24768 16768
rect 23900 16728 23906 16740
rect 15289 16703 15347 16709
rect 15289 16669 15301 16703
rect 15335 16669 15347 16703
rect 16942 16700 16948 16712
rect 16903 16672 16948 16700
rect 15289 16663 15347 16669
rect 16942 16660 16948 16672
rect 17000 16660 17006 16712
rect 19426 16700 19432 16712
rect 19387 16672 19432 16700
rect 19426 16660 19432 16672
rect 19484 16660 19490 16712
rect 21726 16660 21732 16712
rect 21784 16700 21790 16712
rect 21913 16703 21971 16709
rect 21913 16700 21925 16703
rect 21784 16672 21925 16700
rect 21784 16660 21790 16672
rect 21913 16669 21925 16672
rect 21959 16669 21971 16703
rect 21913 16663 21971 16669
rect 22557 16703 22615 16709
rect 22557 16669 22569 16703
rect 22603 16700 22615 16703
rect 23198 16700 23204 16712
rect 22603 16672 23204 16700
rect 22603 16669 22615 16672
rect 22557 16663 22615 16669
rect 23198 16660 23204 16672
rect 23256 16660 23262 16712
rect 24228 16709 24256 16740
rect 24762 16728 24768 16740
rect 24820 16768 24826 16780
rect 24872 16768 24900 16867
rect 24820 16740 24900 16768
rect 24820 16728 24826 16740
rect 24213 16703 24271 16709
rect 24213 16669 24225 16703
rect 24259 16669 24271 16703
rect 24578 16700 24584 16712
rect 24539 16672 24584 16700
rect 24213 16663 24271 16669
rect 24578 16660 24584 16672
rect 24636 16660 24642 16712
rect 1104 16610 26864 16632
rect 1104 16558 10315 16610
rect 10367 16558 10379 16610
rect 10431 16558 10443 16610
rect 10495 16558 10507 16610
rect 10559 16558 19648 16610
rect 19700 16558 19712 16610
rect 19764 16558 19776 16610
rect 19828 16558 19840 16610
rect 19892 16558 26864 16610
rect 1104 16536 26864 16558
rect 13630 16496 13636 16508
rect 13591 16468 13636 16496
rect 13630 16456 13636 16468
rect 13688 16456 13694 16508
rect 14274 16456 14280 16508
rect 14332 16496 14338 16508
rect 15473 16499 15531 16505
rect 15473 16496 15485 16499
rect 14332 16468 15485 16496
rect 14332 16456 14338 16468
rect 15473 16465 15485 16468
rect 15519 16465 15531 16499
rect 15473 16459 15531 16465
rect 15838 16456 15844 16508
rect 15896 16496 15902 16508
rect 16025 16499 16083 16505
rect 16025 16496 16037 16499
rect 15896 16468 16037 16496
rect 15896 16456 15902 16468
rect 16025 16465 16037 16468
rect 16071 16465 16083 16499
rect 16025 16459 16083 16465
rect 16850 16456 16856 16508
rect 16908 16496 16914 16508
rect 17129 16499 17187 16505
rect 17129 16496 17141 16499
rect 16908 16468 17141 16496
rect 16908 16456 16914 16468
rect 17129 16465 17141 16468
rect 17175 16496 17187 16499
rect 17954 16496 17960 16508
rect 17175 16468 17960 16496
rect 17175 16465 17187 16468
rect 17129 16459 17187 16465
rect 17954 16456 17960 16468
rect 18012 16456 18018 16508
rect 19426 16456 19432 16508
rect 19484 16496 19490 16508
rect 20346 16496 20352 16508
rect 19484 16468 20352 16496
rect 19484 16456 19490 16468
rect 20346 16456 20352 16468
rect 20404 16496 20410 16508
rect 20993 16499 21051 16505
rect 20993 16496 21005 16499
rect 20404 16468 21005 16496
rect 20404 16456 20410 16468
rect 20993 16465 21005 16468
rect 21039 16496 21051 16499
rect 21726 16496 21732 16508
rect 21039 16468 21732 16496
rect 21039 16465 21051 16468
rect 20993 16459 21051 16465
rect 21726 16456 21732 16468
rect 21784 16456 21790 16508
rect 21910 16496 21916 16508
rect 21871 16468 21916 16496
rect 21910 16456 21916 16468
rect 21968 16456 21974 16508
rect 23658 16456 23664 16508
rect 23716 16496 23722 16508
rect 24029 16499 24087 16505
rect 24029 16496 24041 16499
rect 23716 16468 24041 16496
rect 23716 16456 23722 16468
rect 24029 16465 24041 16468
rect 24075 16465 24087 16499
rect 24762 16496 24768 16508
rect 24723 16468 24768 16496
rect 24029 16459 24087 16465
rect 24762 16456 24768 16468
rect 24820 16456 24826 16508
rect 25406 16496 25412 16508
rect 25367 16468 25412 16496
rect 25406 16456 25412 16468
rect 25464 16456 25470 16508
rect 14182 16388 14188 16440
rect 14240 16428 14246 16440
rect 14360 16431 14418 16437
rect 14360 16428 14372 16431
rect 14240 16400 14372 16428
rect 14240 16388 14246 16400
rect 14360 16397 14372 16400
rect 14406 16397 14418 16431
rect 14360 16391 14418 16397
rect 14458 16388 14464 16440
rect 14516 16388 14522 16440
rect 19880 16431 19938 16437
rect 19880 16397 19892 16431
rect 19926 16428 19938 16431
rect 20070 16428 20076 16440
rect 19926 16400 20076 16428
rect 19926 16397 19938 16400
rect 19880 16391 19938 16397
rect 20070 16388 20076 16400
rect 20128 16388 20134 16440
rect 21637 16431 21695 16437
rect 21637 16397 21649 16431
rect 21683 16428 21695 16431
rect 21818 16428 21824 16440
rect 21683 16400 21824 16428
rect 21683 16397 21695 16400
rect 21637 16391 21695 16397
rect 21818 16388 21824 16400
rect 21876 16388 21882 16440
rect 21928 16400 22140 16428
rect 14093 16363 14151 16369
rect 14093 16329 14105 16363
rect 14139 16360 14151 16363
rect 14476 16360 14504 16388
rect 21928 16360 21956 16400
rect 14139 16332 14504 16360
rect 19628 16332 21956 16360
rect 14139 16329 14151 16332
rect 14093 16323 14151 16329
rect 19628 16304 19656 16332
rect 22112 16304 22140 16400
rect 24118 16388 24124 16440
rect 24176 16428 24182 16440
rect 24578 16428 24584 16440
rect 24176 16400 24584 16428
rect 24176 16388 24182 16400
rect 24578 16388 24584 16400
rect 24636 16428 24642 16440
rect 25041 16431 25099 16437
rect 25041 16428 25053 16431
rect 24636 16400 25053 16428
rect 24636 16388 24642 16400
rect 25041 16397 25053 16400
rect 25087 16397 25099 16431
rect 25041 16391 25099 16397
rect 22557 16363 22615 16369
rect 22557 16329 22569 16363
rect 22603 16360 22615 16363
rect 23474 16360 23480 16372
rect 22603 16332 23480 16360
rect 22603 16329 22615 16332
rect 22557 16323 22615 16329
rect 23474 16320 23480 16332
rect 23532 16320 23538 16372
rect 23934 16320 23940 16372
rect 23992 16320 23998 16372
rect 24854 16360 24860 16372
rect 24136 16332 24860 16360
rect 19610 16292 19616 16304
rect 19571 16264 19616 16292
rect 19610 16252 19616 16264
rect 19668 16252 19674 16304
rect 22094 16252 22100 16304
rect 22152 16252 22158 16304
rect 23952 16292 23980 16320
rect 24136 16301 24164 16332
rect 24854 16320 24860 16332
rect 24912 16320 24918 16372
rect 25222 16360 25228 16372
rect 25183 16332 25228 16360
rect 25222 16320 25228 16332
rect 25280 16320 25286 16372
rect 24121 16295 24179 16301
rect 24121 16292 24133 16295
rect 23952 16264 24133 16292
rect 24121 16261 24133 16264
rect 24167 16261 24179 16295
rect 24302 16292 24308 16304
rect 24263 16264 24308 16292
rect 24121 16255 24179 16261
rect 24302 16252 24308 16264
rect 24360 16252 24366 16304
rect 23014 16184 23020 16236
rect 23072 16224 23078 16236
rect 24320 16224 24348 16252
rect 23072 16196 24348 16224
rect 23072 16184 23078 16196
rect 23198 16156 23204 16168
rect 23159 16128 23204 16156
rect 23198 16116 23204 16128
rect 23256 16116 23262 16168
rect 23658 16156 23664 16168
rect 23619 16128 23664 16156
rect 23658 16116 23664 16128
rect 23716 16116 23722 16168
rect 1104 16066 26864 16088
rect 1104 16014 5648 16066
rect 5700 16014 5712 16066
rect 5764 16014 5776 16066
rect 5828 16014 5840 16066
rect 5892 16014 14982 16066
rect 15034 16014 15046 16066
rect 15098 16014 15110 16066
rect 15162 16014 15174 16066
rect 15226 16014 24315 16066
rect 24367 16014 24379 16066
rect 24431 16014 24443 16066
rect 24495 16014 24507 16066
rect 24559 16014 26864 16066
rect 1104 15992 26864 16014
rect 14093 15955 14151 15961
rect 14093 15921 14105 15955
rect 14139 15952 14151 15955
rect 14182 15952 14188 15964
rect 14139 15924 14188 15952
rect 14139 15921 14151 15924
rect 14093 15915 14151 15921
rect 14182 15912 14188 15924
rect 14240 15912 14246 15964
rect 14458 15912 14464 15964
rect 14516 15952 14522 15964
rect 14645 15955 14703 15961
rect 14645 15952 14657 15955
rect 14516 15924 14657 15952
rect 14516 15912 14522 15924
rect 14645 15921 14657 15924
rect 14691 15952 14703 15955
rect 16853 15955 16911 15961
rect 16853 15952 16865 15955
rect 14691 15924 16865 15952
rect 14691 15921 14703 15924
rect 14645 15915 14703 15921
rect 16853 15921 16865 15924
rect 16899 15952 16911 15955
rect 16942 15952 16948 15964
rect 16899 15924 16948 15952
rect 16899 15921 16911 15924
rect 16853 15915 16911 15921
rect 16942 15912 16948 15924
rect 17000 15952 17006 15964
rect 17000 15924 17080 15952
rect 17000 15912 17006 15924
rect 15289 15819 15347 15825
rect 15289 15785 15301 15819
rect 15335 15816 15347 15819
rect 15654 15816 15660 15828
rect 15335 15788 15660 15816
rect 15335 15785 15347 15788
rect 15289 15779 15347 15785
rect 15654 15776 15660 15788
rect 15712 15776 15718 15828
rect 17052 15825 17080 15924
rect 17954 15912 17960 15964
rect 18012 15952 18018 15964
rect 18417 15955 18475 15961
rect 18417 15952 18429 15955
rect 18012 15924 18429 15952
rect 18012 15912 18018 15924
rect 18417 15921 18429 15924
rect 18463 15921 18475 15955
rect 18417 15915 18475 15921
rect 20070 15912 20076 15964
rect 20128 15952 20134 15964
rect 20257 15955 20315 15961
rect 20257 15952 20269 15955
rect 20128 15924 20269 15952
rect 20128 15912 20134 15924
rect 20257 15921 20269 15924
rect 20303 15921 20315 15955
rect 20257 15915 20315 15921
rect 22094 15912 22100 15964
rect 22152 15952 22158 15964
rect 23017 15955 23075 15961
rect 23017 15952 23029 15955
rect 22152 15924 23029 15952
rect 22152 15912 22158 15924
rect 23017 15921 23029 15924
rect 23063 15952 23075 15955
rect 23382 15952 23388 15964
rect 23063 15924 23388 15952
rect 23063 15921 23075 15924
rect 23017 15915 23075 15921
rect 23124 15828 23152 15924
rect 23382 15912 23388 15924
rect 23440 15912 23446 15964
rect 24489 15955 24547 15961
rect 24489 15921 24501 15955
rect 24535 15952 24547 15955
rect 24762 15952 24768 15964
rect 24535 15924 24768 15952
rect 24535 15921 24547 15924
rect 24489 15915 24547 15921
rect 24762 15912 24768 15924
rect 24820 15912 24826 15964
rect 25038 15952 25044 15964
rect 24999 15924 25044 15952
rect 25038 15912 25044 15924
rect 25096 15912 25102 15964
rect 25222 15912 25228 15964
rect 25280 15952 25286 15964
rect 25777 15955 25835 15961
rect 25777 15952 25789 15955
rect 25280 15924 25789 15952
rect 25280 15912 25286 15924
rect 25777 15921 25789 15924
rect 25823 15921 25835 15955
rect 25777 15915 25835 15921
rect 24854 15844 24860 15896
rect 24912 15884 24918 15896
rect 25409 15887 25467 15893
rect 25409 15884 25421 15887
rect 24912 15856 25421 15884
rect 24912 15844 24918 15856
rect 25409 15853 25421 15856
rect 25455 15853 25467 15887
rect 25409 15847 25467 15853
rect 17037 15819 17095 15825
rect 17037 15785 17049 15819
rect 17083 15785 17095 15819
rect 17037 15779 17095 15785
rect 19797 15819 19855 15825
rect 19797 15785 19809 15819
rect 19843 15816 19855 15819
rect 20162 15816 20168 15828
rect 19843 15788 20168 15816
rect 19843 15785 19855 15788
rect 19797 15779 19855 15785
rect 11054 15708 11060 15760
rect 11112 15748 11118 15760
rect 12069 15751 12127 15757
rect 12069 15748 12081 15751
rect 11112 15720 12081 15748
rect 11112 15708 11118 15720
rect 12069 15717 12081 15720
rect 12115 15748 12127 15751
rect 12529 15751 12587 15757
rect 12529 15748 12541 15751
rect 12115 15720 12541 15748
rect 12115 15717 12127 15720
rect 12069 15711 12127 15717
rect 12529 15717 12541 15720
rect 12575 15717 12587 15751
rect 12529 15711 12587 15717
rect 13814 15708 13820 15760
rect 13872 15748 13878 15760
rect 14185 15751 14243 15757
rect 14185 15748 14197 15751
rect 13872 15720 14197 15748
rect 13872 15708 13878 15720
rect 14185 15717 14197 15720
rect 14231 15748 14243 15751
rect 15013 15751 15071 15757
rect 15013 15748 15025 15751
rect 14231 15720 15025 15748
rect 14231 15717 14243 15720
rect 14185 15711 14243 15717
rect 15013 15717 15025 15720
rect 15059 15717 15071 15751
rect 17052 15748 17080 15779
rect 20162 15776 20168 15788
rect 20220 15776 20226 15828
rect 21358 15816 21364 15828
rect 21319 15788 21364 15816
rect 21358 15776 21364 15788
rect 21416 15776 21422 15828
rect 21453 15819 21511 15825
rect 21453 15785 21465 15819
rect 21499 15785 21511 15819
rect 23106 15816 23112 15828
rect 23019 15788 23112 15816
rect 21453 15779 21511 15785
rect 17678 15748 17684 15760
rect 17052 15720 17684 15748
rect 15013 15711 15071 15717
rect 17678 15708 17684 15720
rect 17736 15748 17742 15760
rect 19150 15748 19156 15760
rect 17736 15720 19156 15748
rect 17736 15708 17742 15720
rect 19150 15708 19156 15720
rect 19208 15748 19214 15760
rect 19610 15748 19616 15760
rect 19208 15720 19616 15748
rect 19208 15708 19214 15720
rect 19610 15708 19616 15720
rect 19668 15708 19674 15760
rect 21468 15748 21496 15779
rect 23106 15776 23112 15788
rect 23164 15776 23170 15828
rect 20640 15720 21496 15748
rect 17126 15640 17132 15692
rect 17184 15680 17190 15692
rect 17282 15683 17340 15689
rect 17282 15680 17294 15683
rect 17184 15652 17294 15680
rect 17184 15640 17190 15652
rect 17282 15649 17294 15652
rect 17328 15649 17340 15683
rect 17282 15643 17340 15649
rect 20640 15624 20668 15720
rect 20916 15652 22048 15680
rect 12250 15612 12256 15624
rect 12211 15584 12256 15612
rect 12250 15572 12256 15584
rect 12308 15572 12314 15624
rect 14366 15612 14372 15624
rect 14327 15584 14372 15612
rect 14366 15572 14372 15584
rect 14424 15572 14430 15624
rect 20622 15612 20628 15624
rect 20583 15584 20628 15612
rect 20622 15572 20628 15584
rect 20680 15572 20686 15624
rect 20916 15621 20944 15652
rect 20901 15615 20959 15621
rect 20901 15581 20913 15615
rect 20947 15581 20959 15615
rect 20901 15575 20959 15581
rect 20990 15572 20996 15624
rect 21048 15612 21054 15624
rect 21269 15615 21327 15621
rect 21269 15612 21281 15615
rect 21048 15584 21281 15612
rect 21048 15572 21054 15584
rect 21269 15581 21281 15584
rect 21315 15612 21327 15615
rect 21913 15615 21971 15621
rect 21913 15612 21925 15615
rect 21315 15584 21925 15612
rect 21315 15581 21327 15584
rect 21269 15575 21327 15581
rect 21913 15581 21925 15584
rect 21959 15581 21971 15615
rect 22020 15612 22048 15652
rect 23198 15640 23204 15692
rect 23256 15680 23262 15692
rect 23376 15683 23434 15689
rect 23376 15680 23388 15683
rect 23256 15652 23388 15680
rect 23256 15640 23262 15652
rect 23376 15649 23388 15652
rect 23422 15680 23434 15683
rect 24302 15680 24308 15692
rect 23422 15652 24308 15680
rect 23422 15649 23434 15652
rect 23376 15643 23434 15649
rect 24302 15640 24308 15652
rect 24360 15640 24366 15692
rect 22094 15612 22100 15624
rect 22020 15584 22100 15612
rect 21913 15575 21971 15581
rect 22094 15572 22100 15584
rect 22152 15572 22158 15624
rect 1104 15522 26864 15544
rect 1104 15470 10315 15522
rect 10367 15470 10379 15522
rect 10431 15470 10443 15522
rect 10495 15470 10507 15522
rect 10559 15470 19648 15522
rect 19700 15470 19712 15522
rect 19764 15470 19776 15522
rect 19828 15470 19840 15522
rect 19892 15470 26864 15522
rect 1104 15448 26864 15470
rect 12526 15368 12532 15420
rect 12584 15408 12590 15420
rect 12621 15411 12679 15417
rect 12621 15408 12633 15411
rect 12584 15380 12633 15408
rect 12584 15368 12590 15380
rect 12621 15377 12633 15380
rect 12667 15377 12679 15411
rect 12621 15371 12679 15377
rect 14734 15368 14740 15420
rect 14792 15408 14798 15420
rect 14829 15411 14887 15417
rect 14829 15408 14841 15411
rect 14792 15380 14841 15408
rect 14792 15368 14798 15380
rect 14829 15377 14841 15380
rect 14875 15377 14887 15411
rect 17126 15408 17132 15420
rect 17087 15380 17132 15408
rect 14829 15371 14887 15377
rect 17126 15368 17132 15380
rect 17184 15408 17190 15420
rect 20533 15411 20591 15417
rect 20533 15408 20545 15411
rect 17184 15380 20545 15408
rect 17184 15368 17190 15380
rect 20533 15377 20545 15380
rect 20579 15408 20591 15411
rect 20622 15408 20628 15420
rect 20579 15380 20628 15408
rect 20579 15377 20591 15380
rect 20533 15371 20591 15377
rect 20622 15368 20628 15380
rect 20680 15368 20686 15420
rect 21177 15411 21235 15417
rect 21177 15377 21189 15411
rect 21223 15408 21235 15411
rect 21358 15408 21364 15420
rect 21223 15380 21364 15408
rect 21223 15377 21235 15380
rect 21177 15371 21235 15377
rect 21358 15368 21364 15380
rect 21416 15368 21422 15420
rect 23014 15368 23020 15420
rect 23072 15408 23078 15420
rect 23385 15411 23443 15417
rect 23385 15408 23397 15411
rect 23072 15380 23397 15408
rect 23072 15368 23078 15380
rect 23385 15377 23397 15380
rect 23431 15377 23443 15411
rect 23385 15371 23443 15377
rect 23658 15368 23664 15420
rect 23716 15408 23722 15420
rect 24121 15411 24179 15417
rect 24121 15408 24133 15411
rect 23716 15380 24133 15408
rect 23716 15368 23722 15380
rect 24121 15377 24133 15380
rect 24167 15377 24179 15411
rect 24670 15408 24676 15420
rect 24631 15380 24676 15408
rect 24121 15371 24179 15377
rect 24670 15368 24676 15380
rect 24728 15368 24734 15420
rect 25406 15408 25412 15420
rect 25367 15380 25412 15408
rect 25406 15368 25412 15380
rect 25464 15368 25470 15420
rect 23474 15300 23480 15352
rect 23532 15340 23538 15352
rect 24026 15340 24032 15352
rect 23532 15312 24032 15340
rect 23532 15300 23538 15312
rect 24026 15300 24032 15312
rect 24084 15300 24090 15352
rect 12434 15232 12440 15284
rect 12492 15272 12498 15284
rect 14642 15272 14648 15284
rect 12492 15244 12537 15272
rect 14603 15244 14648 15272
rect 12492 15232 12498 15244
rect 14642 15232 14648 15244
rect 14700 15232 14706 15284
rect 19150 15272 19156 15284
rect 19111 15244 19156 15272
rect 19150 15232 19156 15244
rect 19208 15232 19214 15284
rect 19426 15281 19432 15284
rect 19420 15272 19432 15281
rect 19387 15244 19432 15272
rect 19420 15235 19432 15244
rect 19426 15232 19432 15235
rect 19484 15232 19490 15284
rect 25130 15232 25136 15284
rect 25188 15272 25194 15284
rect 25225 15275 25283 15281
rect 25225 15272 25237 15275
rect 25188 15244 25237 15272
rect 25188 15232 25194 15244
rect 25225 15241 25237 15244
rect 25271 15241 25283 15275
rect 25225 15235 25283 15241
rect 24302 15204 24308 15216
rect 24215 15176 24308 15204
rect 24302 15164 24308 15176
rect 24360 15204 24366 15216
rect 24762 15204 24768 15216
rect 24360 15176 24768 15204
rect 24360 15164 24366 15176
rect 24762 15164 24768 15176
rect 24820 15164 24826 15216
rect 23661 15139 23719 15145
rect 23661 15105 23673 15139
rect 23707 15136 23719 15139
rect 24118 15136 24124 15148
rect 23707 15108 24124 15136
rect 23707 15105 23719 15108
rect 23661 15099 23719 15105
rect 24118 15096 24124 15108
rect 24176 15096 24182 15148
rect 12989 15071 13047 15077
rect 12989 15037 13001 15071
rect 13035 15068 13047 15071
rect 13446 15068 13452 15080
rect 13035 15040 13452 15068
rect 13035 15037 13047 15040
rect 12989 15031 13047 15037
rect 13446 15028 13452 15040
rect 13504 15028 13510 15080
rect 15381 15071 15439 15077
rect 15381 15037 15393 15071
rect 15427 15068 15439 15071
rect 15838 15068 15844 15080
rect 15427 15040 15844 15068
rect 15427 15037 15439 15040
rect 15381 15031 15439 15037
rect 15838 15028 15844 15040
rect 15896 15028 15902 15080
rect 1104 14978 26864 15000
rect 1104 14926 5648 14978
rect 5700 14926 5712 14978
rect 5764 14926 5776 14978
rect 5828 14926 5840 14978
rect 5892 14926 14982 14978
rect 15034 14926 15046 14978
rect 15098 14926 15110 14978
rect 15162 14926 15174 14978
rect 15226 14926 24315 14978
rect 24367 14926 24379 14978
rect 24431 14926 24443 14978
rect 24495 14926 24507 14978
rect 24559 14926 26864 14978
rect 1104 14904 26864 14926
rect 12069 14867 12127 14873
rect 12069 14833 12081 14867
rect 12115 14864 12127 14867
rect 12434 14864 12440 14876
rect 12115 14836 12440 14864
rect 12115 14833 12127 14836
rect 12069 14827 12127 14833
rect 12434 14824 12440 14836
rect 12492 14864 12498 14876
rect 12897 14867 12955 14873
rect 12897 14864 12909 14867
rect 12492 14836 12909 14864
rect 12492 14824 12498 14836
rect 12897 14833 12909 14836
rect 12943 14833 12955 14867
rect 17218 14864 17224 14876
rect 17179 14836 17224 14864
rect 12897 14827 12955 14833
rect 17218 14824 17224 14836
rect 17276 14824 17282 14876
rect 19150 14864 19156 14876
rect 19111 14836 19156 14864
rect 19150 14824 19156 14836
rect 19208 14824 19214 14876
rect 19426 14824 19432 14876
rect 19484 14864 19490 14876
rect 19521 14867 19579 14873
rect 19521 14864 19533 14867
rect 19484 14836 19533 14864
rect 19484 14824 19490 14836
rect 19521 14833 19533 14836
rect 19567 14833 19579 14867
rect 19521 14827 19579 14833
rect 21453 14867 21511 14873
rect 21453 14833 21465 14867
rect 21499 14864 21511 14867
rect 21542 14864 21548 14876
rect 21499 14836 21548 14864
rect 21499 14833 21511 14836
rect 21453 14827 21511 14833
rect 21542 14824 21548 14836
rect 21600 14824 21606 14876
rect 23385 14867 23443 14873
rect 23385 14833 23397 14867
rect 23431 14864 23443 14867
rect 23566 14864 23572 14876
rect 23431 14836 23572 14864
rect 23431 14833 23443 14836
rect 23385 14827 23443 14833
rect 23566 14824 23572 14836
rect 23624 14824 23630 14876
rect 23661 14867 23719 14873
rect 23661 14833 23673 14867
rect 23707 14864 23719 14867
rect 24670 14864 24676 14876
rect 23707 14836 24676 14864
rect 23707 14833 23719 14836
rect 23661 14827 23719 14833
rect 24670 14824 24676 14836
rect 24728 14824 24734 14876
rect 25130 14824 25136 14876
rect 25188 14864 25194 14876
rect 25225 14867 25283 14873
rect 25225 14864 25237 14867
rect 25188 14836 25237 14864
rect 25188 14824 25194 14836
rect 25225 14833 25237 14836
rect 25271 14833 25283 14867
rect 25225 14827 25283 14833
rect 14369 14799 14427 14805
rect 14369 14765 14381 14799
rect 14415 14796 14427 14799
rect 14642 14796 14648 14808
rect 14415 14768 14648 14796
rect 14415 14765 14427 14768
rect 14369 14759 14427 14765
rect 14642 14756 14648 14768
rect 14700 14796 14706 14808
rect 15289 14799 15347 14805
rect 15289 14796 15301 14799
rect 14700 14768 15301 14796
rect 14700 14756 14706 14768
rect 15289 14765 15301 14768
rect 15335 14765 15347 14799
rect 24026 14796 24032 14808
rect 23987 14768 24032 14796
rect 15289 14759 15347 14765
rect 24026 14756 24032 14768
rect 24084 14756 24090 14808
rect 24210 14756 24216 14808
rect 24268 14796 24274 14808
rect 24765 14799 24823 14805
rect 24765 14796 24777 14799
rect 24268 14768 24777 14796
rect 24268 14756 24274 14768
rect 24765 14765 24777 14768
rect 24811 14765 24823 14799
rect 24765 14759 24823 14765
rect 13446 14728 13452 14740
rect 13407 14700 13452 14728
rect 13446 14688 13452 14700
rect 13504 14688 13510 14740
rect 15838 14728 15844 14740
rect 15799 14700 15844 14728
rect 15838 14688 15844 14700
rect 15896 14688 15902 14740
rect 23658 14688 23664 14740
rect 23716 14728 23722 14740
rect 25038 14728 25044 14740
rect 23716 14700 25044 14728
rect 23716 14688 23722 14700
rect 25038 14688 25044 14700
rect 25096 14688 25102 14740
rect 17037 14663 17095 14669
rect 17037 14629 17049 14663
rect 17083 14660 17095 14663
rect 18046 14660 18052 14672
rect 17083 14632 17632 14660
rect 18007 14632 18052 14660
rect 17083 14629 17095 14632
rect 17037 14623 17095 14629
rect 12710 14552 12716 14604
rect 12768 14592 12774 14604
rect 12805 14595 12863 14601
rect 12805 14592 12817 14595
rect 12768 14564 12817 14592
rect 12768 14552 12774 14564
rect 12805 14561 12817 14564
rect 12851 14592 12863 14595
rect 13265 14595 13323 14601
rect 13265 14592 13277 14595
rect 12851 14564 13277 14592
rect 12851 14561 12863 14564
rect 12805 14555 12863 14561
rect 13265 14561 13277 14564
rect 13311 14561 13323 14595
rect 13265 14555 13323 14561
rect 15105 14595 15163 14601
rect 15105 14561 15117 14595
rect 15151 14592 15163 14595
rect 15657 14595 15715 14601
rect 15657 14592 15669 14595
rect 15151 14564 15669 14592
rect 15151 14561 15163 14564
rect 15105 14555 15163 14561
rect 15657 14561 15669 14564
rect 15703 14592 15715 14595
rect 16206 14592 16212 14604
rect 15703 14564 16212 14592
rect 15703 14561 15715 14564
rect 15657 14555 15715 14561
rect 16206 14552 16212 14564
rect 16264 14552 16270 14604
rect 17604 14536 17632 14632
rect 18046 14620 18052 14632
rect 18104 14660 18110 14672
rect 18509 14663 18567 14669
rect 18509 14660 18521 14663
rect 18104 14632 18521 14660
rect 18104 14620 18110 14632
rect 18509 14629 18521 14632
rect 18555 14629 18567 14663
rect 18509 14623 18567 14629
rect 20990 14620 20996 14672
rect 21048 14660 21054 14672
rect 21269 14663 21327 14669
rect 21269 14660 21281 14663
rect 21048 14632 21281 14660
rect 21048 14620 21054 14632
rect 21269 14629 21281 14632
rect 21315 14660 21327 14663
rect 21729 14663 21787 14669
rect 21729 14660 21741 14663
rect 21315 14632 21741 14660
rect 21315 14629 21327 14632
rect 21269 14623 21327 14629
rect 21729 14629 21741 14632
rect 21775 14629 21787 14663
rect 23477 14663 23535 14669
rect 23477 14660 23489 14663
rect 21729 14623 21787 14629
rect 22940 14632 23489 14660
rect 22940 14604 22968 14632
rect 23477 14629 23489 14632
rect 23523 14629 23535 14663
rect 23477 14623 23535 14629
rect 23750 14620 23756 14672
rect 23808 14660 23814 14672
rect 24026 14660 24032 14672
rect 23808 14632 24032 14660
rect 23808 14620 23814 14632
rect 24026 14620 24032 14632
rect 24084 14620 24090 14672
rect 24581 14663 24639 14669
rect 24581 14629 24593 14663
rect 24627 14660 24639 14663
rect 24762 14660 24768 14672
rect 24627 14632 24768 14660
rect 24627 14629 24639 14632
rect 24581 14623 24639 14629
rect 24762 14620 24768 14632
rect 24820 14620 24826 14672
rect 22922 14592 22928 14604
rect 22883 14564 22928 14592
rect 22922 14552 22928 14564
rect 22980 14552 22986 14604
rect 26142 14592 26148 14604
rect 23768 14564 26148 14592
rect 23768 14536 23796 14564
rect 26142 14552 26148 14564
rect 26200 14552 26206 14604
rect 12437 14527 12495 14533
rect 12437 14493 12449 14527
rect 12483 14524 12495 14527
rect 12894 14524 12900 14536
rect 12483 14496 12900 14524
rect 12483 14493 12495 14496
rect 12437 14487 12495 14493
rect 12894 14484 12900 14496
rect 12952 14524 12958 14536
rect 13357 14527 13415 14533
rect 13357 14524 13369 14527
rect 12952 14496 13369 14524
rect 12952 14484 12958 14496
rect 13357 14493 13369 14496
rect 13403 14493 13415 14527
rect 13357 14487 13415 14493
rect 14737 14527 14795 14533
rect 14737 14493 14749 14527
rect 14783 14524 14795 14527
rect 15470 14524 15476 14536
rect 14783 14496 15476 14524
rect 14783 14493 14795 14496
rect 14737 14487 14795 14493
rect 15470 14484 15476 14496
rect 15528 14524 15534 14536
rect 15749 14527 15807 14533
rect 15749 14524 15761 14527
rect 15528 14496 15761 14524
rect 15528 14484 15534 14496
rect 15749 14493 15761 14496
rect 15795 14493 15807 14527
rect 17586 14524 17592 14536
rect 17547 14496 17592 14524
rect 15749 14487 15807 14493
rect 17586 14484 17592 14496
rect 17644 14484 17650 14536
rect 18230 14524 18236 14536
rect 18191 14496 18236 14524
rect 18230 14484 18236 14496
rect 18288 14484 18294 14536
rect 23750 14484 23756 14536
rect 23808 14484 23814 14536
rect 24486 14524 24492 14536
rect 24447 14496 24492 14524
rect 24486 14484 24492 14496
rect 24544 14524 24550 14536
rect 24854 14524 24860 14536
rect 24544 14496 24860 14524
rect 24544 14484 24550 14496
rect 24854 14484 24860 14496
rect 24912 14484 24918 14536
rect 1104 14434 26864 14456
rect 1104 14382 10315 14434
rect 10367 14382 10379 14434
rect 10431 14382 10443 14434
rect 10495 14382 10507 14434
rect 10559 14382 19648 14434
rect 19700 14382 19712 14434
rect 19764 14382 19776 14434
rect 19828 14382 19840 14434
rect 19892 14382 26864 14434
rect 1104 14360 26864 14382
rect 12710 14320 12716 14332
rect 12671 14292 12716 14320
rect 12710 14280 12716 14292
rect 12768 14280 12774 14332
rect 16206 14320 16212 14332
rect 16167 14292 16212 14320
rect 16206 14280 16212 14292
rect 16264 14280 16270 14332
rect 17586 14280 17592 14332
rect 17644 14320 17650 14332
rect 18049 14323 18107 14329
rect 18049 14320 18061 14323
rect 17644 14292 18061 14320
rect 17644 14280 17650 14292
rect 18049 14289 18061 14292
rect 18095 14289 18107 14323
rect 20990 14320 20996 14332
rect 20951 14292 20996 14320
rect 18049 14283 18107 14289
rect 20990 14280 20996 14292
rect 21048 14280 21054 14332
rect 24486 14280 24492 14332
rect 24544 14320 24550 14332
rect 25041 14323 25099 14329
rect 25041 14320 25053 14323
rect 24544 14292 25053 14320
rect 24544 14280 24550 14292
rect 25041 14289 25053 14292
rect 25087 14289 25099 14323
rect 25041 14283 25099 14289
rect 13446 14212 13452 14264
rect 13504 14252 13510 14264
rect 13970 14255 14028 14261
rect 13970 14252 13982 14255
rect 13504 14224 13982 14252
rect 13504 14212 13510 14224
rect 13970 14221 13982 14224
rect 14016 14221 14028 14255
rect 13970 14215 14028 14221
rect 23014 14212 23020 14264
rect 23072 14252 23078 14264
rect 23566 14252 23572 14264
rect 23072 14224 23572 14252
rect 23072 14212 23078 14224
rect 23566 14212 23572 14224
rect 23624 14252 23630 14264
rect 23906 14255 23964 14261
rect 23906 14252 23918 14255
rect 23624 14224 23918 14252
rect 23624 14212 23630 14224
rect 23906 14221 23918 14224
rect 23952 14221 23964 14255
rect 23906 14215 23964 14221
rect 13354 14144 13360 14196
rect 13412 14184 13418 14196
rect 13725 14187 13783 14193
rect 13725 14184 13737 14187
rect 13412 14156 13737 14184
rect 13412 14144 13418 14156
rect 13725 14153 13737 14156
rect 13771 14184 13783 14187
rect 14458 14184 14464 14196
rect 13771 14156 14464 14184
rect 13771 14153 13783 14156
rect 13725 14147 13783 14153
rect 14458 14144 14464 14156
rect 14516 14144 14522 14196
rect 18046 14144 18052 14196
rect 18104 14184 18110 14196
rect 18417 14187 18475 14193
rect 18417 14184 18429 14187
rect 18104 14156 18429 14184
rect 18104 14144 18110 14156
rect 18417 14153 18429 14156
rect 18463 14153 18475 14187
rect 21358 14184 21364 14196
rect 21319 14156 21364 14184
rect 18417 14147 18475 14153
rect 21358 14144 21364 14156
rect 21416 14144 21422 14196
rect 22094 14144 22100 14196
rect 22152 14184 22158 14196
rect 22557 14187 22615 14193
rect 22557 14184 22569 14187
rect 22152 14156 22569 14184
rect 22152 14144 22158 14156
rect 22557 14153 22569 14156
rect 22603 14184 22615 14187
rect 22922 14184 22928 14196
rect 22603 14156 22928 14184
rect 22603 14153 22615 14156
rect 22557 14147 22615 14153
rect 22922 14144 22928 14156
rect 22980 14144 22986 14196
rect 23106 14144 23112 14196
rect 23164 14184 23170 14196
rect 23661 14187 23719 14193
rect 23661 14184 23673 14187
rect 23164 14156 23673 14184
rect 23164 14144 23170 14156
rect 23661 14153 23673 14156
rect 23707 14153 23719 14187
rect 23661 14147 23719 14153
rect 18506 14116 18512 14128
rect 18467 14088 18512 14116
rect 18506 14076 18512 14088
rect 18564 14076 18570 14128
rect 18598 14076 18604 14128
rect 18656 14116 18662 14128
rect 21450 14116 21456 14128
rect 18656 14088 18701 14116
rect 21411 14088 21456 14116
rect 18656 14076 18662 14088
rect 21450 14076 21456 14088
rect 21508 14076 21514 14128
rect 21634 14076 21640 14128
rect 21692 14116 21698 14128
rect 21692 14088 21737 14116
rect 21692 14076 21698 14088
rect 22281 14051 22339 14057
rect 22281 14017 22293 14051
rect 22327 14048 22339 14051
rect 22370 14048 22376 14060
rect 22327 14020 22376 14048
rect 22327 14017 22339 14020
rect 22281 14011 22339 14017
rect 22370 14008 22376 14020
rect 22428 14008 22434 14060
rect 15105 13983 15163 13989
rect 15105 13949 15117 13983
rect 15151 13980 15163 13983
rect 15378 13980 15384 13992
rect 15151 13952 15384 13980
rect 15151 13949 15163 13952
rect 15105 13943 15163 13949
rect 15378 13940 15384 13952
rect 15436 13940 15442 13992
rect 22741 13983 22799 13989
rect 22741 13949 22753 13983
rect 22787 13980 22799 13983
rect 23474 13980 23480 13992
rect 22787 13952 23480 13980
rect 22787 13949 22799 13952
rect 22741 13943 22799 13949
rect 23474 13940 23480 13952
rect 23532 13940 23538 13992
rect 1104 13890 26864 13912
rect 1104 13838 5648 13890
rect 5700 13838 5712 13890
rect 5764 13838 5776 13890
rect 5828 13838 5840 13890
rect 5892 13838 14982 13890
rect 15034 13838 15046 13890
rect 15098 13838 15110 13890
rect 15162 13838 15174 13890
rect 15226 13838 24315 13890
rect 24367 13838 24379 13890
rect 24431 13838 24443 13890
rect 24495 13838 24507 13890
rect 24559 13838 26864 13890
rect 1104 13816 26864 13838
rect 12066 13736 12072 13788
rect 12124 13776 12130 13788
rect 13354 13776 13360 13788
rect 12124 13748 13360 13776
rect 12124 13736 12130 13748
rect 13354 13736 13360 13748
rect 13412 13736 13418 13788
rect 13446 13736 13452 13788
rect 13504 13776 13510 13788
rect 13633 13779 13691 13785
rect 13633 13776 13645 13779
rect 13504 13748 13645 13776
rect 13504 13736 13510 13748
rect 13633 13745 13645 13748
rect 13679 13776 13691 13779
rect 14553 13779 14611 13785
rect 14553 13776 14565 13779
rect 13679 13748 14565 13776
rect 13679 13745 13691 13748
rect 13633 13739 13691 13745
rect 14553 13745 14565 13748
rect 14599 13745 14611 13779
rect 14553 13739 14611 13745
rect 15930 13736 15936 13788
rect 15988 13776 15994 13788
rect 16669 13779 16727 13785
rect 16669 13776 16681 13779
rect 15988 13748 16681 13776
rect 15988 13736 15994 13748
rect 16669 13745 16681 13748
rect 16715 13745 16727 13779
rect 16669 13739 16727 13745
rect 17313 13779 17371 13785
rect 17313 13745 17325 13779
rect 17359 13776 17371 13779
rect 18046 13776 18052 13788
rect 17359 13748 18052 13776
rect 17359 13745 17371 13748
rect 17313 13739 17371 13745
rect 14277 13711 14335 13717
rect 14277 13677 14289 13711
rect 14323 13708 14335 13711
rect 14458 13708 14464 13720
rect 14323 13680 14464 13708
rect 14323 13677 14335 13680
rect 14277 13671 14335 13677
rect 14458 13668 14464 13680
rect 14516 13708 14522 13720
rect 15013 13711 15071 13717
rect 15013 13708 15025 13711
rect 14516 13680 15025 13708
rect 14516 13668 14522 13680
rect 15013 13677 15025 13680
rect 15059 13708 15071 13711
rect 15059 13680 15332 13708
rect 15059 13677 15071 13680
rect 15013 13671 15071 13677
rect 15304 13649 15332 13680
rect 15289 13643 15347 13649
rect 11716 13612 12388 13640
rect 11716 13584 11744 13612
rect 11698 13572 11704 13584
rect 11659 13544 11704 13572
rect 11698 13532 11704 13544
rect 11756 13532 11762 13584
rect 12066 13572 12072 13584
rect 12027 13544 12072 13572
rect 12066 13532 12072 13544
rect 12124 13572 12130 13584
rect 12253 13575 12311 13581
rect 12253 13572 12265 13575
rect 12124 13544 12265 13572
rect 12124 13532 12130 13544
rect 12253 13541 12265 13544
rect 12299 13541 12311 13575
rect 12360 13572 12388 13612
rect 15289 13609 15301 13643
rect 15335 13609 15347 13643
rect 16684 13640 16712 13739
rect 18046 13736 18052 13748
rect 18104 13736 18110 13788
rect 21358 13736 21364 13788
rect 21416 13776 21422 13788
rect 21637 13779 21695 13785
rect 21637 13776 21649 13779
rect 21416 13748 21649 13776
rect 21416 13736 21422 13748
rect 21637 13745 21649 13748
rect 21683 13745 21695 13779
rect 21637 13739 21695 13745
rect 22097 13779 22155 13785
rect 22097 13745 22109 13779
rect 22143 13776 22155 13779
rect 23106 13776 23112 13788
rect 22143 13748 23112 13776
rect 22143 13745 22155 13748
rect 22097 13739 22155 13745
rect 17678 13708 17684 13720
rect 17639 13680 17684 13708
rect 17678 13668 17684 13680
rect 17736 13668 17742 13720
rect 21177 13643 21235 13649
rect 16684 13612 17908 13640
rect 15289 13603 15347 13609
rect 17880 13584 17908 13612
rect 21177 13609 21189 13643
rect 21223 13640 21235 13643
rect 21376 13640 21404 13736
rect 22204 13649 22232 13748
rect 23106 13736 23112 13748
rect 23164 13776 23170 13788
rect 24121 13779 24179 13785
rect 24121 13776 24133 13779
rect 23164 13748 24133 13776
rect 23164 13736 23170 13748
rect 24121 13745 24133 13748
rect 24167 13745 24179 13779
rect 24854 13776 24860 13788
rect 24815 13748 24860 13776
rect 24121 13739 24179 13745
rect 24854 13736 24860 13748
rect 24912 13736 24918 13788
rect 23566 13708 23572 13720
rect 23527 13680 23572 13708
rect 23566 13668 23572 13680
rect 23624 13708 23630 13720
rect 24489 13711 24547 13717
rect 24489 13708 24501 13711
rect 23624 13680 24501 13708
rect 23624 13668 23630 13680
rect 24489 13677 24501 13680
rect 24535 13677 24547 13711
rect 24489 13671 24547 13677
rect 21223 13612 21404 13640
rect 22189 13643 22247 13649
rect 21223 13609 21235 13612
rect 21177 13603 21235 13609
rect 22189 13609 22201 13643
rect 22235 13609 22247 13643
rect 22189 13603 22247 13609
rect 12520 13575 12578 13581
rect 12520 13572 12532 13575
rect 12360 13544 12532 13572
rect 12253 13535 12311 13541
rect 12520 13541 12532 13544
rect 12566 13572 12578 13575
rect 13630 13572 13636 13584
rect 12566 13544 13636 13572
rect 12566 13541 12578 13544
rect 12520 13535 12578 13541
rect 13630 13532 13636 13544
rect 13688 13532 13694 13584
rect 15378 13532 15384 13584
rect 15436 13572 15442 13584
rect 15545 13575 15603 13581
rect 15545 13572 15557 13575
rect 15436 13544 15557 13572
rect 15436 13532 15442 13544
rect 15545 13541 15557 13544
rect 15591 13541 15603 13575
rect 15545 13535 15603 13541
rect 17678 13532 17684 13584
rect 17736 13572 17742 13584
rect 17773 13575 17831 13581
rect 17773 13572 17785 13575
rect 17736 13544 17785 13572
rect 17736 13532 17742 13544
rect 17773 13541 17785 13544
rect 17819 13541 17831 13575
rect 17773 13535 17831 13541
rect 17862 13532 17868 13584
rect 17920 13572 17926 13584
rect 18029 13575 18087 13581
rect 18029 13572 18041 13575
rect 17920 13544 18041 13572
rect 17920 13532 17926 13544
rect 18029 13541 18041 13544
rect 18075 13541 18087 13575
rect 18029 13535 18087 13541
rect 20349 13575 20407 13581
rect 20349 13541 20361 13575
rect 20395 13572 20407 13575
rect 21450 13572 21456 13584
rect 20395 13544 21456 13572
rect 20395 13541 20407 13544
rect 20349 13535 20407 13541
rect 21450 13532 21456 13544
rect 21508 13532 21514 13584
rect 24578 13532 24584 13584
rect 24636 13572 24642 13584
rect 24673 13575 24731 13581
rect 24673 13572 24685 13575
rect 24636 13544 24685 13572
rect 24636 13532 24642 13544
rect 24673 13541 24685 13544
rect 24719 13572 24731 13575
rect 25225 13575 25283 13581
rect 25225 13572 25237 13575
rect 24719 13544 25237 13572
rect 24719 13541 24731 13544
rect 24673 13535 24731 13541
rect 25225 13541 25237 13544
rect 25271 13541 25283 13575
rect 25225 13535 25283 13541
rect 20717 13507 20775 13513
rect 20717 13473 20729 13507
rect 20763 13504 20775 13507
rect 21634 13504 21640 13516
rect 20763 13476 21640 13504
rect 20763 13473 20775 13476
rect 20717 13467 20775 13473
rect 21634 13464 21640 13476
rect 21692 13504 21698 13516
rect 22370 13504 22376 13516
rect 21692 13476 22376 13504
rect 21692 13464 21698 13476
rect 22370 13464 22376 13476
rect 22428 13513 22434 13516
rect 22428 13507 22492 13513
rect 22428 13473 22446 13507
rect 22480 13473 22492 13507
rect 22428 13467 22492 13473
rect 22428 13464 22434 13467
rect 19150 13436 19156 13448
rect 19111 13408 19156 13436
rect 19150 13396 19156 13408
rect 19208 13396 19214 13448
rect 1104 13346 26864 13368
rect 1104 13294 10315 13346
rect 10367 13294 10379 13346
rect 10431 13294 10443 13346
rect 10495 13294 10507 13346
rect 10559 13294 19648 13346
rect 19700 13294 19712 13346
rect 19764 13294 19776 13346
rect 19828 13294 19840 13346
rect 19892 13294 26864 13346
rect 1104 13272 26864 13294
rect 2774 13232 2780 13244
rect 2735 13204 2780 13232
rect 2774 13192 2780 13204
rect 2832 13192 2838 13244
rect 12894 13232 12900 13244
rect 12855 13204 12900 13232
rect 12894 13192 12900 13204
rect 12952 13192 12958 13244
rect 15470 13232 15476 13244
rect 15431 13204 15476 13232
rect 15470 13192 15476 13204
rect 15528 13192 15534 13244
rect 17862 13232 17868 13244
rect 17823 13204 17868 13232
rect 17862 13192 17868 13204
rect 17920 13192 17926 13244
rect 18046 13232 18052 13244
rect 18007 13204 18052 13232
rect 18046 13192 18052 13204
rect 18104 13192 18110 13244
rect 18506 13192 18512 13244
rect 18564 13232 18570 13244
rect 18690 13232 18696 13244
rect 18564 13204 18696 13232
rect 18564 13192 18570 13204
rect 18690 13192 18696 13204
rect 18748 13232 18754 13244
rect 18877 13235 18935 13241
rect 18877 13232 18889 13235
rect 18748 13204 18889 13232
rect 18748 13192 18754 13204
rect 18877 13201 18889 13204
rect 18923 13201 18935 13235
rect 18877 13195 18935 13201
rect 21450 13192 21456 13244
rect 21508 13232 21514 13244
rect 21913 13235 21971 13241
rect 21913 13232 21925 13235
rect 21508 13204 21925 13232
rect 21508 13192 21514 13204
rect 21913 13201 21925 13204
rect 21959 13201 21971 13235
rect 22922 13232 22928 13244
rect 22883 13204 22928 13232
rect 21913 13195 21971 13201
rect 22922 13192 22928 13204
rect 22980 13192 22986 13244
rect 24762 13232 24768 13244
rect 24723 13204 24768 13232
rect 24762 13192 24768 13204
rect 24820 13192 24826 13244
rect 2038 13164 2044 13176
rect 1412 13136 2044 13164
rect 1412 13105 1440 13136
rect 2038 13124 2044 13136
rect 2096 13124 2102 13176
rect 15378 13164 15384 13176
rect 15339 13136 15384 13164
rect 15378 13124 15384 13136
rect 15436 13164 15442 13176
rect 18598 13164 18604 13176
rect 15436 13136 16068 13164
rect 18559 13136 18604 13164
rect 15436 13124 15442 13136
rect 1397 13099 1455 13105
rect 1397 13065 1409 13099
rect 1443 13065 1455 13099
rect 1397 13059 1455 13065
rect 1486 13056 1492 13108
rect 1544 13096 1550 13108
rect 1653 13099 1711 13105
rect 1653 13096 1665 13099
rect 1544 13068 1665 13096
rect 1544 13056 1550 13068
rect 1653 13065 1665 13068
rect 1699 13065 1711 13099
rect 13262 13096 13268 13108
rect 13223 13068 13268 13096
rect 1653 13059 1711 13065
rect 13262 13056 13268 13068
rect 13320 13056 13326 13108
rect 15838 13096 15844 13108
rect 15799 13068 15844 13096
rect 15838 13056 15844 13068
rect 15896 13056 15902 13108
rect 13354 13028 13360 13040
rect 13315 13000 13360 13028
rect 13354 12988 13360 13000
rect 13412 12988 13418 13040
rect 13541 13031 13599 13037
rect 13541 12997 13553 13031
rect 13587 13028 13599 13031
rect 13630 13028 13636 13040
rect 13587 13000 13636 13028
rect 13587 12997 13599 13000
rect 13541 12991 13599 12997
rect 13630 12988 13636 13000
rect 13688 12988 13694 13040
rect 15930 13028 15936 13040
rect 15891 13000 15936 13028
rect 15930 12988 15936 13000
rect 15988 12988 15994 13040
rect 16040 13037 16068 13136
rect 18598 13124 18604 13136
rect 18656 13164 18662 13176
rect 19426 13164 19432 13176
rect 18656 13136 19432 13164
rect 18656 13124 18662 13136
rect 19426 13124 19432 13136
rect 19484 13164 19490 13176
rect 19674 13167 19732 13173
rect 19674 13164 19686 13167
rect 19484 13136 19686 13164
rect 19484 13124 19490 13136
rect 19674 13133 19686 13136
rect 19720 13133 19732 13167
rect 19674 13127 19732 13133
rect 22186 13056 22192 13108
rect 22244 13096 22250 13108
rect 22281 13099 22339 13105
rect 22281 13096 22293 13099
rect 22244 13068 22293 13096
rect 22244 13056 22250 13068
rect 22281 13065 22293 13068
rect 22327 13065 22339 13099
rect 24578 13096 24584 13108
rect 24539 13068 24584 13096
rect 22281 13059 22339 13065
rect 24578 13056 24584 13068
rect 24636 13056 24642 13108
rect 16025 13031 16083 13037
rect 16025 12997 16037 13031
rect 16071 13028 16083 13031
rect 16206 13028 16212 13040
rect 16071 13000 16212 13028
rect 16071 12997 16083 13000
rect 16025 12991 16083 12997
rect 16206 12988 16212 13000
rect 16264 12988 16270 13040
rect 19242 12988 19248 13040
rect 19300 13028 19306 13040
rect 19429 13031 19487 13037
rect 19429 13028 19441 13031
rect 19300 13000 19441 13028
rect 19300 12988 19306 13000
rect 19429 12997 19441 13000
rect 19475 12997 19487 13031
rect 22373 13031 22431 13037
rect 22373 13028 22385 13031
rect 19429 12991 19487 12997
rect 22296 13000 22385 13028
rect 22296 12972 22324 13000
rect 22373 12997 22385 13000
rect 22419 12997 22431 13031
rect 22373 12991 22431 12997
rect 22462 12988 22468 13040
rect 22520 13028 22526 13040
rect 22520 13000 22565 13028
rect 22520 12988 22526 13000
rect 22278 12920 22284 12972
rect 22336 12920 22342 12972
rect 20806 12892 20812 12904
rect 20767 12864 20812 12892
rect 20806 12852 20812 12864
rect 20864 12852 20870 12904
rect 1104 12802 26864 12824
rect 1104 12750 5648 12802
rect 5700 12750 5712 12802
rect 5764 12750 5776 12802
rect 5828 12750 5840 12802
rect 5892 12750 14982 12802
rect 15034 12750 15046 12802
rect 15098 12750 15110 12802
rect 15162 12750 15174 12802
rect 15226 12750 24315 12802
rect 24367 12750 24379 12802
rect 24431 12750 24443 12802
rect 24495 12750 24507 12802
rect 24559 12750 26864 12802
rect 1104 12728 26864 12750
rect 1486 12648 1492 12700
rect 1544 12688 1550 12700
rect 1581 12691 1639 12697
rect 1581 12688 1593 12691
rect 1544 12660 1593 12688
rect 1544 12648 1550 12660
rect 1581 12657 1593 12660
rect 1627 12657 1639 12691
rect 2038 12688 2044 12700
rect 1999 12660 2044 12688
rect 1581 12651 1639 12657
rect 2038 12648 2044 12660
rect 2096 12648 2102 12700
rect 12989 12691 13047 12697
rect 12989 12657 13001 12691
rect 13035 12688 13047 12691
rect 13262 12688 13268 12700
rect 13035 12660 13268 12688
rect 13035 12657 13047 12660
rect 12989 12651 13047 12657
rect 13262 12648 13268 12660
rect 13320 12648 13326 12700
rect 13630 12688 13636 12700
rect 13591 12660 13636 12688
rect 13630 12648 13636 12660
rect 13688 12648 13694 12700
rect 15565 12691 15623 12697
rect 15565 12657 15577 12691
rect 15611 12688 15623 12691
rect 15838 12688 15844 12700
rect 15611 12660 15844 12688
rect 15611 12657 15623 12660
rect 15565 12651 15623 12657
rect 15838 12648 15844 12660
rect 15896 12648 15902 12700
rect 16206 12688 16212 12700
rect 16167 12660 16212 12688
rect 16206 12648 16212 12660
rect 16264 12648 16270 12700
rect 17957 12691 18015 12697
rect 17957 12657 17969 12691
rect 18003 12688 18015 12691
rect 18046 12688 18052 12700
rect 18003 12660 18052 12688
rect 18003 12657 18015 12660
rect 17957 12651 18015 12657
rect 18046 12648 18052 12660
rect 18104 12688 18110 12700
rect 19242 12688 19248 12700
rect 18104 12660 19248 12688
rect 18104 12648 18110 12660
rect 19242 12648 19248 12660
rect 19300 12648 19306 12700
rect 19426 12688 19432 12700
rect 19387 12660 19432 12688
rect 19426 12648 19432 12660
rect 19484 12648 19490 12700
rect 22281 12691 22339 12697
rect 22281 12657 22293 12691
rect 22327 12688 22339 12691
rect 22370 12688 22376 12700
rect 22327 12660 22376 12688
rect 22327 12657 22339 12660
rect 22281 12651 22339 12657
rect 22370 12648 22376 12660
rect 22428 12648 22434 12700
rect 23658 12688 23664 12700
rect 23619 12660 23664 12688
rect 23658 12648 23664 12660
rect 23716 12648 23722 12700
rect 24489 12691 24547 12697
rect 24489 12657 24501 12691
rect 24535 12688 24547 12691
rect 24670 12688 24676 12700
rect 24535 12660 24676 12688
rect 24535 12657 24547 12660
rect 24489 12651 24547 12657
rect 24670 12648 24676 12660
rect 24728 12648 24734 12700
rect 19260 12620 19288 12648
rect 19981 12623 20039 12629
rect 19981 12620 19993 12623
rect 19260 12592 19993 12620
rect 19981 12589 19993 12592
rect 20027 12620 20039 12623
rect 20625 12623 20683 12629
rect 20625 12620 20637 12623
rect 20027 12592 20637 12620
rect 20027 12589 20039 12592
rect 19981 12583 20039 12589
rect 20625 12589 20637 12592
rect 20671 12620 20683 12623
rect 24762 12620 24768 12632
rect 20671 12592 20944 12620
rect 24723 12592 24768 12620
rect 20671 12589 20683 12592
rect 20625 12583 20683 12589
rect 20916 12561 20944 12592
rect 24762 12580 24768 12592
rect 24820 12580 24826 12632
rect 17589 12555 17647 12561
rect 17589 12521 17601 12555
rect 17635 12552 17647 12555
rect 20901 12555 20959 12561
rect 17635 12524 18184 12552
rect 17635 12521 17647 12524
rect 17589 12515 17647 12521
rect 13354 12484 13360 12496
rect 13315 12456 13360 12484
rect 13354 12444 13360 12456
rect 13412 12444 13418 12496
rect 15930 12484 15936 12496
rect 15891 12456 15936 12484
rect 15930 12444 15936 12456
rect 15988 12444 15994 12496
rect 18046 12484 18052 12496
rect 18007 12456 18052 12484
rect 18046 12444 18052 12456
rect 18104 12444 18110 12496
rect 18156 12484 18184 12524
rect 20901 12521 20913 12555
rect 20947 12521 20959 12555
rect 20901 12515 20959 12521
rect 18316 12487 18374 12493
rect 18316 12484 18328 12487
rect 18156 12456 18328 12484
rect 18316 12453 18328 12456
rect 18362 12484 18374 12487
rect 19150 12484 19156 12496
rect 18362 12456 19156 12484
rect 18362 12453 18374 12456
rect 18316 12447 18374 12453
rect 19150 12444 19156 12456
rect 19208 12444 19214 12496
rect 20806 12444 20812 12496
rect 20864 12484 20870 12496
rect 21157 12487 21215 12493
rect 21157 12484 21169 12487
rect 20864 12456 21169 12484
rect 20864 12444 20870 12456
rect 21157 12453 21169 12456
rect 21203 12484 21215 12487
rect 22462 12484 22468 12496
rect 21203 12456 22468 12484
rect 21203 12453 21215 12456
rect 21157 12447 21215 12453
rect 22462 12444 22468 12456
rect 22520 12484 22526 12496
rect 22833 12487 22891 12493
rect 22833 12484 22845 12487
rect 22520 12456 22845 12484
rect 22520 12444 22526 12456
rect 22833 12453 22845 12456
rect 22879 12453 22891 12487
rect 23474 12484 23480 12496
rect 23435 12456 23480 12484
rect 22833 12447 22891 12453
rect 23474 12444 23480 12456
rect 23532 12484 23538 12496
rect 24029 12487 24087 12493
rect 24029 12484 24041 12487
rect 23532 12456 24041 12484
rect 23532 12444 23538 12456
rect 24029 12453 24041 12456
rect 24075 12453 24087 12487
rect 24029 12447 24087 12453
rect 24581 12487 24639 12493
rect 24581 12453 24593 12487
rect 24627 12453 24639 12487
rect 24581 12447 24639 12453
rect 24596 12416 24624 12447
rect 25133 12419 25191 12425
rect 25133 12416 25145 12419
rect 23492 12388 25145 12416
rect 23492 12360 23520 12388
rect 25133 12385 25145 12388
rect 25179 12385 25191 12419
rect 25133 12379 25191 12385
rect 23474 12308 23480 12360
rect 23532 12308 23538 12360
rect 1104 12258 26864 12280
rect 1104 12206 10315 12258
rect 10367 12206 10379 12258
rect 10431 12206 10443 12258
rect 10495 12206 10507 12258
rect 10559 12206 19648 12258
rect 19700 12206 19712 12258
rect 19764 12206 19776 12258
rect 19828 12206 19840 12258
rect 19892 12206 26864 12258
rect 1104 12184 26864 12206
rect 18233 12147 18291 12153
rect 18233 12113 18245 12147
rect 18279 12144 18291 12147
rect 18690 12144 18696 12156
rect 18279 12116 18696 12144
rect 18279 12113 18291 12116
rect 18233 12107 18291 12113
rect 18690 12104 18696 12116
rect 18748 12104 18754 12156
rect 19426 12144 19432 12156
rect 19387 12116 19432 12144
rect 19426 12104 19432 12116
rect 19484 12104 19490 12156
rect 20806 12104 20812 12156
rect 20864 12144 20870 12156
rect 20901 12147 20959 12153
rect 20901 12144 20913 12147
rect 20864 12116 20913 12144
rect 20864 12104 20870 12116
rect 20901 12113 20913 12116
rect 20947 12113 20959 12147
rect 22278 12144 22284 12156
rect 22239 12116 22284 12144
rect 20901 12107 20959 12113
rect 22278 12104 22284 12116
rect 22336 12104 22342 12156
rect 22741 12147 22799 12153
rect 22741 12113 22753 12147
rect 22787 12144 22799 12147
rect 23474 12144 23480 12156
rect 22787 12116 23480 12144
rect 22787 12113 22799 12116
rect 22741 12107 22799 12113
rect 23474 12104 23480 12116
rect 23532 12104 23538 12156
rect 24762 12144 24768 12156
rect 24723 12116 24768 12144
rect 24762 12104 24768 12116
rect 24820 12104 24826 12156
rect 18322 11968 18328 12020
rect 18380 12008 18386 12020
rect 18601 12011 18659 12017
rect 18601 12008 18613 12011
rect 18380 11980 18613 12008
rect 18380 11968 18386 11980
rect 18601 11977 18613 11980
rect 18647 11977 18659 12011
rect 18601 11971 18659 11977
rect 22094 11968 22100 12020
rect 22152 12008 22158 12020
rect 22554 12008 22560 12020
rect 22152 11980 22560 12008
rect 22152 11968 22158 11980
rect 22554 11968 22560 11980
rect 22612 11968 22618 12020
rect 24581 12011 24639 12017
rect 24581 11977 24593 12011
rect 24627 12008 24639 12011
rect 24670 12008 24676 12020
rect 24627 11980 24676 12008
rect 24627 11977 24639 11980
rect 24581 11971 24639 11977
rect 24670 11968 24676 11980
rect 24728 11968 24734 12020
rect 18506 11900 18512 11952
rect 18564 11940 18570 11952
rect 18693 11943 18751 11949
rect 18693 11940 18705 11943
rect 18564 11912 18705 11940
rect 18564 11900 18570 11912
rect 18693 11909 18705 11912
rect 18739 11909 18751 11943
rect 18693 11903 18751 11909
rect 18877 11943 18935 11949
rect 18877 11909 18889 11943
rect 18923 11940 18935 11943
rect 19150 11940 19156 11952
rect 18923 11912 19156 11940
rect 18923 11909 18935 11912
rect 18877 11903 18935 11909
rect 19150 11900 19156 11912
rect 19208 11900 19214 11952
rect 22002 11940 22008 11952
rect 21963 11912 22008 11940
rect 22002 11900 22008 11912
rect 22060 11900 22066 11952
rect 1104 11714 26864 11736
rect 1104 11662 5648 11714
rect 5700 11662 5712 11714
rect 5764 11662 5776 11714
rect 5828 11662 5840 11714
rect 5892 11662 14982 11714
rect 15034 11662 15046 11714
rect 15098 11662 15110 11714
rect 15162 11662 15174 11714
rect 15226 11662 24315 11714
rect 24367 11662 24379 11714
rect 24431 11662 24443 11714
rect 24495 11662 24507 11714
rect 24559 11662 26864 11714
rect 1104 11640 26864 11662
rect 18506 11560 18512 11612
rect 18564 11600 18570 11612
rect 18601 11603 18659 11609
rect 18601 11600 18613 11603
rect 18564 11572 18613 11600
rect 18564 11560 18570 11572
rect 18601 11569 18613 11572
rect 18647 11569 18659 11603
rect 18601 11563 18659 11569
rect 19061 11603 19119 11609
rect 19061 11569 19073 11603
rect 19107 11600 19119 11603
rect 19150 11600 19156 11612
rect 19107 11572 19156 11600
rect 19107 11569 19119 11572
rect 19061 11563 19119 11569
rect 19150 11560 19156 11572
rect 19208 11560 19214 11612
rect 22554 11600 22560 11612
rect 22515 11572 22560 11600
rect 22554 11560 22560 11572
rect 22612 11560 22618 11612
rect 23753 11603 23811 11609
rect 23753 11569 23765 11603
rect 23799 11600 23811 11603
rect 24489 11603 24547 11609
rect 24489 11600 24501 11603
rect 23799 11572 24501 11600
rect 23799 11569 23811 11572
rect 23753 11563 23811 11569
rect 24489 11569 24501 11572
rect 24535 11600 24547 11603
rect 24670 11600 24676 11612
rect 24535 11572 24676 11600
rect 24535 11569 24547 11572
rect 24489 11563 24547 11569
rect 24670 11560 24676 11572
rect 24728 11560 24734 11612
rect 24762 11560 24768 11612
rect 24820 11600 24826 11612
rect 24820 11572 24865 11600
rect 24820 11560 24826 11572
rect 23842 11492 23848 11544
rect 23900 11532 23906 11544
rect 24029 11535 24087 11541
rect 24029 11532 24041 11535
rect 23900 11504 24041 11532
rect 23900 11492 23906 11504
rect 24029 11501 24041 11504
rect 24075 11501 24087 11535
rect 24029 11495 24087 11501
rect 23569 11399 23627 11405
rect 23569 11365 23581 11399
rect 23615 11396 23627 11399
rect 23860 11396 23888 11492
rect 25222 11464 25228 11476
rect 24596 11436 25228 11464
rect 24596 11405 24624 11436
rect 25222 11424 25228 11436
rect 25280 11424 25286 11476
rect 23615 11368 23888 11396
rect 24581 11399 24639 11405
rect 23615 11365 23627 11368
rect 23569 11359 23627 11365
rect 24581 11365 24593 11399
rect 24627 11365 24639 11399
rect 24581 11359 24639 11365
rect 18322 11260 18328 11272
rect 18283 11232 18328 11260
rect 18322 11220 18328 11232
rect 18380 11220 18386 11272
rect 1104 11170 26864 11192
rect 1104 11118 10315 11170
rect 10367 11118 10379 11170
rect 10431 11118 10443 11170
rect 10495 11118 10507 11170
rect 10559 11118 19648 11170
rect 19700 11118 19712 11170
rect 19764 11118 19776 11170
rect 19828 11118 19840 11170
rect 19892 11118 26864 11170
rect 1104 11096 26864 11118
rect 23750 11016 23756 11068
rect 23808 11056 23814 11068
rect 24765 11059 24823 11065
rect 24765 11056 24777 11059
rect 23808 11028 24777 11056
rect 23808 11016 23814 11028
rect 24765 11025 24777 11028
rect 24811 11025 24823 11059
rect 24765 11019 24823 11025
rect 24578 10920 24584 10932
rect 24539 10892 24584 10920
rect 24578 10880 24584 10892
rect 24636 10880 24642 10932
rect 1104 10626 26864 10648
rect 1104 10574 5648 10626
rect 5700 10574 5712 10626
rect 5764 10574 5776 10626
rect 5828 10574 5840 10626
rect 5892 10574 14982 10626
rect 15034 10574 15046 10626
rect 15098 10574 15110 10626
rect 15162 10574 15174 10626
rect 15226 10574 24315 10626
rect 24367 10574 24379 10626
rect 24431 10574 24443 10626
rect 24495 10574 24507 10626
rect 24559 10574 26864 10626
rect 1104 10552 26864 10574
rect 24762 10512 24768 10524
rect 24723 10484 24768 10512
rect 24762 10472 24768 10484
rect 24820 10472 24826 10524
rect 24489 10447 24547 10453
rect 24489 10413 24501 10447
rect 24535 10444 24547 10447
rect 24670 10444 24676 10456
rect 24535 10416 24676 10444
rect 24535 10413 24547 10416
rect 24489 10407 24547 10413
rect 24670 10404 24676 10416
rect 24728 10404 24734 10456
rect 24581 10311 24639 10317
rect 24581 10277 24593 10311
rect 24627 10277 24639 10311
rect 24581 10271 24639 10277
rect 24596 10240 24624 10271
rect 25222 10240 25228 10252
rect 24596 10212 25228 10240
rect 25222 10200 25228 10212
rect 25280 10200 25286 10252
rect 1104 10082 26864 10104
rect 1104 10030 10315 10082
rect 10367 10030 10379 10082
rect 10431 10030 10443 10082
rect 10495 10030 10507 10082
rect 10559 10030 19648 10082
rect 19700 10030 19712 10082
rect 19764 10030 19776 10082
rect 19828 10030 19840 10082
rect 19892 10030 26864 10082
rect 1104 10008 26864 10030
rect 24026 9928 24032 9980
rect 24084 9968 24090 9980
rect 24765 9971 24823 9977
rect 24765 9968 24777 9971
rect 24084 9940 24777 9968
rect 24084 9928 24090 9940
rect 24765 9937 24777 9940
rect 24811 9937 24823 9971
rect 24765 9931 24823 9937
rect 24578 9832 24584 9844
rect 24539 9804 24584 9832
rect 24578 9792 24584 9804
rect 24636 9792 24642 9844
rect 1104 9538 26864 9560
rect 1104 9486 5648 9538
rect 5700 9486 5712 9538
rect 5764 9486 5776 9538
rect 5828 9486 5840 9538
rect 5892 9486 14982 9538
rect 15034 9486 15046 9538
rect 15098 9486 15110 9538
rect 15162 9486 15174 9538
rect 15226 9486 24315 9538
rect 24367 9486 24379 9538
rect 24431 9486 24443 9538
rect 24495 9486 24507 9538
rect 24559 9486 26864 9538
rect 1104 9464 26864 9486
rect 18230 9384 18236 9436
rect 18288 9424 18294 9436
rect 18966 9424 18972 9436
rect 18288 9396 18972 9424
rect 18288 9384 18294 9396
rect 18966 9384 18972 9396
rect 19024 9384 19030 9436
rect 24670 9424 24676 9436
rect 24631 9396 24676 9424
rect 24670 9384 24676 9396
rect 24728 9384 24734 9436
rect 23934 9356 23940 9368
rect 23895 9328 23940 9356
rect 23934 9316 23940 9328
rect 23992 9316 23998 9368
rect 23753 9223 23811 9229
rect 23753 9189 23765 9223
rect 23799 9189 23811 9223
rect 23753 9183 23811 9189
rect 23768 9152 23796 9183
rect 24394 9152 24400 9164
rect 23768 9124 24400 9152
rect 24394 9112 24400 9124
rect 24452 9112 24458 9164
rect 1104 8994 26864 9016
rect 1104 8942 10315 8994
rect 10367 8942 10379 8994
rect 10431 8942 10443 8994
rect 10495 8942 10507 8994
rect 10559 8942 19648 8994
rect 19700 8942 19712 8994
rect 19764 8942 19776 8994
rect 19828 8942 19840 8994
rect 19892 8942 26864 8994
rect 1104 8920 26864 8942
rect 24118 8840 24124 8892
rect 24176 8880 24182 8892
rect 24581 8883 24639 8889
rect 24581 8880 24593 8883
rect 24176 8852 24593 8880
rect 24176 8840 24182 8852
rect 24581 8849 24593 8852
rect 24627 8849 24639 8883
rect 24581 8843 24639 8849
rect 24394 8744 24400 8756
rect 24355 8716 24400 8744
rect 24394 8704 24400 8716
rect 24452 8704 24458 8756
rect 16482 8636 16488 8688
rect 16540 8676 16546 8688
rect 16666 8676 16672 8688
rect 16540 8648 16672 8676
rect 16540 8636 16546 8648
rect 16666 8636 16672 8648
rect 16724 8636 16730 8688
rect 1104 8450 26864 8472
rect 1104 8398 5648 8450
rect 5700 8398 5712 8450
rect 5764 8398 5776 8450
rect 5828 8398 5840 8450
rect 5892 8398 14982 8450
rect 15034 8398 15046 8450
rect 15098 8398 15110 8450
rect 15162 8398 15174 8450
rect 15226 8398 24315 8450
rect 24367 8398 24379 8450
rect 24431 8398 24443 8450
rect 24495 8398 24507 8450
rect 24559 8398 26864 8450
rect 1104 8376 26864 8398
rect 24489 8339 24547 8345
rect 24489 8305 24501 8339
rect 24535 8336 24547 8339
rect 24670 8336 24676 8348
rect 24535 8308 24676 8336
rect 24535 8305 24547 8308
rect 24489 8299 24547 8305
rect 24670 8296 24676 8308
rect 24728 8296 24734 8348
rect 1104 7906 26864 7928
rect 1104 7854 10315 7906
rect 10367 7854 10379 7906
rect 10431 7854 10443 7906
rect 10495 7854 10507 7906
rect 10559 7854 19648 7906
rect 19700 7854 19712 7906
rect 19764 7854 19776 7906
rect 19828 7854 19840 7906
rect 19892 7854 26864 7906
rect 1104 7832 26864 7854
rect 23474 7752 23480 7804
rect 23532 7792 23538 7804
rect 24765 7795 24823 7801
rect 24765 7792 24777 7795
rect 23532 7764 24777 7792
rect 23532 7752 23538 7764
rect 24765 7761 24777 7764
rect 24811 7761 24823 7795
rect 24765 7755 24823 7761
rect 24581 7659 24639 7665
rect 24581 7625 24593 7659
rect 24627 7656 24639 7659
rect 24670 7656 24676 7668
rect 24627 7628 24676 7656
rect 24627 7625 24639 7628
rect 24581 7619 24639 7625
rect 24670 7616 24676 7628
rect 24728 7616 24734 7668
rect 1104 7362 26864 7384
rect 1104 7310 5648 7362
rect 5700 7310 5712 7362
rect 5764 7310 5776 7362
rect 5828 7310 5840 7362
rect 5892 7310 14982 7362
rect 15034 7310 15046 7362
rect 15098 7310 15110 7362
rect 15162 7310 15174 7362
rect 15226 7310 24315 7362
rect 24367 7310 24379 7362
rect 24431 7310 24443 7362
rect 24495 7310 24507 7362
rect 24559 7310 26864 7362
rect 1104 7288 26864 7310
rect 21174 7248 21180 7260
rect 21135 7220 21180 7248
rect 21174 7208 21180 7220
rect 21232 7208 21238 7260
rect 24670 7248 24676 7260
rect 24631 7220 24676 7248
rect 24670 7208 24676 7220
rect 24728 7208 24734 7260
rect 20993 7047 21051 7053
rect 20993 7013 21005 7047
rect 21039 7044 21051 7047
rect 21039 7016 21680 7044
rect 21039 7013 21051 7016
rect 20993 7007 21051 7013
rect 21652 6920 21680 7016
rect 21634 6908 21640 6920
rect 21595 6880 21640 6908
rect 21634 6868 21640 6880
rect 21692 6868 21698 6920
rect 1104 6818 26864 6840
rect 1104 6766 10315 6818
rect 10367 6766 10379 6818
rect 10431 6766 10443 6818
rect 10495 6766 10507 6818
rect 10559 6766 19648 6818
rect 19700 6766 19712 6818
rect 19764 6766 19776 6818
rect 19828 6766 19840 6818
rect 19892 6766 26864 6818
rect 1104 6744 26864 6766
rect 20346 6568 20352 6580
rect 20307 6540 20352 6568
rect 20346 6528 20352 6540
rect 20404 6528 20410 6580
rect 20533 6435 20591 6441
rect 20533 6401 20545 6435
rect 20579 6432 20591 6435
rect 21266 6432 21272 6444
rect 20579 6404 21272 6432
rect 20579 6401 20591 6404
rect 20533 6395 20591 6401
rect 21266 6392 21272 6404
rect 21324 6392 21330 6444
rect 1104 6274 26864 6296
rect 1104 6222 5648 6274
rect 5700 6222 5712 6274
rect 5764 6222 5776 6274
rect 5828 6222 5840 6274
rect 5892 6222 14982 6274
rect 15034 6222 15046 6274
rect 15098 6222 15110 6274
rect 15162 6222 15174 6274
rect 15226 6222 24315 6274
rect 24367 6222 24379 6274
rect 24431 6222 24443 6274
rect 24495 6222 24507 6274
rect 24559 6222 26864 6274
rect 1104 6200 26864 6222
rect 19797 6163 19855 6169
rect 19797 6129 19809 6163
rect 19843 6160 19855 6163
rect 19978 6160 19984 6172
rect 19843 6132 19984 6160
rect 19843 6129 19855 6132
rect 19797 6123 19855 6129
rect 19978 6120 19984 6132
rect 20036 6120 20042 6172
rect 20346 6160 20352 6172
rect 20307 6132 20352 6160
rect 20346 6120 20352 6132
rect 20404 6120 20410 6172
rect 19613 5959 19671 5965
rect 19613 5925 19625 5959
rect 19659 5925 19671 5959
rect 19613 5919 19671 5925
rect 19521 5823 19579 5829
rect 19521 5789 19533 5823
rect 19567 5820 19579 5823
rect 19628 5820 19656 5919
rect 20070 5820 20076 5832
rect 19567 5792 20076 5820
rect 19567 5789 19579 5792
rect 19521 5783 19579 5789
rect 20070 5780 20076 5792
rect 20128 5780 20134 5832
rect 1104 5730 26864 5752
rect 1104 5678 10315 5730
rect 10367 5678 10379 5730
rect 10431 5678 10443 5730
rect 10495 5678 10507 5730
rect 10559 5678 19648 5730
rect 19700 5678 19712 5730
rect 19764 5678 19776 5730
rect 19828 5678 19840 5730
rect 19892 5678 26864 5730
rect 1104 5656 26864 5678
rect 1104 5186 26864 5208
rect 1104 5134 5648 5186
rect 5700 5134 5712 5186
rect 5764 5134 5776 5186
rect 5828 5134 5840 5186
rect 5892 5134 14982 5186
rect 15034 5134 15046 5186
rect 15098 5134 15110 5186
rect 15162 5134 15174 5186
rect 15226 5134 24315 5186
rect 24367 5134 24379 5186
rect 24431 5134 24443 5186
rect 24495 5134 24507 5186
rect 24559 5134 26864 5186
rect 1104 5112 26864 5134
rect 23474 5032 23480 5084
rect 23532 5072 23538 5084
rect 24765 5075 24823 5081
rect 24765 5072 24777 5075
rect 23532 5044 24777 5072
rect 23532 5032 23538 5044
rect 24765 5041 24777 5044
rect 24811 5041 24823 5075
rect 25222 5072 25228 5084
rect 25183 5044 25228 5072
rect 24765 5035 24823 5041
rect 25222 5032 25228 5044
rect 25280 5032 25286 5084
rect 24581 4871 24639 4877
rect 24581 4837 24593 4871
rect 24627 4868 24639 4871
rect 25222 4868 25228 4880
rect 24627 4840 25228 4868
rect 24627 4837 24639 4840
rect 24581 4831 24639 4837
rect 25222 4828 25228 4840
rect 25280 4828 25286 4880
rect 1104 4642 26864 4664
rect 1104 4590 10315 4642
rect 10367 4590 10379 4642
rect 10431 4590 10443 4642
rect 10495 4590 10507 4642
rect 10559 4590 19648 4642
rect 19700 4590 19712 4642
rect 19764 4590 19776 4642
rect 19828 4590 19840 4642
rect 19892 4590 26864 4642
rect 1104 4568 26864 4590
rect 24762 4528 24768 4540
rect 24723 4500 24768 4528
rect 24762 4488 24768 4500
rect 24820 4488 24826 4540
rect 24578 4392 24584 4404
rect 24539 4364 24584 4392
rect 24578 4352 24584 4364
rect 24636 4352 24642 4404
rect 1104 4098 26864 4120
rect 1104 4046 5648 4098
rect 5700 4046 5712 4098
rect 5764 4046 5776 4098
rect 5828 4046 5840 4098
rect 5892 4046 14982 4098
rect 15034 4046 15046 4098
rect 15098 4046 15110 4098
rect 15162 4046 15174 4098
rect 15226 4046 24315 4098
rect 24367 4046 24379 4098
rect 24431 4046 24443 4098
rect 24495 4046 24507 4098
rect 24559 4046 26864 4098
rect 1104 4024 26864 4046
rect 24489 3987 24547 3993
rect 24489 3953 24501 3987
rect 24535 3984 24547 3987
rect 24670 3984 24676 3996
rect 24535 3956 24676 3984
rect 24535 3953 24547 3956
rect 24489 3947 24547 3953
rect 24670 3944 24676 3956
rect 24728 3944 24734 3996
rect 25222 3848 25228 3860
rect 24596 3820 25228 3848
rect 24596 3789 24624 3820
rect 25222 3808 25228 3820
rect 25280 3808 25286 3860
rect 24581 3783 24639 3789
rect 24581 3749 24593 3783
rect 24627 3749 24639 3783
rect 24581 3743 24639 3749
rect 24762 3644 24768 3656
rect 24723 3616 24768 3644
rect 24762 3604 24768 3616
rect 24820 3604 24826 3656
rect 1104 3554 26864 3576
rect 1104 3502 10315 3554
rect 10367 3502 10379 3554
rect 10431 3502 10443 3554
rect 10495 3502 10507 3554
rect 10559 3502 19648 3554
rect 19700 3502 19712 3554
rect 19764 3502 19776 3554
rect 19828 3502 19840 3554
rect 19892 3502 26864 3554
rect 1104 3480 26864 3502
rect 1104 3010 26864 3032
rect 1104 2958 5648 3010
rect 5700 2958 5712 3010
rect 5764 2958 5776 3010
rect 5828 2958 5840 3010
rect 5892 2958 14982 3010
rect 15034 2958 15046 3010
rect 15098 2958 15110 3010
rect 15162 2958 15174 3010
rect 15226 2958 24315 3010
rect 24367 2958 24379 3010
rect 24431 2958 24443 3010
rect 24495 2958 24507 3010
rect 24559 2958 26864 3010
rect 1104 2936 26864 2958
rect 16301 2899 16359 2905
rect 16301 2865 16313 2899
rect 16347 2896 16359 2899
rect 16482 2896 16488 2908
rect 16347 2868 16488 2896
rect 16347 2865 16359 2868
rect 16301 2859 16359 2865
rect 16482 2856 16488 2868
rect 16540 2856 16546 2908
rect 24762 2896 24768 2908
rect 24723 2868 24768 2896
rect 24762 2856 24768 2868
rect 24820 2856 24826 2908
rect 16758 2760 16764 2772
rect 16132 2732 16764 2760
rect 16132 2701 16160 2732
rect 16758 2720 16764 2732
rect 16816 2720 16822 2772
rect 16117 2695 16175 2701
rect 16117 2661 16129 2695
rect 16163 2661 16175 2695
rect 16117 2655 16175 2661
rect 24581 2695 24639 2701
rect 24581 2661 24593 2695
rect 24627 2692 24639 2695
rect 24670 2692 24676 2704
rect 24627 2664 24676 2692
rect 24627 2661 24639 2664
rect 24581 2655 24639 2661
rect 24670 2652 24676 2664
rect 24728 2692 24734 2704
rect 25133 2695 25191 2701
rect 25133 2692 25145 2695
rect 24728 2664 25145 2692
rect 24728 2652 24734 2664
rect 25133 2661 25145 2664
rect 25179 2661 25191 2695
rect 25133 2655 25191 2661
rect 1104 2466 26864 2488
rect 1104 2414 10315 2466
rect 10367 2414 10379 2466
rect 10431 2414 10443 2466
rect 10495 2414 10507 2466
rect 10559 2414 19648 2466
rect 19700 2414 19712 2466
rect 19764 2414 19776 2466
rect 19828 2414 19840 2466
rect 19892 2414 26864 2466
rect 1104 2392 26864 2414
rect 24581 2219 24639 2225
rect 24581 2185 24593 2219
rect 24627 2216 24639 2219
rect 25222 2216 25228 2228
rect 24627 2188 25228 2216
rect 24627 2185 24639 2188
rect 24581 2179 24639 2185
rect 25222 2176 25228 2188
rect 25280 2176 25286 2228
rect 24762 2080 24768 2092
rect 24723 2052 24768 2080
rect 24762 2040 24768 2052
rect 24820 2040 24826 2092
rect 25222 2012 25228 2024
rect 25183 1984 25228 2012
rect 25222 1972 25228 1984
rect 25280 1972 25286 2024
rect 1104 1922 26864 1944
rect 1104 1870 5648 1922
rect 5700 1870 5712 1922
rect 5764 1870 5776 1922
rect 5828 1870 5840 1922
rect 5892 1870 14982 1922
rect 15034 1870 15046 1922
rect 15098 1870 15110 1922
rect 15162 1870 15174 1922
rect 15226 1870 24315 1922
rect 24367 1870 24379 1922
rect 24431 1870 24443 1922
rect 24495 1870 24507 1922
rect 24559 1870 26864 1922
rect 1104 1848 26864 1870
<< via1 >>
rect 19984 26248 20036 26300
rect 24768 26248 24820 26300
rect 10315 25262 10367 25314
rect 10379 25262 10431 25314
rect 10443 25262 10495 25314
rect 10507 25262 10559 25314
rect 19648 25262 19700 25314
rect 19712 25262 19764 25314
rect 19776 25262 19828 25314
rect 19840 25262 19892 25314
rect 23940 24820 23992 24872
rect 5648 24718 5700 24770
rect 5712 24718 5764 24770
rect 5776 24718 5828 24770
rect 5840 24718 5892 24770
rect 14982 24718 15034 24770
rect 15046 24718 15098 24770
rect 15110 24718 15162 24770
rect 15174 24718 15226 24770
rect 24315 24718 24367 24770
rect 24379 24718 24431 24770
rect 24443 24718 24495 24770
rect 24507 24718 24559 24770
rect 21732 24548 21784 24600
rect 24768 24548 24820 24600
rect 15292 24480 15344 24532
rect 16488 24480 16540 24532
rect 17960 24480 18012 24532
rect 18880 24480 18932 24532
rect 23940 24523 23992 24532
rect 23940 24489 23949 24523
rect 23949 24489 23983 24523
rect 23983 24489 23992 24523
rect 23940 24480 23992 24489
rect 20720 24412 20772 24464
rect 21272 24412 21324 24464
rect 23756 24455 23808 24464
rect 23756 24421 23765 24455
rect 23765 24421 23799 24455
rect 23799 24421 23808 24455
rect 23756 24412 23808 24421
rect 24952 24455 25004 24464
rect 24952 24421 24961 24455
rect 24961 24421 24995 24455
rect 24995 24421 25004 24455
rect 24952 24412 25004 24421
rect 23204 24387 23256 24396
rect 23204 24353 23213 24387
rect 23213 24353 23247 24387
rect 23247 24353 23256 24387
rect 23204 24344 23256 24353
rect 23572 24276 23624 24328
rect 25136 24319 25188 24328
rect 25136 24285 25145 24319
rect 25145 24285 25179 24319
rect 25179 24285 25188 24319
rect 25136 24276 25188 24285
rect 10315 24174 10367 24226
rect 10379 24174 10431 24226
rect 10443 24174 10495 24226
rect 10507 24174 10559 24226
rect 19648 24174 19700 24226
rect 19712 24174 19764 24226
rect 19776 24174 19828 24226
rect 19840 24174 19892 24226
rect 17316 24072 17368 24124
rect 23756 24072 23808 24124
rect 23848 24072 23900 24124
rect 24216 24072 24268 24124
rect 19340 24004 19392 24056
rect 20444 24004 20496 24056
rect 11152 23936 11204 23988
rect 12900 23936 12952 23988
rect 15108 23936 15160 23988
rect 17224 23936 17276 23988
rect 19892 23979 19944 23988
rect 19892 23945 19926 23979
rect 19926 23945 19944 23979
rect 19892 23936 19944 23945
rect 23296 23936 23348 23988
rect 13728 23911 13780 23920
rect 13728 23877 13737 23911
rect 13737 23877 13771 23911
rect 13771 23877 13780 23911
rect 13728 23868 13780 23877
rect 19616 23911 19668 23920
rect 19616 23877 19625 23911
rect 19625 23877 19659 23911
rect 19659 23877 19668 23911
rect 19616 23868 19668 23877
rect 23572 23868 23624 23920
rect 24676 23911 24728 23920
rect 24676 23877 24685 23911
rect 24685 23877 24719 23911
rect 24719 23877 24728 23911
rect 24676 23868 24728 23877
rect 23756 23800 23808 23852
rect 12348 23732 12400 23784
rect 14464 23732 14516 23784
rect 16764 23732 16816 23784
rect 17224 23775 17276 23784
rect 17224 23741 17233 23775
rect 17233 23741 17267 23775
rect 17267 23741 17276 23775
rect 17224 23732 17276 23741
rect 19892 23732 19944 23784
rect 24032 23732 24084 23784
rect 5648 23630 5700 23682
rect 5712 23630 5764 23682
rect 5776 23630 5828 23682
rect 5840 23630 5892 23682
rect 14982 23630 15034 23682
rect 15046 23630 15098 23682
rect 15110 23630 15162 23682
rect 15174 23630 15226 23682
rect 24315 23630 24367 23682
rect 24379 23630 24431 23682
rect 24443 23630 24495 23682
rect 24507 23630 24559 23682
rect 11152 23528 11204 23580
rect 12900 23571 12952 23580
rect 12900 23537 12909 23571
rect 12909 23537 12943 23571
rect 12943 23537 12952 23571
rect 12900 23528 12952 23537
rect 13728 23528 13780 23580
rect 14556 23528 14608 23580
rect 15936 23528 15988 23580
rect 16304 23571 16356 23580
rect 16304 23537 16313 23571
rect 16313 23537 16347 23571
rect 16347 23537 16356 23571
rect 17868 23571 17920 23580
rect 16304 23528 16356 23537
rect 17868 23537 17877 23571
rect 17877 23537 17911 23571
rect 17911 23537 17920 23571
rect 17868 23528 17920 23537
rect 19800 23528 19852 23580
rect 22744 23528 22796 23580
rect 23296 23571 23348 23580
rect 23296 23537 23305 23571
rect 23305 23537 23339 23571
rect 23339 23537 23348 23571
rect 23296 23528 23348 23537
rect 23664 23528 23716 23580
rect 23940 23528 23992 23580
rect 24676 23528 24728 23580
rect 19616 23460 19668 23512
rect 20168 23460 20220 23512
rect 19892 23435 19944 23444
rect 19892 23401 19901 23435
rect 19901 23401 19935 23435
rect 19935 23401 19944 23435
rect 19892 23392 19944 23401
rect 9772 23324 9824 23376
rect 10784 23367 10836 23376
rect 10784 23333 10793 23367
rect 10793 23333 10827 23367
rect 10827 23333 10836 23367
rect 10784 23324 10836 23333
rect 11888 23367 11940 23376
rect 11888 23333 11897 23367
rect 11897 23333 11931 23367
rect 11931 23333 11940 23367
rect 11888 23324 11940 23333
rect 12532 23324 12584 23376
rect 14096 23367 14148 23376
rect 14096 23333 14105 23367
rect 14105 23333 14139 23367
rect 14139 23333 14148 23367
rect 14096 23324 14148 23333
rect 15292 23367 15344 23376
rect 15292 23333 15301 23367
rect 15301 23333 15335 23367
rect 15335 23333 15344 23367
rect 15292 23324 15344 23333
rect 16764 23367 16816 23376
rect 16764 23333 16798 23367
rect 16798 23333 16816 23367
rect 16764 23324 16816 23333
rect 19432 23324 19484 23376
rect 19984 23324 20036 23376
rect 20352 23324 20404 23376
rect 19064 23299 19116 23308
rect 19064 23265 19073 23299
rect 19073 23265 19107 23299
rect 19107 23265 19116 23299
rect 19064 23256 19116 23265
rect 24032 23299 24084 23308
rect 24032 23265 24066 23299
rect 24066 23265 24084 23299
rect 24032 23256 24084 23265
rect 25044 23256 25096 23308
rect 9864 23231 9916 23240
rect 9864 23197 9873 23231
rect 9873 23197 9907 23231
rect 9907 23197 9916 23231
rect 9864 23188 9916 23197
rect 10968 23231 11020 23240
rect 10968 23197 10977 23231
rect 10977 23197 11011 23231
rect 11011 23197 11020 23231
rect 10968 23188 11020 23197
rect 12072 23231 12124 23240
rect 12072 23197 12081 23231
rect 12081 23197 12115 23231
rect 12115 23197 12124 23231
rect 12072 23188 12124 23197
rect 14280 23188 14332 23240
rect 19340 23188 19392 23240
rect 21548 23188 21600 23240
rect 23664 23231 23716 23240
rect 23664 23197 23673 23231
rect 23673 23197 23707 23231
rect 23707 23197 23716 23231
rect 23664 23188 23716 23197
rect 10315 23086 10367 23138
rect 10379 23086 10431 23138
rect 10443 23086 10495 23138
rect 10507 23086 10559 23138
rect 19648 23086 19700 23138
rect 19712 23086 19764 23138
rect 19776 23086 19828 23138
rect 19840 23086 19892 23138
rect 18972 22984 19024 23036
rect 19432 22984 19484 23036
rect 23572 22984 23624 23036
rect 25044 23027 25096 23036
rect 25044 22993 25053 23027
rect 25053 22993 25087 23027
rect 25087 22993 25096 23027
rect 25044 22984 25096 22993
rect 19984 22916 20036 22968
rect 14188 22891 14240 22900
rect 14188 22857 14197 22891
rect 14197 22857 14231 22891
rect 14231 22857 14240 22891
rect 14188 22848 14240 22857
rect 14280 22891 14332 22900
rect 14280 22857 14289 22891
rect 14289 22857 14323 22891
rect 14323 22857 14332 22891
rect 14280 22848 14332 22857
rect 17500 22848 17552 22900
rect 18236 22848 18288 22900
rect 19708 22848 19760 22900
rect 20168 22848 20220 22900
rect 22652 22848 22704 22900
rect 23756 22848 23808 22900
rect 24216 22848 24268 22900
rect 14096 22780 14148 22832
rect 14464 22823 14516 22832
rect 14464 22789 14473 22823
rect 14473 22789 14507 22823
rect 14507 22789 14516 22823
rect 14464 22780 14516 22789
rect 16120 22780 16172 22832
rect 16764 22712 16816 22764
rect 17960 22780 18012 22832
rect 18604 22823 18656 22832
rect 18604 22789 18613 22823
rect 18613 22789 18647 22823
rect 18647 22789 18656 22823
rect 18604 22780 18656 22789
rect 23664 22823 23716 22832
rect 23664 22789 23673 22823
rect 23673 22789 23707 22823
rect 23707 22789 23716 22823
rect 23664 22780 23716 22789
rect 17684 22712 17736 22764
rect 11336 22644 11388 22696
rect 13636 22687 13688 22696
rect 13636 22653 13645 22687
rect 13645 22653 13679 22687
rect 13679 22653 13688 22687
rect 13636 22644 13688 22653
rect 13820 22687 13872 22696
rect 13820 22653 13829 22687
rect 13829 22653 13863 22687
rect 13863 22653 13872 22687
rect 13820 22644 13872 22653
rect 16856 22644 16908 22696
rect 18052 22687 18104 22696
rect 18052 22653 18061 22687
rect 18061 22653 18095 22687
rect 18095 22653 18104 22687
rect 18052 22644 18104 22653
rect 20536 22644 20588 22696
rect 22008 22687 22060 22696
rect 22008 22653 22017 22687
rect 22017 22653 22051 22687
rect 22051 22653 22060 22687
rect 22008 22644 22060 22653
rect 22744 22687 22796 22696
rect 22744 22653 22753 22687
rect 22753 22653 22787 22687
rect 22787 22653 22796 22687
rect 22744 22644 22796 22653
rect 5648 22542 5700 22594
rect 5712 22542 5764 22594
rect 5776 22542 5828 22594
rect 5840 22542 5892 22594
rect 14982 22542 15034 22594
rect 15046 22542 15098 22594
rect 15110 22542 15162 22594
rect 15174 22542 15226 22594
rect 24315 22542 24367 22594
rect 24379 22542 24431 22594
rect 24443 22542 24495 22594
rect 24507 22542 24559 22594
rect 13544 22483 13596 22492
rect 13544 22449 13553 22483
rect 13553 22449 13587 22483
rect 13587 22449 13596 22483
rect 13544 22440 13596 22449
rect 14188 22440 14240 22492
rect 14280 22440 14332 22492
rect 17500 22440 17552 22492
rect 17684 22483 17736 22492
rect 17684 22449 17693 22483
rect 17693 22449 17727 22483
rect 17727 22449 17736 22483
rect 17684 22440 17736 22449
rect 18604 22483 18656 22492
rect 18604 22449 18613 22483
rect 18613 22449 18647 22483
rect 18647 22449 18656 22483
rect 18604 22440 18656 22449
rect 18972 22483 19024 22492
rect 18972 22449 18981 22483
rect 18981 22449 19015 22483
rect 19015 22449 19024 22483
rect 18972 22440 19024 22449
rect 19432 22440 19484 22492
rect 19708 22483 19760 22492
rect 19708 22449 19717 22483
rect 19717 22449 19751 22483
rect 19751 22449 19760 22483
rect 19708 22440 19760 22449
rect 19984 22440 20036 22492
rect 25228 22440 25280 22492
rect 16120 22415 16172 22424
rect 16120 22381 16129 22415
rect 16129 22381 16163 22415
rect 16163 22381 16172 22415
rect 16120 22372 16172 22381
rect 13820 22304 13872 22356
rect 16304 22347 16356 22356
rect 10876 22236 10928 22288
rect 13636 22236 13688 22288
rect 16304 22313 16313 22347
rect 16313 22313 16347 22347
rect 16347 22313 16356 22347
rect 16304 22304 16356 22313
rect 16856 22236 16908 22288
rect 20628 22236 20680 22288
rect 11336 22168 11388 22220
rect 12164 22143 12216 22152
rect 12164 22109 12173 22143
rect 12173 22109 12207 22143
rect 12207 22109 12216 22143
rect 12164 22100 12216 22109
rect 13728 22100 13780 22152
rect 14188 22168 14240 22220
rect 22008 22236 22060 22288
rect 23664 22236 23716 22288
rect 24584 22279 24636 22288
rect 24584 22245 24593 22279
rect 24593 22245 24627 22279
rect 24627 22245 24636 22279
rect 24584 22236 24636 22245
rect 14096 22100 14148 22152
rect 18236 22143 18288 22152
rect 18236 22109 18245 22143
rect 18245 22109 18279 22143
rect 18279 22109 18288 22143
rect 18236 22100 18288 22109
rect 20168 22100 20220 22152
rect 24216 22143 24268 22152
rect 24216 22109 24225 22143
rect 24225 22109 24259 22143
rect 24259 22109 24268 22143
rect 24216 22100 24268 22109
rect 24676 22100 24728 22152
rect 10315 21998 10367 22050
rect 10379 21998 10431 22050
rect 10443 21998 10495 22050
rect 10507 21998 10559 22050
rect 19648 21998 19700 22050
rect 19712 21998 19764 22050
rect 19776 21998 19828 22050
rect 19840 21998 19892 22050
rect 13636 21896 13688 21948
rect 16304 21939 16356 21948
rect 16304 21905 16313 21939
rect 16313 21905 16347 21939
rect 16347 21905 16356 21939
rect 16304 21896 16356 21905
rect 18236 21896 18288 21948
rect 20168 21939 20220 21948
rect 20168 21905 20177 21939
rect 20177 21905 20211 21939
rect 20211 21905 20220 21939
rect 20168 21896 20220 21905
rect 21732 21939 21784 21948
rect 21732 21905 21741 21939
rect 21741 21905 21775 21939
rect 21775 21905 21784 21939
rect 21732 21896 21784 21905
rect 22652 21939 22704 21948
rect 22652 21905 22661 21939
rect 22661 21905 22695 21939
rect 22695 21905 22704 21939
rect 22652 21896 22704 21905
rect 11152 21871 11204 21880
rect 11152 21837 11161 21871
rect 11161 21837 11195 21871
rect 11195 21837 11204 21871
rect 11152 21828 11204 21837
rect 14096 21828 14148 21880
rect 17684 21828 17736 21880
rect 18052 21803 18104 21812
rect 18052 21769 18061 21803
rect 18061 21769 18095 21803
rect 18095 21769 18104 21803
rect 18052 21760 18104 21769
rect 10508 21692 10560 21744
rect 11336 21735 11388 21744
rect 11336 21701 11345 21735
rect 11345 21701 11379 21735
rect 11379 21701 11388 21735
rect 13636 21735 13688 21744
rect 11336 21692 11388 21701
rect 13636 21701 13645 21735
rect 13645 21701 13679 21735
rect 13679 21701 13688 21735
rect 13636 21692 13688 21701
rect 19340 21692 19392 21744
rect 19524 21692 19576 21744
rect 25228 21803 25280 21812
rect 20536 21692 20588 21744
rect 21364 21692 21416 21744
rect 22008 21735 22060 21744
rect 22008 21701 22017 21735
rect 22017 21701 22051 21735
rect 22051 21701 22060 21735
rect 22008 21692 22060 21701
rect 23480 21692 23532 21744
rect 24216 21735 24268 21744
rect 24216 21701 24225 21735
rect 24225 21701 24259 21735
rect 24259 21701 24268 21735
rect 24216 21692 24268 21701
rect 18236 21667 18288 21676
rect 18236 21633 18245 21667
rect 18245 21633 18279 21667
rect 18279 21633 18288 21667
rect 18236 21624 18288 21633
rect 20628 21624 20680 21676
rect 24032 21624 24084 21676
rect 25228 21769 25237 21803
rect 25237 21769 25271 21803
rect 25271 21769 25280 21803
rect 25228 21760 25280 21769
rect 10600 21599 10652 21608
rect 10600 21565 10609 21599
rect 10609 21565 10643 21599
rect 10643 21565 10652 21599
rect 10600 21556 10652 21565
rect 10692 21556 10744 21608
rect 23480 21556 23532 21608
rect 23664 21599 23716 21608
rect 23664 21565 23673 21599
rect 23673 21565 23707 21599
rect 23707 21565 23716 21599
rect 23664 21556 23716 21565
rect 24860 21556 24912 21608
rect 5648 21454 5700 21506
rect 5712 21454 5764 21506
rect 5776 21454 5828 21506
rect 5840 21454 5892 21506
rect 14982 21454 15034 21506
rect 15046 21454 15098 21506
rect 15110 21454 15162 21506
rect 15174 21454 15226 21506
rect 24315 21454 24367 21506
rect 24379 21454 24431 21506
rect 24443 21454 24495 21506
rect 24507 21454 24559 21506
rect 9128 21352 9180 21404
rect 10508 21395 10560 21404
rect 10508 21361 10517 21395
rect 10517 21361 10551 21395
rect 10551 21361 10560 21395
rect 10508 21352 10560 21361
rect 11336 21352 11388 21404
rect 13636 21395 13688 21404
rect 13636 21361 13645 21395
rect 13645 21361 13679 21395
rect 13679 21361 13688 21395
rect 13636 21352 13688 21361
rect 13820 21352 13872 21404
rect 14096 21395 14148 21404
rect 14096 21361 14105 21395
rect 14105 21361 14139 21395
rect 14139 21361 14148 21395
rect 14096 21352 14148 21361
rect 18052 21352 18104 21404
rect 18144 21395 18196 21404
rect 18144 21361 18153 21395
rect 18153 21361 18187 21395
rect 18187 21361 18196 21395
rect 18144 21352 18196 21361
rect 20168 21352 20220 21404
rect 20720 21395 20772 21404
rect 20720 21361 20729 21395
rect 20729 21361 20763 21395
rect 20763 21361 20772 21395
rect 20720 21352 20772 21361
rect 22008 21352 22060 21404
rect 23480 21352 23532 21404
rect 24032 21352 24084 21404
rect 24216 21395 24268 21404
rect 24216 21361 24225 21395
rect 24225 21361 24259 21395
rect 24259 21361 24268 21395
rect 24216 21352 24268 21361
rect 25228 21395 25280 21404
rect 25228 21361 25237 21395
rect 25237 21361 25271 21395
rect 25271 21361 25280 21395
rect 25228 21352 25280 21361
rect 24216 21216 24268 21268
rect 24676 21216 24728 21268
rect 10784 21148 10836 21200
rect 23664 21148 23716 21200
rect 10600 21080 10652 21132
rect 9680 21055 9732 21064
rect 9680 21021 9689 21055
rect 9689 21021 9723 21055
rect 9723 21021 9732 21055
rect 9680 21012 9732 21021
rect 14556 21012 14608 21064
rect 17776 21055 17828 21064
rect 17776 21021 17785 21055
rect 17785 21021 17819 21055
rect 17819 21021 17828 21055
rect 17776 21012 17828 21021
rect 20168 21012 20220 21064
rect 24676 21012 24728 21064
rect 10315 20910 10367 20962
rect 10379 20910 10431 20962
rect 10443 20910 10495 20962
rect 10507 20910 10559 20962
rect 19648 20910 19700 20962
rect 19712 20910 19764 20962
rect 19776 20910 19828 20962
rect 19840 20910 19892 20962
rect 11336 20808 11388 20860
rect 14188 20851 14240 20860
rect 14188 20817 14197 20851
rect 14197 20817 14231 20851
rect 14231 20817 14240 20851
rect 14188 20808 14240 20817
rect 18512 20851 18564 20860
rect 18512 20817 18521 20851
rect 18521 20817 18555 20851
rect 18555 20817 18564 20851
rect 18512 20808 18564 20817
rect 19524 20851 19576 20860
rect 19524 20817 19533 20851
rect 19533 20817 19567 20851
rect 19567 20817 19576 20851
rect 19524 20808 19576 20817
rect 21364 20851 21416 20860
rect 21364 20817 21373 20851
rect 21373 20817 21407 20851
rect 21407 20817 21416 20851
rect 21364 20808 21416 20817
rect 21732 20851 21784 20860
rect 21732 20817 21741 20851
rect 21741 20817 21775 20851
rect 21775 20817 21784 20851
rect 21732 20808 21784 20817
rect 22008 20808 22060 20860
rect 23940 20808 23992 20860
rect 25136 20808 25188 20860
rect 11060 20740 11112 20792
rect 9680 20672 9732 20724
rect 10140 20604 10192 20656
rect 10692 20604 10744 20656
rect 12164 20740 12216 20792
rect 12440 20715 12492 20724
rect 12440 20681 12449 20715
rect 12449 20681 12483 20715
rect 12483 20681 12492 20715
rect 14556 20715 14608 20724
rect 12440 20672 12492 20681
rect 14556 20681 14565 20715
rect 14565 20681 14599 20715
rect 14599 20681 14608 20715
rect 14556 20672 14608 20681
rect 16764 20715 16816 20724
rect 16764 20681 16773 20715
rect 16773 20681 16807 20715
rect 16807 20681 16816 20715
rect 16764 20672 16816 20681
rect 18420 20715 18472 20724
rect 18420 20681 18429 20715
rect 18429 20681 18463 20715
rect 18463 20681 18472 20715
rect 18420 20672 18472 20681
rect 19984 20715 20036 20724
rect 19984 20681 19993 20715
rect 19993 20681 20027 20715
rect 20027 20681 20036 20715
rect 19984 20672 20036 20681
rect 14648 20647 14700 20656
rect 14648 20613 14657 20647
rect 14657 20613 14691 20647
rect 14691 20613 14700 20647
rect 14648 20604 14700 20613
rect 12440 20536 12492 20588
rect 12624 20579 12676 20588
rect 12624 20545 12633 20579
rect 12633 20545 12667 20579
rect 12667 20545 12676 20579
rect 12624 20536 12676 20545
rect 14096 20536 14148 20588
rect 16028 20604 16080 20656
rect 11152 20468 11204 20520
rect 16212 20511 16264 20520
rect 16212 20477 16221 20511
rect 16221 20477 16255 20511
rect 16255 20477 16264 20511
rect 16212 20468 16264 20477
rect 16672 20468 16724 20520
rect 16856 20468 16908 20520
rect 17776 20604 17828 20656
rect 20168 20647 20220 20656
rect 20168 20613 20177 20647
rect 20177 20613 20211 20647
rect 20211 20613 20220 20647
rect 20168 20604 20220 20613
rect 24032 20604 24084 20656
rect 24952 20672 25004 20724
rect 25320 20715 25372 20724
rect 25320 20681 25329 20715
rect 25329 20681 25363 20715
rect 25363 20681 25372 20715
rect 25320 20672 25372 20681
rect 24860 20647 24912 20656
rect 24860 20613 24869 20647
rect 24869 20613 24903 20647
rect 24903 20613 24912 20647
rect 24860 20604 24912 20613
rect 20260 20536 20312 20588
rect 19248 20468 19300 20520
rect 20720 20468 20772 20520
rect 23940 20468 23992 20520
rect 5648 20366 5700 20418
rect 5712 20366 5764 20418
rect 5776 20366 5828 20418
rect 5840 20366 5892 20418
rect 14982 20366 15034 20418
rect 15046 20366 15098 20418
rect 15110 20366 15162 20418
rect 15174 20366 15226 20418
rect 24315 20366 24367 20418
rect 24379 20366 24431 20418
rect 24443 20366 24495 20418
rect 24507 20366 24559 20418
rect 9680 20264 9732 20316
rect 12440 20264 12492 20316
rect 14096 20307 14148 20316
rect 14096 20273 14105 20307
rect 14105 20273 14139 20307
rect 14139 20273 14148 20307
rect 14096 20264 14148 20273
rect 14556 20264 14608 20316
rect 16028 20307 16080 20316
rect 16028 20273 16037 20307
rect 16037 20273 16071 20307
rect 16071 20273 16080 20307
rect 16028 20264 16080 20273
rect 18512 20264 18564 20316
rect 19800 20307 19852 20316
rect 10140 20239 10192 20248
rect 10140 20205 10149 20239
rect 10149 20205 10183 20239
rect 10183 20205 10192 20239
rect 10140 20196 10192 20205
rect 14648 20239 14700 20248
rect 14648 20205 14657 20239
rect 14657 20205 14691 20239
rect 14691 20205 14700 20239
rect 14648 20196 14700 20205
rect 10048 20128 10100 20180
rect 10968 20128 11020 20180
rect 18420 20128 18472 20180
rect 19800 20273 19809 20307
rect 19809 20273 19843 20307
rect 19843 20273 19852 20307
rect 19800 20264 19852 20273
rect 19984 20264 20036 20316
rect 20168 20264 20220 20316
rect 24032 20264 24084 20316
rect 25136 20307 25188 20316
rect 25136 20273 25145 20307
rect 25145 20273 25179 20307
rect 25179 20273 25188 20307
rect 25136 20264 25188 20273
rect 19248 20171 19300 20180
rect 19248 20137 19257 20171
rect 19257 20137 19291 20171
rect 19291 20137 19300 20171
rect 19248 20128 19300 20137
rect 22652 20128 22704 20180
rect 24308 20171 24360 20180
rect 10876 20060 10928 20112
rect 12256 20060 12308 20112
rect 14464 20060 14516 20112
rect 16212 20103 16264 20112
rect 16212 20069 16221 20103
rect 16221 20069 16255 20103
rect 16255 20069 16264 20103
rect 16212 20060 16264 20069
rect 19064 20103 19116 20112
rect 19064 20069 19073 20103
rect 19073 20069 19107 20103
rect 19107 20069 19116 20103
rect 19064 20060 19116 20069
rect 20720 20060 20772 20112
rect 24308 20137 24317 20171
rect 24317 20137 24351 20171
rect 24351 20137 24360 20171
rect 24308 20128 24360 20137
rect 11796 19992 11848 20044
rect 15844 19992 15896 20044
rect 23480 20035 23532 20044
rect 23480 20001 23489 20035
rect 23489 20001 23523 20035
rect 23523 20001 23532 20035
rect 23480 19992 23532 20001
rect 25320 20060 25372 20112
rect 12808 19967 12860 19976
rect 12808 19933 12817 19967
rect 12817 19933 12851 19967
rect 12851 19933 12860 19967
rect 12808 19924 12860 19933
rect 14188 19967 14240 19976
rect 14188 19933 14197 19967
rect 14197 19933 14231 19967
rect 14231 19933 14240 19967
rect 14188 19924 14240 19933
rect 17776 19924 17828 19976
rect 18696 19967 18748 19976
rect 18696 19933 18705 19967
rect 18705 19933 18739 19967
rect 18739 19933 18748 19967
rect 18696 19924 18748 19933
rect 21088 19967 21140 19976
rect 21088 19933 21097 19967
rect 21097 19933 21131 19967
rect 21131 19933 21140 19967
rect 21088 19924 21140 19933
rect 23388 19924 23440 19976
rect 23664 19967 23716 19976
rect 23664 19933 23673 19967
rect 23673 19933 23707 19967
rect 23707 19933 23716 19967
rect 23664 19924 23716 19933
rect 25504 19992 25556 20044
rect 25412 19967 25464 19976
rect 25412 19933 25421 19967
rect 25421 19933 25455 19967
rect 25455 19933 25464 19967
rect 25412 19924 25464 19933
rect 25780 19967 25832 19976
rect 25780 19933 25789 19967
rect 25789 19933 25823 19967
rect 25823 19933 25832 19967
rect 25780 19924 25832 19933
rect 10315 19822 10367 19874
rect 10379 19822 10431 19874
rect 10443 19822 10495 19874
rect 10507 19822 10559 19874
rect 19648 19822 19700 19874
rect 19712 19822 19764 19874
rect 19776 19822 19828 19874
rect 19840 19822 19892 19874
rect 11244 19763 11296 19772
rect 11244 19729 11253 19763
rect 11253 19729 11287 19763
rect 11287 19729 11296 19763
rect 11244 19720 11296 19729
rect 13636 19763 13688 19772
rect 13636 19729 13645 19763
rect 13645 19729 13679 19763
rect 13679 19729 13688 19763
rect 13636 19720 13688 19729
rect 13728 19720 13780 19772
rect 15844 19763 15896 19772
rect 15844 19729 15853 19763
rect 15853 19729 15887 19763
rect 15887 19729 15896 19763
rect 15844 19720 15896 19729
rect 16396 19763 16448 19772
rect 16396 19729 16405 19763
rect 16405 19729 16439 19763
rect 16439 19729 16448 19763
rect 16396 19720 16448 19729
rect 16856 19763 16908 19772
rect 16856 19729 16865 19763
rect 16865 19729 16899 19763
rect 16899 19729 16908 19763
rect 16856 19720 16908 19729
rect 17776 19763 17828 19772
rect 17776 19729 17785 19763
rect 17785 19729 17819 19763
rect 17819 19729 17828 19763
rect 17776 19720 17828 19729
rect 18696 19720 18748 19772
rect 19984 19720 20036 19772
rect 20260 19720 20312 19772
rect 11152 19695 11204 19704
rect 11152 19661 11161 19695
rect 11161 19661 11195 19695
rect 11195 19661 11204 19695
rect 11152 19652 11204 19661
rect 19064 19695 19116 19704
rect 19064 19661 19073 19695
rect 19073 19661 19107 19695
rect 19107 19661 19116 19695
rect 19064 19652 19116 19661
rect 14096 19584 14148 19636
rect 12348 19516 12400 19568
rect 13820 19516 13872 19568
rect 14464 19559 14516 19568
rect 14464 19525 14473 19559
rect 14473 19525 14507 19559
rect 14507 19525 14516 19559
rect 14464 19516 14516 19525
rect 17960 19516 18012 19568
rect 20904 19516 20956 19568
rect 21364 19627 21416 19636
rect 21364 19593 21398 19627
rect 21398 19593 21416 19627
rect 24032 19627 24084 19636
rect 21364 19584 21416 19593
rect 24032 19593 24041 19627
rect 24041 19593 24075 19627
rect 24075 19593 24084 19627
rect 24032 19584 24084 19593
rect 24308 19627 24360 19636
rect 23572 19516 23624 19568
rect 24308 19593 24342 19627
rect 24342 19593 24360 19627
rect 24308 19584 24360 19593
rect 24860 19584 24912 19636
rect 25780 19584 25832 19636
rect 11060 19380 11112 19432
rect 11796 19423 11848 19432
rect 11796 19389 11805 19423
rect 11805 19389 11839 19423
rect 11839 19389 11848 19423
rect 11796 19380 11848 19389
rect 17316 19380 17368 19432
rect 18052 19423 18104 19432
rect 18052 19389 18061 19423
rect 18061 19389 18095 19423
rect 18095 19389 18104 19423
rect 18052 19380 18104 19389
rect 20996 19423 21048 19432
rect 20996 19389 21005 19423
rect 21005 19389 21039 19423
rect 21039 19389 21048 19423
rect 20996 19380 21048 19389
rect 22560 19380 22612 19432
rect 25504 19380 25556 19432
rect 5648 19278 5700 19330
rect 5712 19278 5764 19330
rect 5776 19278 5828 19330
rect 5840 19278 5892 19330
rect 14982 19278 15034 19330
rect 15046 19278 15098 19330
rect 15110 19278 15162 19330
rect 15174 19278 15226 19330
rect 24315 19278 24367 19330
rect 24379 19278 24431 19330
rect 24443 19278 24495 19330
rect 24507 19278 24559 19330
rect 14464 19176 14516 19228
rect 22100 19176 22152 19228
rect 23296 19176 23348 19228
rect 23572 19176 23624 19228
rect 24032 19176 24084 19228
rect 24492 19108 24544 19160
rect 25872 19108 25924 19160
rect 11244 19040 11296 19092
rect 15936 19083 15988 19092
rect 15936 19049 15945 19083
rect 15945 19049 15979 19083
rect 15979 19049 15988 19083
rect 15936 19040 15988 19049
rect 17316 19040 17368 19092
rect 11060 18972 11112 19024
rect 12256 18972 12308 19024
rect 10968 18904 11020 18956
rect 11244 18904 11296 18956
rect 12348 18904 12400 18956
rect 12808 18972 12860 19024
rect 16672 19015 16724 19024
rect 16672 18981 16681 19015
rect 16681 18981 16715 19015
rect 16715 18981 16724 19015
rect 16672 18972 16724 18981
rect 17868 18972 17920 19024
rect 19524 18972 19576 19024
rect 23664 19040 23716 19092
rect 20904 19015 20956 19024
rect 20904 18981 20913 19015
rect 20913 18981 20947 19015
rect 20947 18981 20956 19015
rect 20904 18972 20956 18981
rect 20996 18972 21048 19024
rect 23940 19015 23992 19024
rect 23940 18981 23949 19015
rect 23949 18981 23983 19015
rect 23983 18981 23992 19015
rect 23940 18972 23992 18981
rect 24308 19040 24360 19092
rect 25136 19015 25188 19024
rect 25136 18981 25145 19015
rect 25145 18981 25179 19015
rect 25179 18981 25188 19015
rect 25136 18972 25188 18981
rect 13820 18904 13872 18956
rect 15016 18947 15068 18956
rect 15016 18913 15025 18947
rect 15025 18913 15059 18947
rect 15059 18913 15068 18947
rect 15016 18904 15068 18913
rect 17500 18947 17552 18956
rect 17500 18913 17509 18947
rect 17509 18913 17543 18947
rect 17543 18913 17552 18947
rect 17500 18904 17552 18913
rect 11060 18836 11112 18888
rect 14096 18879 14148 18888
rect 14096 18845 14105 18879
rect 14105 18845 14139 18879
rect 14139 18845 14148 18879
rect 14096 18836 14148 18845
rect 15384 18836 15436 18888
rect 16396 18879 16448 18888
rect 16396 18845 16405 18879
rect 16405 18845 16439 18879
rect 16439 18845 16448 18879
rect 16396 18836 16448 18845
rect 17316 18836 17368 18888
rect 17592 18879 17644 18888
rect 17592 18845 17601 18879
rect 17601 18845 17635 18879
rect 17635 18845 17644 18879
rect 17592 18836 17644 18845
rect 17684 18836 17736 18888
rect 18144 18836 18196 18888
rect 18972 18836 19024 18888
rect 19800 18904 19852 18956
rect 21364 18904 21416 18956
rect 24308 18904 24360 18956
rect 19248 18879 19300 18888
rect 19248 18845 19257 18879
rect 19257 18845 19291 18879
rect 19291 18845 19300 18879
rect 19248 18836 19300 18845
rect 19340 18836 19392 18888
rect 20168 18836 20220 18888
rect 22284 18879 22336 18888
rect 22284 18845 22293 18879
rect 22293 18845 22327 18879
rect 22327 18845 22336 18879
rect 22284 18836 22336 18845
rect 23572 18879 23624 18888
rect 23572 18845 23581 18879
rect 23581 18845 23615 18879
rect 23615 18845 23624 18879
rect 23572 18836 23624 18845
rect 25320 18879 25372 18888
rect 25320 18845 25329 18879
rect 25329 18845 25363 18879
rect 25363 18845 25372 18879
rect 25320 18836 25372 18845
rect 10315 18734 10367 18786
rect 10379 18734 10431 18786
rect 10443 18734 10495 18786
rect 10507 18734 10559 18786
rect 19648 18734 19700 18786
rect 19712 18734 19764 18786
rect 19776 18734 19828 18786
rect 19840 18734 19892 18786
rect 11244 18675 11296 18684
rect 11244 18641 11253 18675
rect 11253 18641 11287 18675
rect 11287 18641 11296 18675
rect 11244 18632 11296 18641
rect 12808 18675 12860 18684
rect 12808 18641 12817 18675
rect 12817 18641 12851 18675
rect 12851 18641 12860 18675
rect 12808 18632 12860 18641
rect 14188 18632 14240 18684
rect 14832 18632 14884 18684
rect 15936 18675 15988 18684
rect 15936 18641 15945 18675
rect 15945 18641 15979 18675
rect 15979 18641 15988 18675
rect 15936 18632 15988 18641
rect 17684 18675 17736 18684
rect 17684 18641 17693 18675
rect 17693 18641 17727 18675
rect 17727 18641 17736 18675
rect 17684 18632 17736 18641
rect 18052 18632 18104 18684
rect 19064 18632 19116 18684
rect 19340 18675 19392 18684
rect 19340 18641 19349 18675
rect 19349 18641 19383 18675
rect 19383 18641 19392 18675
rect 19340 18632 19392 18641
rect 21364 18632 21416 18684
rect 23572 18632 23624 18684
rect 23664 18632 23716 18684
rect 24492 18632 24544 18684
rect 14096 18564 14148 18616
rect 17592 18564 17644 18616
rect 18604 18564 18656 18616
rect 21732 18564 21784 18616
rect 23940 18564 23992 18616
rect 15384 18471 15436 18480
rect 15384 18437 15393 18471
rect 15393 18437 15427 18471
rect 15427 18437 15436 18471
rect 15384 18428 15436 18437
rect 15844 18428 15896 18480
rect 18236 18428 18288 18480
rect 20536 18428 20588 18480
rect 19524 18360 19576 18412
rect 20168 18360 20220 18412
rect 22284 18428 22336 18480
rect 22560 18471 22612 18480
rect 22560 18437 22569 18471
rect 22569 18437 22603 18471
rect 22603 18437 22612 18471
rect 22560 18428 22612 18437
rect 23388 18496 23440 18548
rect 24952 18496 25004 18548
rect 25044 18496 25096 18548
rect 24308 18471 24360 18480
rect 24308 18437 24317 18471
rect 24317 18437 24351 18471
rect 24351 18437 24360 18471
rect 24308 18428 24360 18437
rect 25504 18428 25556 18480
rect 10876 18335 10928 18344
rect 10876 18301 10885 18335
rect 10885 18301 10919 18335
rect 10919 18301 10928 18335
rect 10876 18292 10928 18301
rect 14188 18292 14240 18344
rect 15292 18292 15344 18344
rect 18052 18335 18104 18344
rect 18052 18301 18061 18335
rect 18061 18301 18095 18335
rect 18095 18301 18104 18335
rect 18052 18292 18104 18301
rect 20720 18292 20772 18344
rect 22008 18335 22060 18344
rect 22008 18301 22017 18335
rect 22017 18301 22051 18335
rect 22051 18301 22060 18335
rect 22008 18292 22060 18301
rect 24216 18292 24268 18344
rect 25412 18335 25464 18344
rect 25412 18301 25421 18335
rect 25421 18301 25455 18335
rect 25455 18301 25464 18335
rect 25412 18292 25464 18301
rect 5648 18190 5700 18242
rect 5712 18190 5764 18242
rect 5776 18190 5828 18242
rect 5840 18190 5892 18242
rect 14982 18190 15034 18242
rect 15046 18190 15098 18242
rect 15110 18190 15162 18242
rect 15174 18190 15226 18242
rect 24315 18190 24367 18242
rect 24379 18190 24431 18242
rect 24443 18190 24495 18242
rect 24507 18190 24559 18242
rect 12256 18088 12308 18140
rect 12440 18131 12492 18140
rect 12440 18097 12449 18131
rect 12449 18097 12483 18131
rect 12483 18097 12492 18131
rect 12440 18088 12492 18097
rect 14832 18088 14884 18140
rect 15384 18088 15436 18140
rect 19064 18131 19116 18140
rect 19064 18097 19073 18131
rect 19073 18097 19107 18131
rect 19107 18097 19116 18131
rect 19064 18088 19116 18097
rect 20168 18131 20220 18140
rect 20168 18097 20177 18131
rect 20177 18097 20211 18131
rect 20211 18097 20220 18131
rect 20168 18088 20220 18097
rect 20996 18088 21048 18140
rect 24952 18131 25004 18140
rect 24952 18097 24961 18131
rect 24961 18097 24995 18131
rect 24995 18097 25004 18131
rect 24952 18088 25004 18097
rect 25044 18088 25096 18140
rect 15844 18063 15896 18072
rect 15844 18029 15853 18063
rect 15853 18029 15887 18063
rect 15887 18029 15896 18063
rect 15844 18020 15896 18029
rect 21732 18020 21784 18072
rect 23480 18020 23532 18072
rect 25504 18020 25556 18072
rect 14188 17995 14240 18004
rect 14188 17961 14197 17995
rect 14197 17961 14231 17995
rect 14231 17961 14240 17995
rect 14188 17952 14240 17961
rect 24216 17952 24268 18004
rect 13544 17884 13596 17936
rect 15292 17927 15344 17936
rect 15292 17893 15301 17927
rect 15301 17893 15335 17927
rect 15335 17893 15344 17927
rect 15292 17884 15344 17893
rect 11152 17816 11204 17868
rect 13452 17859 13504 17868
rect 13452 17825 13461 17859
rect 13461 17825 13495 17859
rect 13495 17825 13504 17859
rect 13452 17816 13504 17825
rect 22468 17884 22520 17936
rect 23204 17884 23256 17936
rect 23664 17884 23716 17936
rect 23848 17927 23900 17936
rect 23848 17893 23857 17927
rect 23857 17893 23891 17927
rect 23891 17893 23900 17927
rect 23848 17884 23900 17893
rect 25688 17884 25740 17936
rect 17316 17816 17368 17868
rect 22192 17859 22244 17868
rect 22192 17825 22201 17859
rect 22201 17825 22235 17859
rect 22235 17825 22244 17859
rect 22192 17816 22244 17825
rect 13636 17791 13688 17800
rect 13636 17757 13645 17791
rect 13645 17757 13679 17791
rect 13679 17757 13688 17791
rect 13636 17748 13688 17757
rect 15476 17791 15528 17800
rect 15476 17757 15485 17791
rect 15485 17757 15519 17791
rect 15519 17757 15528 17791
rect 15476 17748 15528 17757
rect 16948 17791 17000 17800
rect 16948 17757 16957 17791
rect 16957 17757 16991 17791
rect 16991 17757 17000 17791
rect 16948 17748 17000 17757
rect 18236 17748 18288 17800
rect 20536 17791 20588 17800
rect 20536 17757 20545 17791
rect 20545 17757 20579 17791
rect 20579 17757 20588 17791
rect 20536 17748 20588 17757
rect 22744 17748 22796 17800
rect 23940 17748 23992 17800
rect 10315 17646 10367 17698
rect 10379 17646 10431 17698
rect 10443 17646 10495 17698
rect 10507 17646 10559 17698
rect 19648 17646 19700 17698
rect 19712 17646 19764 17698
rect 19776 17646 19828 17698
rect 19840 17646 19892 17698
rect 13544 17544 13596 17596
rect 18604 17587 18656 17596
rect 18604 17553 18613 17587
rect 18613 17553 18647 17587
rect 18647 17553 18656 17587
rect 18604 17544 18656 17553
rect 20720 17544 20772 17596
rect 21916 17544 21968 17596
rect 22468 17587 22520 17596
rect 22468 17553 22477 17587
rect 22477 17553 22511 17587
rect 22511 17553 22520 17587
rect 22468 17544 22520 17553
rect 22744 17587 22796 17596
rect 22744 17553 22753 17587
rect 22753 17553 22787 17587
rect 22787 17553 22796 17587
rect 22744 17544 22796 17553
rect 23388 17544 23440 17596
rect 23940 17587 23992 17596
rect 23940 17553 23949 17587
rect 23949 17553 23983 17587
rect 23983 17553 23992 17587
rect 23940 17544 23992 17553
rect 25780 17544 25832 17596
rect 15108 17476 15160 17528
rect 18236 17519 18288 17528
rect 18236 17485 18245 17519
rect 18245 17485 18279 17519
rect 18279 17485 18288 17519
rect 18236 17476 18288 17485
rect 20352 17476 20404 17528
rect 20904 17519 20956 17528
rect 20904 17485 20913 17519
rect 20913 17485 20947 17519
rect 20947 17485 20956 17519
rect 20904 17476 20956 17485
rect 21824 17519 21876 17528
rect 21824 17485 21833 17519
rect 21833 17485 21867 17519
rect 21867 17485 21876 17519
rect 21824 17476 21876 17485
rect 13820 17408 13872 17460
rect 14372 17408 14424 17460
rect 20168 17451 20220 17460
rect 20168 17417 20177 17451
rect 20177 17417 20211 17451
rect 20211 17417 20220 17451
rect 20168 17408 20220 17417
rect 24768 17408 24820 17460
rect 19156 17340 19208 17392
rect 20260 17383 20312 17392
rect 20260 17349 20269 17383
rect 20269 17349 20303 17383
rect 20303 17349 20312 17383
rect 20260 17340 20312 17349
rect 20352 17383 20404 17392
rect 20352 17349 20361 17383
rect 20361 17349 20395 17383
rect 20395 17349 20404 17383
rect 20352 17340 20404 17349
rect 21732 17340 21784 17392
rect 24032 17340 24084 17392
rect 20996 17272 21048 17324
rect 11152 17247 11204 17256
rect 11152 17213 11161 17247
rect 11161 17213 11195 17247
rect 11195 17213 11204 17247
rect 11152 17204 11204 17213
rect 14188 17204 14240 17256
rect 15844 17204 15896 17256
rect 17316 17204 17368 17256
rect 21364 17247 21416 17256
rect 21364 17213 21373 17247
rect 21373 17213 21407 17247
rect 21407 17213 21416 17247
rect 21364 17204 21416 17213
rect 5648 17102 5700 17154
rect 5712 17102 5764 17154
rect 5776 17102 5828 17154
rect 5840 17102 5892 17154
rect 14982 17102 15034 17154
rect 15046 17102 15098 17154
rect 15110 17102 15162 17154
rect 15174 17102 15226 17154
rect 24315 17102 24367 17154
rect 24379 17102 24431 17154
rect 24443 17102 24495 17154
rect 24507 17102 24559 17154
rect 14648 17000 14700 17052
rect 11152 16932 11204 16984
rect 13636 16864 13688 16916
rect 14280 16907 14332 16916
rect 14280 16873 14289 16907
rect 14289 16873 14323 16907
rect 14323 16873 14332 16907
rect 14280 16864 14332 16873
rect 14372 16864 14424 16916
rect 17316 17000 17368 17052
rect 19156 17043 19208 17052
rect 19156 17009 19165 17043
rect 19165 17009 19199 17043
rect 19199 17009 19208 17043
rect 19156 17000 19208 17009
rect 20168 17000 20220 17052
rect 20260 17000 20312 17052
rect 23480 17000 23532 17052
rect 24032 17043 24084 17052
rect 24032 17009 24041 17043
rect 24041 17009 24075 17043
rect 24075 17009 24084 17043
rect 24032 17000 24084 17009
rect 15844 16907 15896 16916
rect 15844 16873 15853 16907
rect 15853 16873 15887 16907
rect 15887 16873 15896 16907
rect 15844 16864 15896 16873
rect 16948 16864 17000 16916
rect 20076 16864 20128 16916
rect 23204 16907 23256 16916
rect 23204 16873 23213 16907
rect 23213 16873 23247 16907
rect 23247 16873 23256 16907
rect 23204 16864 23256 16873
rect 26240 16932 26292 16984
rect 27528 16932 27580 16984
rect 15752 16839 15804 16848
rect 15752 16805 15761 16839
rect 15761 16805 15795 16839
rect 15795 16805 15804 16839
rect 15752 16796 15804 16805
rect 16856 16796 16908 16848
rect 20720 16839 20772 16848
rect 20720 16805 20729 16839
rect 20729 16805 20763 16839
rect 20763 16805 20772 16839
rect 20720 16796 20772 16805
rect 20904 16796 20956 16848
rect 21640 16796 21692 16848
rect 23388 16796 23440 16848
rect 15660 16771 15712 16780
rect 13820 16660 13872 16712
rect 15660 16737 15669 16771
rect 15669 16737 15703 16771
rect 15703 16737 15712 16771
rect 15660 16728 15712 16737
rect 22744 16728 22796 16780
rect 23848 16728 23900 16780
rect 16948 16703 17000 16712
rect 16948 16669 16957 16703
rect 16957 16669 16991 16703
rect 16991 16669 17000 16703
rect 16948 16660 17000 16669
rect 19432 16703 19484 16712
rect 19432 16669 19441 16703
rect 19441 16669 19475 16703
rect 19475 16669 19484 16703
rect 19432 16660 19484 16669
rect 21732 16660 21784 16712
rect 23204 16660 23256 16712
rect 24768 16728 24820 16780
rect 24584 16703 24636 16712
rect 24584 16669 24593 16703
rect 24593 16669 24627 16703
rect 24627 16669 24636 16703
rect 24584 16660 24636 16669
rect 10315 16558 10367 16610
rect 10379 16558 10431 16610
rect 10443 16558 10495 16610
rect 10507 16558 10559 16610
rect 19648 16558 19700 16610
rect 19712 16558 19764 16610
rect 19776 16558 19828 16610
rect 19840 16558 19892 16610
rect 13636 16499 13688 16508
rect 13636 16465 13645 16499
rect 13645 16465 13679 16499
rect 13679 16465 13688 16499
rect 13636 16456 13688 16465
rect 14280 16456 14332 16508
rect 15844 16456 15896 16508
rect 16856 16456 16908 16508
rect 17960 16456 18012 16508
rect 19432 16456 19484 16508
rect 20352 16456 20404 16508
rect 21732 16456 21784 16508
rect 21916 16499 21968 16508
rect 21916 16465 21925 16499
rect 21925 16465 21959 16499
rect 21959 16465 21968 16499
rect 21916 16456 21968 16465
rect 23664 16456 23716 16508
rect 24768 16499 24820 16508
rect 24768 16465 24777 16499
rect 24777 16465 24811 16499
rect 24811 16465 24820 16499
rect 24768 16456 24820 16465
rect 25412 16499 25464 16508
rect 25412 16465 25421 16499
rect 25421 16465 25455 16499
rect 25455 16465 25464 16499
rect 25412 16456 25464 16465
rect 14188 16388 14240 16440
rect 14464 16388 14516 16440
rect 20076 16388 20128 16440
rect 21824 16388 21876 16440
rect 24124 16388 24176 16440
rect 24584 16388 24636 16440
rect 23480 16320 23532 16372
rect 23940 16320 23992 16372
rect 19616 16295 19668 16304
rect 19616 16261 19625 16295
rect 19625 16261 19659 16295
rect 19659 16261 19668 16295
rect 19616 16252 19668 16261
rect 22100 16252 22152 16304
rect 24860 16320 24912 16372
rect 25228 16363 25280 16372
rect 25228 16329 25237 16363
rect 25237 16329 25271 16363
rect 25271 16329 25280 16363
rect 25228 16320 25280 16329
rect 24308 16295 24360 16304
rect 24308 16261 24317 16295
rect 24317 16261 24351 16295
rect 24351 16261 24360 16295
rect 24308 16252 24360 16261
rect 23020 16184 23072 16236
rect 23204 16159 23256 16168
rect 23204 16125 23213 16159
rect 23213 16125 23247 16159
rect 23247 16125 23256 16159
rect 23204 16116 23256 16125
rect 23664 16159 23716 16168
rect 23664 16125 23673 16159
rect 23673 16125 23707 16159
rect 23707 16125 23716 16159
rect 23664 16116 23716 16125
rect 5648 16014 5700 16066
rect 5712 16014 5764 16066
rect 5776 16014 5828 16066
rect 5840 16014 5892 16066
rect 14982 16014 15034 16066
rect 15046 16014 15098 16066
rect 15110 16014 15162 16066
rect 15174 16014 15226 16066
rect 24315 16014 24367 16066
rect 24379 16014 24431 16066
rect 24443 16014 24495 16066
rect 24507 16014 24559 16066
rect 14188 15912 14240 15964
rect 14464 15912 14516 15964
rect 16948 15912 17000 15964
rect 15660 15776 15712 15828
rect 17960 15912 18012 15964
rect 20076 15912 20128 15964
rect 22100 15912 22152 15964
rect 23388 15912 23440 15964
rect 24768 15912 24820 15964
rect 25044 15955 25096 15964
rect 25044 15921 25053 15955
rect 25053 15921 25087 15955
rect 25087 15921 25096 15955
rect 25044 15912 25096 15921
rect 25228 15912 25280 15964
rect 24860 15844 24912 15896
rect 11060 15708 11112 15760
rect 13820 15708 13872 15760
rect 20168 15776 20220 15828
rect 21364 15819 21416 15828
rect 21364 15785 21373 15819
rect 21373 15785 21407 15819
rect 21407 15785 21416 15819
rect 21364 15776 21416 15785
rect 23112 15819 23164 15828
rect 17684 15708 17736 15760
rect 19156 15708 19208 15760
rect 19616 15751 19668 15760
rect 19616 15717 19625 15751
rect 19625 15717 19659 15751
rect 19659 15717 19668 15751
rect 19616 15708 19668 15717
rect 23112 15785 23121 15819
rect 23121 15785 23155 15819
rect 23155 15785 23164 15819
rect 23112 15776 23164 15785
rect 17132 15640 17184 15692
rect 12256 15615 12308 15624
rect 12256 15581 12265 15615
rect 12265 15581 12299 15615
rect 12299 15581 12308 15615
rect 12256 15572 12308 15581
rect 14372 15615 14424 15624
rect 14372 15581 14381 15615
rect 14381 15581 14415 15615
rect 14415 15581 14424 15615
rect 14372 15572 14424 15581
rect 20628 15615 20680 15624
rect 20628 15581 20637 15615
rect 20637 15581 20671 15615
rect 20671 15581 20680 15615
rect 20628 15572 20680 15581
rect 20996 15572 21048 15624
rect 23204 15640 23256 15692
rect 24308 15640 24360 15692
rect 22100 15572 22152 15624
rect 10315 15470 10367 15522
rect 10379 15470 10431 15522
rect 10443 15470 10495 15522
rect 10507 15470 10559 15522
rect 19648 15470 19700 15522
rect 19712 15470 19764 15522
rect 19776 15470 19828 15522
rect 19840 15470 19892 15522
rect 12532 15368 12584 15420
rect 14740 15368 14792 15420
rect 17132 15411 17184 15420
rect 17132 15377 17141 15411
rect 17141 15377 17175 15411
rect 17175 15377 17184 15411
rect 17132 15368 17184 15377
rect 20628 15368 20680 15420
rect 21364 15368 21416 15420
rect 23020 15368 23072 15420
rect 23664 15368 23716 15420
rect 24676 15411 24728 15420
rect 24676 15377 24685 15411
rect 24685 15377 24719 15411
rect 24719 15377 24728 15411
rect 24676 15368 24728 15377
rect 25412 15411 25464 15420
rect 25412 15377 25421 15411
rect 25421 15377 25455 15411
rect 25455 15377 25464 15411
rect 25412 15368 25464 15377
rect 23480 15300 23532 15352
rect 24032 15343 24084 15352
rect 24032 15309 24041 15343
rect 24041 15309 24075 15343
rect 24075 15309 24084 15343
rect 24032 15300 24084 15309
rect 12440 15275 12492 15284
rect 12440 15241 12449 15275
rect 12449 15241 12483 15275
rect 12483 15241 12492 15275
rect 14648 15275 14700 15284
rect 12440 15232 12492 15241
rect 14648 15241 14657 15275
rect 14657 15241 14691 15275
rect 14691 15241 14700 15275
rect 14648 15232 14700 15241
rect 19156 15275 19208 15284
rect 19156 15241 19165 15275
rect 19165 15241 19199 15275
rect 19199 15241 19208 15275
rect 19156 15232 19208 15241
rect 19432 15275 19484 15284
rect 19432 15241 19466 15275
rect 19466 15241 19484 15275
rect 19432 15232 19484 15241
rect 25136 15232 25188 15284
rect 24308 15207 24360 15216
rect 24308 15173 24317 15207
rect 24317 15173 24351 15207
rect 24351 15173 24360 15207
rect 24308 15164 24360 15173
rect 24768 15164 24820 15216
rect 24124 15096 24176 15148
rect 13452 15028 13504 15080
rect 15844 15028 15896 15080
rect 5648 14926 5700 14978
rect 5712 14926 5764 14978
rect 5776 14926 5828 14978
rect 5840 14926 5892 14978
rect 14982 14926 15034 14978
rect 15046 14926 15098 14978
rect 15110 14926 15162 14978
rect 15174 14926 15226 14978
rect 24315 14926 24367 14978
rect 24379 14926 24431 14978
rect 24443 14926 24495 14978
rect 24507 14926 24559 14978
rect 12440 14824 12492 14876
rect 17224 14867 17276 14876
rect 17224 14833 17233 14867
rect 17233 14833 17267 14867
rect 17267 14833 17276 14867
rect 17224 14824 17276 14833
rect 19156 14867 19208 14876
rect 19156 14833 19165 14867
rect 19165 14833 19199 14867
rect 19199 14833 19208 14867
rect 19156 14824 19208 14833
rect 19432 14824 19484 14876
rect 21548 14824 21600 14876
rect 23572 14824 23624 14876
rect 24676 14824 24728 14876
rect 25136 14824 25188 14876
rect 14648 14756 14700 14808
rect 24032 14799 24084 14808
rect 24032 14765 24041 14799
rect 24041 14765 24075 14799
rect 24075 14765 24084 14799
rect 24032 14756 24084 14765
rect 24216 14756 24268 14808
rect 13452 14731 13504 14740
rect 13452 14697 13461 14731
rect 13461 14697 13495 14731
rect 13495 14697 13504 14731
rect 13452 14688 13504 14697
rect 15844 14731 15896 14740
rect 15844 14697 15853 14731
rect 15853 14697 15887 14731
rect 15887 14697 15896 14731
rect 15844 14688 15896 14697
rect 23664 14688 23716 14740
rect 25044 14688 25096 14740
rect 18052 14663 18104 14672
rect 12716 14552 12768 14604
rect 16212 14552 16264 14604
rect 18052 14629 18061 14663
rect 18061 14629 18095 14663
rect 18095 14629 18104 14663
rect 18052 14620 18104 14629
rect 20996 14620 21048 14672
rect 23756 14620 23808 14672
rect 24032 14620 24084 14672
rect 24768 14620 24820 14672
rect 22928 14595 22980 14604
rect 22928 14561 22937 14595
rect 22937 14561 22971 14595
rect 22971 14561 22980 14595
rect 22928 14552 22980 14561
rect 26148 14552 26200 14604
rect 12900 14484 12952 14536
rect 15476 14484 15528 14536
rect 17592 14527 17644 14536
rect 17592 14493 17601 14527
rect 17601 14493 17635 14527
rect 17635 14493 17644 14527
rect 17592 14484 17644 14493
rect 18236 14527 18288 14536
rect 18236 14493 18245 14527
rect 18245 14493 18279 14527
rect 18279 14493 18288 14527
rect 18236 14484 18288 14493
rect 23756 14484 23808 14536
rect 24492 14527 24544 14536
rect 24492 14493 24501 14527
rect 24501 14493 24535 14527
rect 24535 14493 24544 14527
rect 24492 14484 24544 14493
rect 24860 14484 24912 14536
rect 10315 14382 10367 14434
rect 10379 14382 10431 14434
rect 10443 14382 10495 14434
rect 10507 14382 10559 14434
rect 19648 14382 19700 14434
rect 19712 14382 19764 14434
rect 19776 14382 19828 14434
rect 19840 14382 19892 14434
rect 12716 14323 12768 14332
rect 12716 14289 12725 14323
rect 12725 14289 12759 14323
rect 12759 14289 12768 14323
rect 12716 14280 12768 14289
rect 16212 14323 16264 14332
rect 16212 14289 16221 14323
rect 16221 14289 16255 14323
rect 16255 14289 16264 14323
rect 16212 14280 16264 14289
rect 17592 14280 17644 14332
rect 20996 14323 21048 14332
rect 20996 14289 21005 14323
rect 21005 14289 21039 14323
rect 21039 14289 21048 14323
rect 20996 14280 21048 14289
rect 24492 14280 24544 14332
rect 13452 14212 13504 14264
rect 23020 14212 23072 14264
rect 23572 14212 23624 14264
rect 13360 14144 13412 14196
rect 14464 14144 14516 14196
rect 18052 14144 18104 14196
rect 21364 14187 21416 14196
rect 21364 14153 21373 14187
rect 21373 14153 21407 14187
rect 21407 14153 21416 14187
rect 21364 14144 21416 14153
rect 22100 14144 22152 14196
rect 22928 14144 22980 14196
rect 23112 14144 23164 14196
rect 18512 14119 18564 14128
rect 18512 14085 18521 14119
rect 18521 14085 18555 14119
rect 18555 14085 18564 14119
rect 18512 14076 18564 14085
rect 18604 14119 18656 14128
rect 18604 14085 18613 14119
rect 18613 14085 18647 14119
rect 18647 14085 18656 14119
rect 21456 14119 21508 14128
rect 18604 14076 18656 14085
rect 21456 14085 21465 14119
rect 21465 14085 21499 14119
rect 21499 14085 21508 14119
rect 21456 14076 21508 14085
rect 21640 14119 21692 14128
rect 21640 14085 21649 14119
rect 21649 14085 21683 14119
rect 21683 14085 21692 14119
rect 21640 14076 21692 14085
rect 22376 14008 22428 14060
rect 15384 13940 15436 13992
rect 23480 13940 23532 13992
rect 5648 13838 5700 13890
rect 5712 13838 5764 13890
rect 5776 13838 5828 13890
rect 5840 13838 5892 13890
rect 14982 13838 15034 13890
rect 15046 13838 15098 13890
rect 15110 13838 15162 13890
rect 15174 13838 15226 13890
rect 24315 13838 24367 13890
rect 24379 13838 24431 13890
rect 24443 13838 24495 13890
rect 24507 13838 24559 13890
rect 12072 13736 12124 13788
rect 13360 13736 13412 13788
rect 13452 13736 13504 13788
rect 15936 13736 15988 13788
rect 14464 13668 14516 13720
rect 11704 13575 11756 13584
rect 11704 13541 11713 13575
rect 11713 13541 11747 13575
rect 11747 13541 11756 13575
rect 11704 13532 11756 13541
rect 12072 13575 12124 13584
rect 12072 13541 12081 13575
rect 12081 13541 12115 13575
rect 12115 13541 12124 13575
rect 12072 13532 12124 13541
rect 18052 13736 18104 13788
rect 21364 13736 21416 13788
rect 17684 13711 17736 13720
rect 17684 13677 17693 13711
rect 17693 13677 17727 13711
rect 17727 13677 17736 13711
rect 17684 13668 17736 13677
rect 23112 13736 23164 13788
rect 24860 13779 24912 13788
rect 24860 13745 24869 13779
rect 24869 13745 24903 13779
rect 24903 13745 24912 13779
rect 24860 13736 24912 13745
rect 23572 13711 23624 13720
rect 23572 13677 23581 13711
rect 23581 13677 23615 13711
rect 23615 13677 23624 13711
rect 23572 13668 23624 13677
rect 13636 13532 13688 13584
rect 15384 13532 15436 13584
rect 17684 13532 17736 13584
rect 17868 13532 17920 13584
rect 21456 13532 21508 13584
rect 24584 13532 24636 13584
rect 21640 13464 21692 13516
rect 22376 13464 22428 13516
rect 19156 13439 19208 13448
rect 19156 13405 19165 13439
rect 19165 13405 19199 13439
rect 19199 13405 19208 13439
rect 19156 13396 19208 13405
rect 10315 13294 10367 13346
rect 10379 13294 10431 13346
rect 10443 13294 10495 13346
rect 10507 13294 10559 13346
rect 19648 13294 19700 13346
rect 19712 13294 19764 13346
rect 19776 13294 19828 13346
rect 19840 13294 19892 13346
rect 2780 13235 2832 13244
rect 2780 13201 2789 13235
rect 2789 13201 2823 13235
rect 2823 13201 2832 13235
rect 2780 13192 2832 13201
rect 12900 13235 12952 13244
rect 12900 13201 12909 13235
rect 12909 13201 12943 13235
rect 12943 13201 12952 13235
rect 12900 13192 12952 13201
rect 15476 13235 15528 13244
rect 15476 13201 15485 13235
rect 15485 13201 15519 13235
rect 15519 13201 15528 13235
rect 15476 13192 15528 13201
rect 17868 13235 17920 13244
rect 17868 13201 17877 13235
rect 17877 13201 17911 13235
rect 17911 13201 17920 13235
rect 17868 13192 17920 13201
rect 18052 13235 18104 13244
rect 18052 13201 18061 13235
rect 18061 13201 18095 13235
rect 18095 13201 18104 13235
rect 18052 13192 18104 13201
rect 18512 13192 18564 13244
rect 18696 13192 18748 13244
rect 21456 13192 21508 13244
rect 22928 13235 22980 13244
rect 22928 13201 22937 13235
rect 22937 13201 22971 13235
rect 22971 13201 22980 13235
rect 22928 13192 22980 13201
rect 24768 13235 24820 13244
rect 24768 13201 24777 13235
rect 24777 13201 24811 13235
rect 24811 13201 24820 13235
rect 24768 13192 24820 13201
rect 2044 13124 2096 13176
rect 15384 13167 15436 13176
rect 15384 13133 15393 13167
rect 15393 13133 15427 13167
rect 15427 13133 15436 13167
rect 18604 13167 18656 13176
rect 15384 13124 15436 13133
rect 1492 13056 1544 13108
rect 13268 13099 13320 13108
rect 13268 13065 13277 13099
rect 13277 13065 13311 13099
rect 13311 13065 13320 13099
rect 13268 13056 13320 13065
rect 15844 13099 15896 13108
rect 15844 13065 15853 13099
rect 15853 13065 15887 13099
rect 15887 13065 15896 13099
rect 15844 13056 15896 13065
rect 13360 13031 13412 13040
rect 13360 12997 13369 13031
rect 13369 12997 13403 13031
rect 13403 12997 13412 13031
rect 13360 12988 13412 12997
rect 13636 12988 13688 13040
rect 15936 13031 15988 13040
rect 15936 12997 15945 13031
rect 15945 12997 15979 13031
rect 15979 12997 15988 13031
rect 15936 12988 15988 12997
rect 18604 13133 18613 13167
rect 18613 13133 18647 13167
rect 18647 13133 18656 13167
rect 18604 13124 18656 13133
rect 19432 13124 19484 13176
rect 22192 13056 22244 13108
rect 24584 13099 24636 13108
rect 24584 13065 24593 13099
rect 24593 13065 24627 13099
rect 24627 13065 24636 13099
rect 24584 13056 24636 13065
rect 16212 12988 16264 13040
rect 19248 12988 19300 13040
rect 22468 13031 22520 13040
rect 22468 12997 22477 13031
rect 22477 12997 22511 13031
rect 22511 12997 22520 13031
rect 22468 12988 22520 12997
rect 22284 12920 22336 12972
rect 20812 12895 20864 12904
rect 20812 12861 20821 12895
rect 20821 12861 20855 12895
rect 20855 12861 20864 12895
rect 20812 12852 20864 12861
rect 5648 12750 5700 12802
rect 5712 12750 5764 12802
rect 5776 12750 5828 12802
rect 5840 12750 5892 12802
rect 14982 12750 15034 12802
rect 15046 12750 15098 12802
rect 15110 12750 15162 12802
rect 15174 12750 15226 12802
rect 24315 12750 24367 12802
rect 24379 12750 24431 12802
rect 24443 12750 24495 12802
rect 24507 12750 24559 12802
rect 1492 12648 1544 12700
rect 2044 12691 2096 12700
rect 2044 12657 2053 12691
rect 2053 12657 2087 12691
rect 2087 12657 2096 12691
rect 2044 12648 2096 12657
rect 13268 12648 13320 12700
rect 13636 12691 13688 12700
rect 13636 12657 13645 12691
rect 13645 12657 13679 12691
rect 13679 12657 13688 12691
rect 13636 12648 13688 12657
rect 15844 12648 15896 12700
rect 16212 12691 16264 12700
rect 16212 12657 16221 12691
rect 16221 12657 16255 12691
rect 16255 12657 16264 12691
rect 16212 12648 16264 12657
rect 18052 12648 18104 12700
rect 19248 12648 19300 12700
rect 19432 12691 19484 12700
rect 19432 12657 19441 12691
rect 19441 12657 19475 12691
rect 19475 12657 19484 12691
rect 19432 12648 19484 12657
rect 22376 12648 22428 12700
rect 23664 12691 23716 12700
rect 23664 12657 23673 12691
rect 23673 12657 23707 12691
rect 23707 12657 23716 12691
rect 23664 12648 23716 12657
rect 24676 12648 24728 12700
rect 24768 12623 24820 12632
rect 24768 12589 24777 12623
rect 24777 12589 24811 12623
rect 24811 12589 24820 12623
rect 24768 12580 24820 12589
rect 13360 12487 13412 12496
rect 13360 12453 13369 12487
rect 13369 12453 13403 12487
rect 13403 12453 13412 12487
rect 13360 12444 13412 12453
rect 15936 12487 15988 12496
rect 15936 12453 15945 12487
rect 15945 12453 15979 12487
rect 15979 12453 15988 12487
rect 15936 12444 15988 12453
rect 18052 12487 18104 12496
rect 18052 12453 18061 12487
rect 18061 12453 18095 12487
rect 18095 12453 18104 12487
rect 18052 12444 18104 12453
rect 19156 12444 19208 12496
rect 20812 12444 20864 12496
rect 22468 12444 22520 12496
rect 23480 12487 23532 12496
rect 23480 12453 23489 12487
rect 23489 12453 23523 12487
rect 23523 12453 23532 12487
rect 23480 12444 23532 12453
rect 23480 12308 23532 12360
rect 10315 12206 10367 12258
rect 10379 12206 10431 12258
rect 10443 12206 10495 12258
rect 10507 12206 10559 12258
rect 19648 12206 19700 12258
rect 19712 12206 19764 12258
rect 19776 12206 19828 12258
rect 19840 12206 19892 12258
rect 18696 12104 18748 12156
rect 19432 12147 19484 12156
rect 19432 12113 19441 12147
rect 19441 12113 19475 12147
rect 19475 12113 19484 12147
rect 19432 12104 19484 12113
rect 20812 12104 20864 12156
rect 22284 12147 22336 12156
rect 22284 12113 22293 12147
rect 22293 12113 22327 12147
rect 22327 12113 22336 12147
rect 22284 12104 22336 12113
rect 23480 12104 23532 12156
rect 24768 12147 24820 12156
rect 24768 12113 24777 12147
rect 24777 12113 24811 12147
rect 24811 12113 24820 12147
rect 24768 12104 24820 12113
rect 18328 11968 18380 12020
rect 22100 11968 22152 12020
rect 22560 12011 22612 12020
rect 22560 11977 22569 12011
rect 22569 11977 22603 12011
rect 22603 11977 22612 12011
rect 22560 11968 22612 11977
rect 24676 11968 24728 12020
rect 18512 11900 18564 11952
rect 19156 11900 19208 11952
rect 22008 11943 22060 11952
rect 22008 11909 22017 11943
rect 22017 11909 22051 11943
rect 22051 11909 22060 11943
rect 22008 11900 22060 11909
rect 5648 11662 5700 11714
rect 5712 11662 5764 11714
rect 5776 11662 5828 11714
rect 5840 11662 5892 11714
rect 14982 11662 15034 11714
rect 15046 11662 15098 11714
rect 15110 11662 15162 11714
rect 15174 11662 15226 11714
rect 24315 11662 24367 11714
rect 24379 11662 24431 11714
rect 24443 11662 24495 11714
rect 24507 11662 24559 11714
rect 18512 11560 18564 11612
rect 19156 11560 19208 11612
rect 22560 11603 22612 11612
rect 22560 11569 22569 11603
rect 22569 11569 22603 11603
rect 22603 11569 22612 11603
rect 22560 11560 22612 11569
rect 24676 11560 24728 11612
rect 24768 11603 24820 11612
rect 24768 11569 24777 11603
rect 24777 11569 24811 11603
rect 24811 11569 24820 11603
rect 24768 11560 24820 11569
rect 23848 11492 23900 11544
rect 25228 11467 25280 11476
rect 25228 11433 25237 11467
rect 25237 11433 25271 11467
rect 25271 11433 25280 11467
rect 25228 11424 25280 11433
rect 18328 11263 18380 11272
rect 18328 11229 18337 11263
rect 18337 11229 18371 11263
rect 18371 11229 18380 11263
rect 18328 11220 18380 11229
rect 10315 11118 10367 11170
rect 10379 11118 10431 11170
rect 10443 11118 10495 11170
rect 10507 11118 10559 11170
rect 19648 11118 19700 11170
rect 19712 11118 19764 11170
rect 19776 11118 19828 11170
rect 19840 11118 19892 11170
rect 23756 11016 23808 11068
rect 24584 10923 24636 10932
rect 24584 10889 24593 10923
rect 24593 10889 24627 10923
rect 24627 10889 24636 10923
rect 24584 10880 24636 10889
rect 5648 10574 5700 10626
rect 5712 10574 5764 10626
rect 5776 10574 5828 10626
rect 5840 10574 5892 10626
rect 14982 10574 15034 10626
rect 15046 10574 15098 10626
rect 15110 10574 15162 10626
rect 15174 10574 15226 10626
rect 24315 10574 24367 10626
rect 24379 10574 24431 10626
rect 24443 10574 24495 10626
rect 24507 10574 24559 10626
rect 24768 10515 24820 10524
rect 24768 10481 24777 10515
rect 24777 10481 24811 10515
rect 24811 10481 24820 10515
rect 24768 10472 24820 10481
rect 24676 10404 24728 10456
rect 25228 10243 25280 10252
rect 25228 10209 25237 10243
rect 25237 10209 25271 10243
rect 25271 10209 25280 10243
rect 25228 10200 25280 10209
rect 10315 10030 10367 10082
rect 10379 10030 10431 10082
rect 10443 10030 10495 10082
rect 10507 10030 10559 10082
rect 19648 10030 19700 10082
rect 19712 10030 19764 10082
rect 19776 10030 19828 10082
rect 19840 10030 19892 10082
rect 24032 9928 24084 9980
rect 24584 9835 24636 9844
rect 24584 9801 24593 9835
rect 24593 9801 24627 9835
rect 24627 9801 24636 9835
rect 24584 9792 24636 9801
rect 5648 9486 5700 9538
rect 5712 9486 5764 9538
rect 5776 9486 5828 9538
rect 5840 9486 5892 9538
rect 14982 9486 15034 9538
rect 15046 9486 15098 9538
rect 15110 9486 15162 9538
rect 15174 9486 15226 9538
rect 24315 9486 24367 9538
rect 24379 9486 24431 9538
rect 24443 9486 24495 9538
rect 24507 9486 24559 9538
rect 18236 9384 18288 9436
rect 18972 9384 19024 9436
rect 24676 9427 24728 9436
rect 24676 9393 24685 9427
rect 24685 9393 24719 9427
rect 24719 9393 24728 9427
rect 24676 9384 24728 9393
rect 23940 9359 23992 9368
rect 23940 9325 23949 9359
rect 23949 9325 23983 9359
rect 23983 9325 23992 9359
rect 23940 9316 23992 9325
rect 24400 9155 24452 9164
rect 24400 9121 24409 9155
rect 24409 9121 24443 9155
rect 24443 9121 24452 9155
rect 24400 9112 24452 9121
rect 10315 8942 10367 8994
rect 10379 8942 10431 8994
rect 10443 8942 10495 8994
rect 10507 8942 10559 8994
rect 19648 8942 19700 8994
rect 19712 8942 19764 8994
rect 19776 8942 19828 8994
rect 19840 8942 19892 8994
rect 24124 8840 24176 8892
rect 24400 8747 24452 8756
rect 24400 8713 24409 8747
rect 24409 8713 24443 8747
rect 24443 8713 24452 8747
rect 24400 8704 24452 8713
rect 16488 8636 16540 8688
rect 16672 8636 16724 8688
rect 5648 8398 5700 8450
rect 5712 8398 5764 8450
rect 5776 8398 5828 8450
rect 5840 8398 5892 8450
rect 14982 8398 15034 8450
rect 15046 8398 15098 8450
rect 15110 8398 15162 8450
rect 15174 8398 15226 8450
rect 24315 8398 24367 8450
rect 24379 8398 24431 8450
rect 24443 8398 24495 8450
rect 24507 8398 24559 8450
rect 24676 8296 24728 8348
rect 10315 7854 10367 7906
rect 10379 7854 10431 7906
rect 10443 7854 10495 7906
rect 10507 7854 10559 7906
rect 19648 7854 19700 7906
rect 19712 7854 19764 7906
rect 19776 7854 19828 7906
rect 19840 7854 19892 7906
rect 23480 7752 23532 7804
rect 24676 7616 24728 7668
rect 5648 7310 5700 7362
rect 5712 7310 5764 7362
rect 5776 7310 5828 7362
rect 5840 7310 5892 7362
rect 14982 7310 15034 7362
rect 15046 7310 15098 7362
rect 15110 7310 15162 7362
rect 15174 7310 15226 7362
rect 24315 7310 24367 7362
rect 24379 7310 24431 7362
rect 24443 7310 24495 7362
rect 24507 7310 24559 7362
rect 21180 7251 21232 7260
rect 21180 7217 21189 7251
rect 21189 7217 21223 7251
rect 21223 7217 21232 7251
rect 21180 7208 21232 7217
rect 24676 7251 24728 7260
rect 24676 7217 24685 7251
rect 24685 7217 24719 7251
rect 24719 7217 24728 7251
rect 24676 7208 24728 7217
rect 21640 6911 21692 6920
rect 21640 6877 21649 6911
rect 21649 6877 21683 6911
rect 21683 6877 21692 6911
rect 21640 6868 21692 6877
rect 10315 6766 10367 6818
rect 10379 6766 10431 6818
rect 10443 6766 10495 6818
rect 10507 6766 10559 6818
rect 19648 6766 19700 6818
rect 19712 6766 19764 6818
rect 19776 6766 19828 6818
rect 19840 6766 19892 6818
rect 20352 6571 20404 6580
rect 20352 6537 20361 6571
rect 20361 6537 20395 6571
rect 20395 6537 20404 6571
rect 20352 6528 20404 6537
rect 21272 6392 21324 6444
rect 5648 6222 5700 6274
rect 5712 6222 5764 6274
rect 5776 6222 5828 6274
rect 5840 6222 5892 6274
rect 14982 6222 15034 6274
rect 15046 6222 15098 6274
rect 15110 6222 15162 6274
rect 15174 6222 15226 6274
rect 24315 6222 24367 6274
rect 24379 6222 24431 6274
rect 24443 6222 24495 6274
rect 24507 6222 24559 6274
rect 19984 6120 20036 6172
rect 20352 6163 20404 6172
rect 20352 6129 20361 6163
rect 20361 6129 20395 6163
rect 20395 6129 20404 6163
rect 20352 6120 20404 6129
rect 20076 5780 20128 5832
rect 10315 5678 10367 5730
rect 10379 5678 10431 5730
rect 10443 5678 10495 5730
rect 10507 5678 10559 5730
rect 19648 5678 19700 5730
rect 19712 5678 19764 5730
rect 19776 5678 19828 5730
rect 19840 5678 19892 5730
rect 5648 5134 5700 5186
rect 5712 5134 5764 5186
rect 5776 5134 5828 5186
rect 5840 5134 5892 5186
rect 14982 5134 15034 5186
rect 15046 5134 15098 5186
rect 15110 5134 15162 5186
rect 15174 5134 15226 5186
rect 24315 5134 24367 5186
rect 24379 5134 24431 5186
rect 24443 5134 24495 5186
rect 24507 5134 24559 5186
rect 23480 5032 23532 5084
rect 25228 5075 25280 5084
rect 25228 5041 25237 5075
rect 25237 5041 25271 5075
rect 25271 5041 25280 5075
rect 25228 5032 25280 5041
rect 25228 4828 25280 4880
rect 10315 4590 10367 4642
rect 10379 4590 10431 4642
rect 10443 4590 10495 4642
rect 10507 4590 10559 4642
rect 19648 4590 19700 4642
rect 19712 4590 19764 4642
rect 19776 4590 19828 4642
rect 19840 4590 19892 4642
rect 24768 4531 24820 4540
rect 24768 4497 24777 4531
rect 24777 4497 24811 4531
rect 24811 4497 24820 4531
rect 24768 4488 24820 4497
rect 24584 4395 24636 4404
rect 24584 4361 24593 4395
rect 24593 4361 24627 4395
rect 24627 4361 24636 4395
rect 24584 4352 24636 4361
rect 5648 4046 5700 4098
rect 5712 4046 5764 4098
rect 5776 4046 5828 4098
rect 5840 4046 5892 4098
rect 14982 4046 15034 4098
rect 15046 4046 15098 4098
rect 15110 4046 15162 4098
rect 15174 4046 15226 4098
rect 24315 4046 24367 4098
rect 24379 4046 24431 4098
rect 24443 4046 24495 4098
rect 24507 4046 24559 4098
rect 24676 3944 24728 3996
rect 25228 3851 25280 3860
rect 25228 3817 25237 3851
rect 25237 3817 25271 3851
rect 25271 3817 25280 3851
rect 25228 3808 25280 3817
rect 24768 3647 24820 3656
rect 24768 3613 24777 3647
rect 24777 3613 24811 3647
rect 24811 3613 24820 3647
rect 24768 3604 24820 3613
rect 10315 3502 10367 3554
rect 10379 3502 10431 3554
rect 10443 3502 10495 3554
rect 10507 3502 10559 3554
rect 19648 3502 19700 3554
rect 19712 3502 19764 3554
rect 19776 3502 19828 3554
rect 19840 3502 19892 3554
rect 5648 2958 5700 3010
rect 5712 2958 5764 3010
rect 5776 2958 5828 3010
rect 5840 2958 5892 3010
rect 14982 2958 15034 3010
rect 15046 2958 15098 3010
rect 15110 2958 15162 3010
rect 15174 2958 15226 3010
rect 24315 2958 24367 3010
rect 24379 2958 24431 3010
rect 24443 2958 24495 3010
rect 24507 2958 24559 3010
rect 16488 2856 16540 2908
rect 24768 2899 24820 2908
rect 24768 2865 24777 2899
rect 24777 2865 24811 2899
rect 24811 2865 24820 2899
rect 24768 2856 24820 2865
rect 16764 2763 16816 2772
rect 16764 2729 16773 2763
rect 16773 2729 16807 2763
rect 16807 2729 16816 2763
rect 16764 2720 16816 2729
rect 24676 2652 24728 2704
rect 10315 2414 10367 2466
rect 10379 2414 10431 2466
rect 10443 2414 10495 2466
rect 10507 2414 10559 2466
rect 19648 2414 19700 2466
rect 19712 2414 19764 2466
rect 19776 2414 19828 2466
rect 19840 2414 19892 2466
rect 25228 2176 25280 2228
rect 24768 2083 24820 2092
rect 24768 2049 24777 2083
rect 24777 2049 24811 2083
rect 24811 2049 24820 2083
rect 24768 2040 24820 2049
rect 25228 2015 25280 2024
rect 25228 1981 25237 2015
rect 25237 1981 25271 2015
rect 25271 1981 25280 2015
rect 25228 1972 25280 1981
rect 5648 1870 5700 1922
rect 5712 1870 5764 1922
rect 5776 1870 5828 1922
rect 5840 1870 5892 1922
rect 14982 1870 15034 1922
rect 15046 1870 15098 1922
rect 15110 1870 15162 1922
rect 15174 1870 15226 1922
rect 24315 1870 24367 1922
rect 24379 1870 24431 1922
rect 24443 1870 24495 1922
rect 24507 1870 24559 1922
<< metal2 >>
rect 294 27240 350 27720
rect 938 27240 994 27720
rect 1582 27240 1638 27720
rect 2318 27240 2374 27720
rect 2962 27240 3018 27720
rect 3698 27240 3754 27720
rect 4342 27240 4398 27720
rect 4986 27240 5042 27720
rect 5722 27240 5778 27720
rect 6366 27240 6422 27720
rect 7102 27240 7158 27720
rect 7746 27240 7802 27720
rect 8390 27240 8446 27720
rect 9126 27240 9182 27720
rect 9770 27240 9826 27720
rect 10506 27240 10562 27720
rect 11150 27240 11206 27720
rect 11886 27240 11942 27720
rect 12530 27240 12586 27720
rect 13174 27240 13230 27720
rect 13910 27240 13966 27720
rect 14554 27240 14610 27720
rect 15290 27240 15346 27720
rect 15934 27240 15990 27720
rect 16578 27240 16634 27720
rect 17314 27240 17370 27720
rect 17958 27240 18014 27720
rect 18694 27240 18750 27720
rect 19338 27240 19394 27720
rect 20074 27240 20130 27720
rect 20718 27240 20774 27720
rect 21362 27240 21418 27720
rect 22098 27240 22154 27720
rect 22742 27240 22798 27720
rect 23478 27240 23534 27720
rect 24122 27240 24178 27720
rect 24766 27240 24822 27720
rect 25502 27240 25558 27720
rect 25870 27424 25926 27433
rect 25870 27359 25926 27368
rect 308 27138 336 27240
rect 308 27110 428 27138
rect 400 13153 428 27110
rect 952 20089 980 27240
rect 938 20080 994 20089
rect 938 20015 994 20024
rect 1596 18593 1624 27240
rect 2332 21313 2360 27240
rect 2318 21304 2374 21313
rect 2318 21239 2374 21248
rect 1582 18584 1638 18593
rect 1582 18519 1638 18528
rect 2976 17913 3004 27240
rect 3712 20225 3740 27240
rect 3698 20216 3754 20225
rect 3698 20151 3754 20160
rect 4356 19001 4384 27240
rect 5000 22401 5028 27240
rect 5736 24962 5764 27240
rect 5736 24934 6040 24962
rect 5622 24772 5918 24792
rect 5678 24770 5702 24772
rect 5758 24770 5782 24772
rect 5838 24770 5862 24772
rect 5700 24718 5702 24770
rect 5764 24718 5776 24770
rect 5838 24718 5840 24770
rect 5678 24716 5702 24718
rect 5758 24716 5782 24718
rect 5838 24716 5862 24718
rect 5622 24696 5918 24716
rect 6012 23897 6040 24934
rect 6380 24441 6408 27240
rect 6366 24432 6422 24441
rect 6366 24367 6422 24376
rect 5998 23888 6054 23897
rect 5998 23823 6054 23832
rect 5622 23684 5918 23704
rect 5678 23682 5702 23684
rect 5758 23682 5782 23684
rect 5838 23682 5862 23684
rect 5700 23630 5702 23682
rect 5764 23630 5776 23682
rect 5838 23630 5840 23682
rect 5678 23628 5702 23630
rect 5758 23628 5782 23630
rect 5838 23628 5862 23630
rect 5622 23608 5918 23628
rect 7116 23353 7144 27240
rect 7102 23344 7158 23353
rect 7102 23279 7158 23288
rect 7760 22809 7788 27240
rect 8404 22945 8432 27240
rect 8390 22936 8446 22945
rect 8390 22871 8446 22880
rect 7746 22800 7802 22809
rect 7746 22735 7802 22744
rect 5622 22596 5918 22616
rect 5678 22594 5702 22596
rect 5758 22594 5782 22596
rect 5838 22594 5862 22596
rect 5700 22542 5702 22594
rect 5764 22542 5776 22594
rect 5838 22542 5840 22594
rect 5678 22540 5702 22542
rect 5758 22540 5782 22542
rect 5838 22540 5862 22542
rect 5622 22520 5918 22540
rect 4986 22392 5042 22401
rect 4986 22327 5042 22336
rect 5622 21508 5918 21528
rect 5678 21506 5702 21508
rect 5758 21506 5782 21508
rect 5838 21506 5862 21508
rect 5700 21454 5702 21506
rect 5764 21454 5776 21506
rect 5838 21454 5840 21506
rect 5678 21452 5702 21454
rect 5758 21452 5782 21454
rect 5838 21452 5862 21454
rect 5622 21432 5918 21452
rect 9140 21410 9168 27240
rect 9784 23382 9812 27240
rect 10520 25506 10548 27240
rect 10520 25478 10824 25506
rect 10289 25316 10585 25336
rect 10345 25314 10369 25316
rect 10425 25314 10449 25316
rect 10505 25314 10529 25316
rect 10367 25262 10369 25314
rect 10431 25262 10443 25314
rect 10505 25262 10507 25314
rect 10345 25260 10369 25262
rect 10425 25260 10449 25262
rect 10505 25260 10529 25262
rect 10289 25240 10585 25260
rect 10289 24228 10585 24248
rect 10345 24226 10369 24228
rect 10425 24226 10449 24228
rect 10505 24226 10529 24228
rect 10367 24174 10369 24226
rect 10431 24174 10443 24226
rect 10505 24174 10507 24226
rect 10345 24172 10369 24174
rect 10425 24172 10449 24174
rect 10505 24172 10529 24174
rect 10289 24152 10585 24172
rect 10796 23382 10824 25478
rect 11164 23994 11192 27240
rect 11152 23988 11204 23994
rect 11152 23930 11204 23936
rect 11164 23586 11192 23930
rect 11152 23580 11204 23586
rect 11152 23522 11204 23528
rect 11900 23382 11928 27240
rect 12348 23784 12400 23790
rect 12348 23726 12400 23732
rect 9772 23376 9824 23382
rect 9772 23318 9824 23324
rect 10784 23376 10836 23382
rect 10784 23318 10836 23324
rect 11888 23376 11940 23382
rect 11888 23318 11940 23324
rect 9864 23240 9916 23246
rect 10968 23240 11020 23246
rect 9864 23182 9916 23188
rect 10966 23208 10968 23217
rect 12072 23240 12124 23246
rect 11020 23208 11022 23217
rect 9128 21404 9180 21410
rect 9128 21346 9180 21352
rect 9680 21064 9732 21070
rect 9680 21006 9732 21012
rect 9692 20730 9720 21006
rect 9680 20724 9732 20730
rect 9680 20666 9732 20672
rect 5622 20420 5918 20440
rect 5678 20418 5702 20420
rect 5758 20418 5782 20420
rect 5838 20418 5862 20420
rect 5700 20366 5702 20418
rect 5764 20366 5776 20418
rect 5838 20366 5840 20418
rect 5678 20364 5702 20366
rect 5758 20364 5782 20366
rect 5838 20364 5862 20366
rect 5622 20344 5918 20364
rect 9692 20322 9720 20666
rect 9680 20316 9732 20322
rect 9680 20258 9732 20264
rect 5622 19332 5918 19352
rect 5678 19330 5702 19332
rect 5758 19330 5782 19332
rect 5838 19330 5862 19332
rect 5700 19278 5702 19330
rect 5764 19278 5776 19330
rect 5838 19278 5840 19330
rect 5678 19276 5702 19278
rect 5758 19276 5782 19278
rect 5838 19276 5862 19278
rect 5622 19256 5918 19276
rect 9876 19137 9904 23182
rect 10289 23140 10585 23160
rect 12072 23182 12124 23188
rect 10966 23143 11022 23152
rect 10345 23138 10369 23140
rect 10425 23138 10449 23140
rect 10505 23138 10529 23140
rect 10367 23086 10369 23138
rect 10431 23086 10443 23138
rect 10505 23086 10507 23138
rect 10345 23084 10369 23086
rect 10425 23084 10449 23086
rect 10505 23084 10529 23086
rect 10289 23064 10585 23084
rect 11336 22696 11388 22702
rect 11336 22638 11388 22644
rect 10876 22288 10928 22294
rect 10876 22230 10928 22236
rect 10289 22052 10585 22072
rect 10345 22050 10369 22052
rect 10425 22050 10449 22052
rect 10505 22050 10529 22052
rect 10367 21998 10369 22050
rect 10431 21998 10443 22050
rect 10505 21998 10507 22050
rect 10345 21996 10369 21998
rect 10425 21996 10449 21998
rect 10505 21996 10529 21998
rect 10289 21976 10585 21996
rect 10046 21848 10102 21857
rect 10046 21783 10102 21792
rect 10598 21848 10654 21857
rect 10598 21783 10654 21792
rect 10060 20186 10088 21783
rect 10508 21744 10560 21750
rect 10508 21686 10560 21692
rect 10520 21410 10548 21686
rect 10612 21614 10640 21783
rect 10600 21608 10652 21614
rect 10600 21550 10652 21556
rect 10692 21608 10744 21614
rect 10692 21550 10744 21556
rect 10508 21404 10560 21410
rect 10508 21346 10560 21352
rect 10612 21138 10640 21550
rect 10600 21132 10652 21138
rect 10600 21074 10652 21080
rect 10289 20964 10585 20984
rect 10345 20962 10369 20964
rect 10425 20962 10449 20964
rect 10505 20962 10529 20964
rect 10367 20910 10369 20962
rect 10431 20910 10443 20962
rect 10505 20910 10507 20962
rect 10345 20908 10369 20910
rect 10425 20908 10449 20910
rect 10505 20908 10529 20910
rect 10289 20888 10585 20908
rect 10704 20662 10732 21550
rect 10784 21200 10836 21206
rect 10888 21154 10916 22230
rect 11348 22226 11376 22638
rect 11336 22220 11388 22226
rect 11336 22162 11388 22168
rect 11152 21880 11204 21886
rect 11152 21822 11204 21828
rect 10836 21148 10916 21154
rect 10784 21142 10916 21148
rect 10796 21126 10916 21142
rect 10140 20656 10192 20662
rect 10140 20598 10192 20604
rect 10692 20656 10744 20662
rect 10692 20598 10744 20604
rect 10152 20254 10180 20598
rect 10140 20248 10192 20254
rect 10140 20190 10192 20196
rect 10048 20180 10100 20186
rect 10048 20122 10100 20128
rect 10888 20118 10916 21126
rect 11060 20792 11112 20798
rect 10980 20740 11060 20746
rect 10980 20734 11112 20740
rect 10980 20718 11100 20734
rect 10980 20186 11008 20718
rect 11164 20526 11192 21822
rect 11348 21750 11376 22162
rect 11336 21744 11388 21750
rect 11336 21686 11388 21692
rect 11348 21410 11376 21686
rect 11336 21404 11388 21410
rect 11336 21346 11388 21352
rect 11348 20866 11376 21346
rect 11336 20860 11388 20866
rect 11336 20802 11388 20808
rect 12084 20769 12112 23182
rect 12164 22152 12216 22158
rect 12164 22094 12216 22100
rect 12176 20798 12204 22094
rect 12360 21041 12388 23726
rect 12544 23382 12572 27240
rect 13188 24577 13216 27240
rect 13174 24568 13230 24577
rect 13174 24503 13230 24512
rect 12900 23988 12952 23994
rect 12900 23930 12952 23936
rect 12912 23586 12940 23930
rect 13728 23920 13780 23926
rect 13728 23862 13780 23868
rect 13740 23586 13768 23862
rect 12900 23580 12952 23586
rect 12900 23522 12952 23528
rect 13728 23580 13780 23586
rect 13728 23522 13780 23528
rect 12532 23376 12584 23382
rect 12532 23318 12584 23324
rect 12530 23072 12586 23081
rect 12530 23007 12586 23016
rect 12346 21032 12402 21041
rect 12346 20967 12402 20976
rect 12164 20792 12216 20798
rect 12070 20760 12126 20769
rect 12164 20734 12216 20740
rect 12070 20695 12126 20704
rect 12440 20724 12492 20730
rect 12440 20666 12492 20672
rect 12452 20594 12480 20666
rect 12440 20588 12492 20594
rect 12440 20530 12492 20536
rect 11152 20520 11204 20526
rect 11152 20462 11204 20468
rect 10968 20180 11020 20186
rect 10968 20122 11020 20128
rect 10876 20112 10928 20118
rect 10876 20054 10928 20060
rect 10289 19876 10585 19896
rect 10345 19874 10369 19876
rect 10425 19874 10449 19876
rect 10505 19874 10529 19876
rect 10367 19822 10369 19874
rect 10431 19822 10443 19874
rect 10505 19822 10507 19874
rect 10345 19820 10369 19822
rect 10425 19820 10449 19822
rect 10505 19820 10529 19822
rect 10289 19800 10585 19820
rect 11164 19817 11192 20462
rect 12452 20322 12480 20530
rect 12440 20316 12492 20322
rect 12440 20258 12492 20264
rect 11242 20216 11298 20225
rect 11242 20151 11298 20160
rect 11150 19808 11206 19817
rect 11256 19778 11284 20151
rect 12256 20112 12308 20118
rect 12256 20054 12308 20060
rect 11796 20044 11848 20050
rect 11796 19986 11848 19992
rect 11150 19743 11206 19752
rect 11244 19772 11296 19778
rect 11164 19710 11192 19743
rect 11244 19714 11296 19720
rect 11152 19704 11204 19710
rect 11152 19646 11204 19652
rect 11164 19522 11192 19646
rect 10980 19494 11192 19522
rect 9862 19128 9918 19137
rect 9862 19063 9918 19072
rect 4342 18992 4398 19001
rect 10980 18962 11008 19494
rect 11060 19432 11112 19438
rect 11060 19374 11112 19380
rect 11072 19030 11100 19374
rect 11256 19098 11284 19714
rect 11808 19438 11836 19986
rect 11796 19432 11848 19438
rect 11796 19374 11848 19380
rect 11244 19092 11296 19098
rect 11244 19034 11296 19040
rect 11060 19024 11112 19030
rect 11060 18966 11112 18972
rect 4342 18927 4398 18936
rect 10968 18956 11020 18962
rect 10968 18898 11020 18904
rect 11244 18956 11296 18962
rect 11244 18898 11296 18904
rect 11060 18888 11112 18894
rect 11060 18830 11112 18836
rect 10289 18788 10585 18808
rect 10345 18786 10369 18788
rect 10425 18786 10449 18788
rect 10505 18786 10529 18788
rect 10367 18734 10369 18786
rect 10431 18734 10443 18786
rect 10505 18734 10507 18786
rect 10345 18732 10369 18734
rect 10425 18732 10449 18734
rect 10505 18732 10529 18734
rect 10289 18712 10585 18732
rect 10876 18344 10928 18350
rect 10874 18312 10876 18321
rect 10928 18312 10930 18321
rect 5622 18244 5918 18264
rect 10874 18247 10930 18256
rect 5678 18242 5702 18244
rect 5758 18242 5782 18244
rect 5838 18242 5862 18244
rect 5700 18190 5702 18242
rect 5764 18190 5776 18242
rect 5838 18190 5840 18242
rect 5678 18188 5702 18190
rect 5758 18188 5782 18190
rect 5838 18188 5862 18190
rect 5622 18168 5918 18188
rect 2962 17904 3018 17913
rect 2962 17839 3018 17848
rect 10289 17700 10585 17720
rect 10345 17698 10369 17700
rect 10425 17698 10449 17700
rect 10505 17698 10529 17700
rect 10367 17646 10369 17698
rect 10431 17646 10443 17698
rect 10505 17646 10507 17698
rect 10345 17644 10369 17646
rect 10425 17644 10449 17646
rect 10505 17644 10529 17646
rect 10289 17624 10585 17644
rect 5622 17156 5918 17176
rect 5678 17154 5702 17156
rect 5758 17154 5782 17156
rect 5838 17154 5862 17156
rect 5700 17102 5702 17154
rect 5764 17102 5776 17154
rect 5838 17102 5840 17154
rect 5678 17100 5702 17102
rect 5758 17100 5782 17102
rect 5838 17100 5862 17102
rect 5622 17080 5918 17100
rect 10289 16612 10585 16632
rect 10345 16610 10369 16612
rect 10425 16610 10449 16612
rect 10505 16610 10529 16612
rect 10367 16558 10369 16610
rect 10431 16558 10443 16610
rect 10505 16558 10507 16610
rect 10345 16556 10369 16558
rect 10425 16556 10449 16558
rect 10505 16556 10529 16558
rect 10289 16536 10585 16556
rect 5622 16068 5918 16088
rect 5678 16066 5702 16068
rect 5758 16066 5782 16068
rect 5838 16066 5862 16068
rect 5700 16014 5702 16066
rect 5764 16014 5776 16066
rect 5838 16014 5840 16066
rect 5678 16012 5702 16014
rect 5758 16012 5782 16014
rect 5838 16012 5862 16014
rect 5622 15992 5918 16012
rect 11072 15766 11100 18830
rect 11256 18690 11284 18898
rect 11244 18684 11296 18690
rect 11244 18626 11296 18632
rect 11808 18321 11836 19374
rect 12268 19030 12296 20054
rect 12348 19568 12400 19574
rect 12348 19510 12400 19516
rect 12256 19024 12308 19030
rect 12256 18966 12308 18972
rect 11794 18312 11850 18321
rect 11794 18247 11850 18256
rect 12268 18146 12296 18966
rect 12360 18962 12388 19510
rect 12348 18956 12400 18962
rect 12348 18898 12400 18904
rect 12438 18312 12494 18321
rect 12438 18247 12494 18256
rect 12452 18146 12480 18247
rect 12256 18140 12308 18146
rect 12256 18082 12308 18088
rect 12440 18140 12492 18146
rect 12440 18082 12492 18088
rect 11152 17868 11204 17874
rect 11152 17810 11204 17816
rect 11164 17262 11192 17810
rect 11152 17256 11204 17262
rect 11152 17198 11204 17204
rect 11164 16990 11192 17198
rect 11152 16984 11204 16990
rect 11152 16926 11204 16932
rect 11060 15760 11112 15766
rect 11060 15702 11112 15708
rect 12256 15624 12308 15630
rect 12256 15566 12308 15572
rect 10289 15524 10585 15544
rect 10345 15522 10369 15524
rect 10425 15522 10449 15524
rect 10505 15522 10529 15524
rect 10367 15470 10369 15522
rect 10431 15470 10443 15522
rect 10505 15470 10507 15522
rect 10345 15468 10369 15470
rect 10425 15468 10449 15470
rect 10505 15468 10529 15470
rect 10289 15448 10585 15468
rect 5622 14980 5918 15000
rect 5678 14978 5702 14980
rect 5758 14978 5782 14980
rect 5838 14978 5862 14980
rect 5700 14926 5702 14978
rect 5764 14926 5776 14978
rect 5838 14926 5840 14978
rect 5678 14924 5702 14926
rect 5758 14924 5782 14926
rect 5838 14924 5862 14926
rect 5622 14904 5918 14924
rect 12268 14649 12296 15566
rect 12544 15426 12572 23007
rect 13636 22696 13688 22702
rect 13636 22638 13688 22644
rect 13820 22696 13872 22702
rect 13820 22638 13872 22644
rect 13544 22492 13596 22498
rect 13544 22434 13596 22440
rect 12622 20624 12678 20633
rect 12622 20559 12624 20568
rect 12676 20559 12678 20568
rect 12624 20530 12676 20536
rect 12808 19976 12860 19982
rect 12808 19918 12860 19924
rect 12820 19030 12848 19918
rect 12808 19024 12860 19030
rect 12808 18966 12860 18972
rect 12820 18690 12848 18966
rect 13556 18729 13584 22434
rect 13648 22294 13676 22638
rect 13832 22362 13860 22638
rect 13820 22356 13872 22362
rect 13820 22298 13872 22304
rect 13636 22288 13688 22294
rect 13636 22230 13688 22236
rect 13648 21954 13676 22230
rect 13728 22152 13780 22158
rect 13728 22094 13780 22100
rect 13636 21948 13688 21954
rect 13636 21890 13688 21896
rect 13648 21857 13676 21890
rect 13634 21848 13690 21857
rect 13634 21783 13690 21792
rect 13636 21744 13688 21750
rect 13636 21686 13688 21692
rect 13648 21410 13676 21686
rect 13636 21404 13688 21410
rect 13636 21346 13688 21352
rect 13740 19778 13768 22094
rect 13820 21404 13872 21410
rect 13820 21346 13872 21352
rect 13636 19772 13688 19778
rect 13636 19714 13688 19720
rect 13728 19772 13780 19778
rect 13728 19714 13780 19720
rect 13648 19681 13676 19714
rect 13634 19672 13690 19681
rect 13634 19607 13690 19616
rect 13832 19574 13860 21346
rect 13820 19568 13872 19574
rect 13820 19510 13872 19516
rect 13832 18962 13860 19510
rect 13820 18956 13872 18962
rect 13820 18898 13872 18904
rect 13542 18720 13598 18729
rect 12808 18684 12860 18690
rect 13542 18655 13598 18664
rect 12808 18626 12860 18632
rect 13556 17942 13584 18655
rect 13544 17936 13596 17942
rect 13450 17904 13506 17913
rect 13544 17878 13596 17884
rect 13450 17839 13452 17848
rect 13504 17839 13506 17848
rect 13452 17810 13504 17816
rect 13556 17602 13584 17878
rect 13636 17800 13688 17806
rect 13636 17742 13688 17748
rect 13544 17596 13596 17602
rect 13544 17538 13596 17544
rect 13648 16922 13676 17742
rect 13832 17466 13860 18898
rect 13924 18049 13952 27240
rect 14464 23784 14516 23790
rect 14464 23726 14516 23732
rect 14096 23376 14148 23382
rect 14096 23318 14148 23324
rect 14108 23081 14136 23318
rect 14280 23240 14332 23246
rect 14280 23182 14332 23188
rect 14292 23081 14320 23182
rect 14094 23072 14150 23081
rect 14094 23007 14150 23016
rect 14278 23072 14334 23081
rect 14278 23007 14334 23016
rect 14278 22936 14334 22945
rect 14188 22900 14240 22906
rect 14278 22871 14280 22880
rect 14188 22842 14240 22848
rect 14332 22871 14334 22880
rect 14280 22842 14332 22848
rect 14096 22832 14148 22838
rect 14096 22774 14148 22780
rect 14108 22158 14136 22774
rect 14200 22498 14228 22842
rect 14292 22498 14320 22842
rect 14476 22838 14504 23726
rect 14568 23586 14596 27240
rect 14956 24772 15252 24792
rect 15012 24770 15036 24772
rect 15092 24770 15116 24772
rect 15172 24770 15196 24772
rect 15034 24718 15036 24770
rect 15098 24718 15110 24770
rect 15172 24718 15174 24770
rect 15012 24716 15036 24718
rect 15092 24716 15116 24718
rect 15172 24716 15196 24718
rect 14956 24696 15252 24716
rect 15304 24538 15332 27240
rect 15292 24532 15344 24538
rect 15292 24474 15344 24480
rect 15108 23988 15160 23994
rect 15108 23930 15160 23936
rect 15120 23897 15148 23930
rect 15106 23888 15162 23897
rect 15106 23823 15162 23832
rect 14956 23684 15252 23704
rect 15012 23682 15036 23684
rect 15092 23682 15116 23684
rect 15172 23682 15196 23684
rect 15034 23630 15036 23682
rect 15098 23630 15110 23682
rect 15172 23630 15174 23682
rect 15012 23628 15036 23630
rect 15092 23628 15116 23630
rect 15172 23628 15196 23630
rect 14956 23608 15252 23628
rect 15948 23586 15976 27240
rect 16488 24532 16540 24538
rect 16488 24474 16540 24480
rect 14556 23580 14608 23586
rect 14556 23522 14608 23528
rect 15936 23580 15988 23586
rect 15936 23522 15988 23528
rect 16304 23580 16356 23586
rect 16304 23522 16356 23528
rect 15292 23376 15344 23382
rect 15292 23318 15344 23324
rect 14464 22832 14516 22838
rect 14464 22774 14516 22780
rect 14956 22596 15252 22616
rect 15012 22594 15036 22596
rect 15092 22594 15116 22596
rect 15172 22594 15196 22596
rect 15034 22542 15036 22594
rect 15098 22542 15110 22594
rect 15172 22542 15174 22594
rect 15012 22540 15036 22542
rect 15092 22540 15116 22542
rect 15172 22540 15196 22542
rect 14956 22520 15252 22540
rect 14188 22492 14240 22498
rect 14188 22434 14240 22440
rect 14280 22492 14332 22498
rect 14280 22434 14332 22440
rect 14188 22220 14240 22226
rect 14188 22162 14240 22168
rect 14096 22152 14148 22158
rect 14096 22094 14148 22100
rect 14108 21886 14136 22094
rect 14096 21880 14148 21886
rect 14096 21822 14148 21828
rect 14108 21410 14136 21822
rect 14096 21404 14148 21410
rect 14096 21346 14148 21352
rect 14108 20594 14136 21346
rect 14200 20866 14228 22162
rect 14956 21508 15252 21528
rect 15012 21506 15036 21508
rect 15092 21506 15116 21508
rect 15172 21506 15196 21508
rect 15034 21454 15036 21506
rect 15098 21454 15110 21506
rect 15172 21454 15174 21506
rect 15012 21452 15036 21454
rect 15092 21452 15116 21454
rect 15172 21452 15196 21454
rect 14956 21432 15252 21452
rect 14556 21064 14608 21070
rect 14556 21006 14608 21012
rect 14188 20860 14240 20866
rect 14188 20802 14240 20808
rect 14568 20730 14596 21006
rect 14556 20724 14608 20730
rect 14556 20666 14608 20672
rect 14096 20588 14148 20594
rect 14096 20530 14148 20536
rect 14108 20322 14136 20530
rect 14568 20322 14596 20666
rect 14648 20656 14700 20662
rect 14648 20598 14700 20604
rect 14096 20316 14148 20322
rect 14096 20258 14148 20264
rect 14556 20316 14608 20322
rect 14556 20258 14608 20264
rect 14660 20254 14688 20598
rect 14956 20420 15252 20440
rect 15012 20418 15036 20420
rect 15092 20418 15116 20420
rect 15172 20418 15196 20420
rect 15034 20366 15036 20418
rect 15098 20366 15110 20418
rect 15172 20366 15174 20418
rect 15012 20364 15036 20366
rect 15092 20364 15116 20366
rect 15172 20364 15196 20366
rect 14956 20344 15252 20364
rect 14648 20248 14700 20254
rect 14648 20190 14700 20196
rect 14464 20112 14516 20118
rect 14464 20054 14516 20060
rect 14188 19976 14240 19982
rect 14188 19918 14240 19924
rect 14096 19636 14148 19642
rect 14096 19578 14148 19584
rect 14108 18894 14136 19578
rect 14096 18888 14148 18894
rect 14096 18830 14148 18836
rect 14108 18622 14136 18830
rect 14200 18690 14228 19918
rect 14476 19574 14504 20054
rect 14464 19568 14516 19574
rect 14464 19510 14516 19516
rect 14476 19234 14504 19510
rect 14464 19228 14516 19234
rect 14464 19170 14516 19176
rect 14188 18684 14240 18690
rect 14188 18626 14240 18632
rect 14096 18616 14148 18622
rect 14096 18558 14148 18564
rect 14188 18344 14240 18350
rect 14188 18286 14240 18292
rect 13910 18040 13966 18049
rect 14200 18010 14228 18286
rect 13910 17975 13966 17984
rect 14188 18004 14240 18010
rect 14188 17946 14240 17952
rect 13820 17460 13872 17466
rect 13820 17402 13872 17408
rect 14200 17262 14228 17946
rect 14372 17460 14424 17466
rect 14372 17402 14424 17408
rect 14188 17256 14240 17262
rect 14188 17198 14240 17204
rect 13636 16916 13688 16922
rect 13636 16858 13688 16864
rect 13648 16514 13676 16858
rect 13820 16712 13872 16718
rect 13820 16654 13872 16660
rect 13636 16508 13688 16514
rect 13636 16450 13688 16456
rect 13832 15766 13860 16654
rect 14200 16446 14228 17198
rect 14384 16922 14412 17402
rect 14660 17058 14688 20190
rect 14956 19332 15252 19352
rect 15012 19330 15036 19332
rect 15092 19330 15116 19332
rect 15172 19330 15196 19332
rect 15034 19278 15036 19330
rect 15098 19278 15110 19330
rect 15172 19278 15174 19330
rect 15012 19276 15036 19278
rect 15092 19276 15116 19278
rect 15172 19276 15196 19278
rect 14956 19256 15252 19276
rect 15304 19137 15332 23318
rect 16132 22838 16160 22869
rect 16120 22832 16172 22838
rect 16118 22800 16120 22809
rect 16172 22800 16174 22809
rect 16118 22735 16174 22744
rect 16132 22430 16160 22735
rect 16120 22424 16172 22430
rect 16120 22366 16172 22372
rect 16316 22362 16344 23522
rect 16304 22356 16356 22362
rect 16304 22298 16356 22304
rect 16316 21954 16344 22298
rect 16304 21948 16356 21954
rect 16304 21890 16356 21896
rect 16316 21449 16344 21890
rect 16302 21440 16358 21449
rect 16302 21375 16358 21384
rect 16026 21304 16082 21313
rect 16026 21239 16082 21248
rect 16040 20662 16068 21239
rect 16028 20656 16080 20662
rect 16316 20610 16344 21375
rect 16028 20598 16080 20604
rect 16040 20322 16068 20598
rect 16224 20582 16344 20610
rect 16224 20526 16252 20582
rect 16212 20520 16264 20526
rect 16212 20462 16264 20468
rect 16028 20316 16080 20322
rect 16028 20258 16080 20264
rect 16224 20118 16252 20462
rect 16212 20112 16264 20118
rect 16212 20054 16264 20060
rect 15844 20044 15896 20050
rect 15844 19986 15896 19992
rect 15856 19778 15884 19986
rect 16394 19808 16450 19817
rect 15844 19772 15896 19778
rect 16394 19743 16396 19752
rect 15844 19714 15896 19720
rect 16448 19743 16450 19752
rect 16396 19714 16448 19720
rect 14738 19128 14794 19137
rect 14738 19063 14794 19072
rect 15290 19128 15346 19137
rect 15290 19063 15346 19072
rect 14648 17052 14700 17058
rect 14648 16994 14700 17000
rect 14280 16916 14332 16922
rect 14280 16858 14332 16864
rect 14372 16916 14424 16922
rect 14372 16858 14424 16864
rect 14292 16514 14320 16858
rect 14384 16530 14412 16858
rect 14280 16508 14332 16514
rect 14384 16502 14504 16530
rect 14280 16450 14332 16456
rect 14476 16446 14504 16502
rect 14188 16440 14240 16446
rect 14188 16382 14240 16388
rect 14464 16440 14516 16446
rect 14464 16382 14516 16388
rect 14200 15970 14228 16382
rect 14476 15970 14504 16382
rect 14188 15964 14240 15970
rect 14188 15906 14240 15912
rect 14464 15964 14516 15970
rect 14464 15906 14516 15912
rect 13820 15760 13872 15766
rect 13820 15702 13872 15708
rect 14372 15624 14424 15630
rect 14372 15566 14424 15572
rect 12532 15420 12584 15426
rect 12532 15362 12584 15368
rect 12440 15284 12492 15290
rect 12440 15226 12492 15232
rect 12452 14882 12480 15226
rect 13452 15080 13504 15086
rect 13452 15022 13504 15028
rect 12440 14876 12492 14882
rect 12440 14818 12492 14824
rect 13464 14746 13492 15022
rect 13452 14740 13504 14746
rect 13452 14682 13504 14688
rect 12254 14640 12310 14649
rect 12254 14575 12310 14584
rect 12716 14604 12768 14610
rect 12716 14546 12768 14552
rect 10289 14436 10585 14456
rect 10345 14434 10369 14436
rect 10425 14434 10449 14436
rect 10505 14434 10529 14436
rect 10367 14382 10369 14434
rect 10431 14382 10443 14434
rect 10505 14382 10507 14434
rect 10345 14380 10369 14382
rect 10425 14380 10449 14382
rect 10505 14380 10529 14382
rect 10289 14360 10585 14380
rect 12728 14338 12756 14546
rect 12900 14536 12952 14542
rect 12900 14478 12952 14484
rect 12716 14332 12768 14338
rect 12716 14274 12768 14280
rect 5622 13892 5918 13912
rect 5678 13890 5702 13892
rect 5758 13890 5782 13892
rect 5838 13890 5862 13892
rect 5700 13838 5702 13890
rect 5764 13838 5776 13890
rect 5838 13838 5840 13890
rect 5678 13836 5702 13838
rect 5758 13836 5782 13838
rect 5838 13836 5862 13838
rect 5622 13816 5918 13836
rect 12072 13788 12124 13794
rect 12072 13730 12124 13736
rect 1490 13688 1546 13697
rect 1490 13623 1546 13632
rect 386 13144 442 13153
rect 1504 13114 1532 13623
rect 12084 13590 12112 13730
rect 11704 13584 11756 13590
rect 2778 13552 2834 13561
rect 2778 13487 2834 13496
rect 11702 13552 11704 13561
rect 12072 13584 12124 13590
rect 11756 13552 11758 13561
rect 12072 13526 12124 13532
rect 11702 13487 11758 13496
rect 2792 13250 2820 13487
rect 10289 13348 10585 13368
rect 10345 13346 10369 13348
rect 10425 13346 10449 13348
rect 10505 13346 10529 13348
rect 10367 13294 10369 13346
rect 10431 13294 10443 13346
rect 10505 13294 10507 13346
rect 10345 13292 10369 13294
rect 10425 13292 10449 13294
rect 10505 13292 10529 13294
rect 10289 13272 10585 13292
rect 2780 13244 2832 13250
rect 2780 13186 2832 13192
rect 2044 13176 2096 13182
rect 2044 13118 2096 13124
rect 386 13079 442 13088
rect 1492 13108 1544 13114
rect 1492 13050 1544 13056
rect 1504 12706 1532 13050
rect 2056 13017 2084 13118
rect 12084 13017 12112 13526
rect 12912 13250 12940 14478
rect 13464 14270 13492 14682
rect 13452 14264 13504 14270
rect 13452 14206 13504 14212
rect 13360 14196 13412 14202
rect 13360 14138 13412 14144
rect 13372 13794 13400 14138
rect 13464 13794 13492 14206
rect 13360 13788 13412 13794
rect 13360 13730 13412 13736
rect 13452 13788 13504 13794
rect 13452 13730 13504 13736
rect 14384 13697 14412 15566
rect 14476 14202 14504 15906
rect 14752 15426 14780 19063
rect 15014 18992 15070 19001
rect 15014 18927 15016 18936
rect 15068 18927 15070 18936
rect 15016 18898 15068 18904
rect 15384 18888 15436 18894
rect 15384 18830 15436 18836
rect 14832 18684 14884 18690
rect 14832 18626 14884 18632
rect 14844 18146 14872 18626
rect 15396 18486 15424 18830
rect 15856 18486 15884 19714
rect 15936 19092 15988 19098
rect 15936 19034 15988 19040
rect 15948 18690 15976 19034
rect 16396 18888 16448 18894
rect 16396 18830 16448 18836
rect 15936 18684 15988 18690
rect 15936 18626 15988 18632
rect 15384 18480 15436 18486
rect 15384 18422 15436 18428
rect 15844 18480 15896 18486
rect 16408 18457 16436 18830
rect 15844 18422 15896 18428
rect 16394 18448 16450 18457
rect 15292 18344 15344 18350
rect 15292 18286 15344 18292
rect 14956 18244 15252 18264
rect 15012 18242 15036 18244
rect 15092 18242 15116 18244
rect 15172 18242 15196 18244
rect 15034 18190 15036 18242
rect 15098 18190 15110 18242
rect 15172 18190 15174 18242
rect 15012 18188 15036 18190
rect 15092 18188 15116 18190
rect 15172 18188 15196 18190
rect 14956 18168 15252 18188
rect 14832 18140 14884 18146
rect 14832 18082 14884 18088
rect 15304 17942 15332 18286
rect 15396 18146 15424 18422
rect 15384 18140 15436 18146
rect 15384 18082 15436 18088
rect 15856 18078 15884 18422
rect 16394 18383 16450 18392
rect 15844 18072 15896 18078
rect 15844 18014 15896 18020
rect 15292 17936 15344 17942
rect 15292 17878 15344 17884
rect 15476 17800 15528 17806
rect 15476 17742 15528 17748
rect 15108 17528 15160 17534
rect 15106 17496 15108 17505
rect 15160 17496 15162 17505
rect 15106 17431 15162 17440
rect 14956 17156 15252 17176
rect 15012 17154 15036 17156
rect 15092 17154 15116 17156
rect 15172 17154 15196 17156
rect 15034 17102 15036 17154
rect 15098 17102 15110 17154
rect 15172 17102 15174 17154
rect 15012 17100 15036 17102
rect 15092 17100 15116 17102
rect 15172 17100 15196 17102
rect 14956 17080 15252 17100
rect 15488 16961 15516 17742
rect 15844 17256 15896 17262
rect 15844 17198 15896 17204
rect 15474 16952 15530 16961
rect 15856 16922 15884 17198
rect 15474 16887 15530 16896
rect 15844 16916 15896 16922
rect 15844 16858 15896 16864
rect 15752 16848 15804 16854
rect 15750 16816 15752 16825
rect 15804 16816 15806 16825
rect 15660 16780 15712 16786
rect 15750 16751 15806 16760
rect 15660 16722 15712 16728
rect 14956 16068 15252 16088
rect 15012 16066 15036 16068
rect 15092 16066 15116 16068
rect 15172 16066 15196 16068
rect 15034 16014 15036 16066
rect 15098 16014 15110 16066
rect 15172 16014 15174 16066
rect 15012 16012 15036 16014
rect 15092 16012 15116 16014
rect 15172 16012 15196 16014
rect 14956 15992 15252 16012
rect 15672 15834 15700 16722
rect 15856 16514 15884 16858
rect 15844 16508 15896 16514
rect 15844 16450 15896 16456
rect 15660 15828 15712 15834
rect 15660 15770 15712 15776
rect 14740 15420 14792 15426
rect 14740 15362 14792 15368
rect 14648 15284 14700 15290
rect 14648 15226 14700 15232
rect 14660 14814 14688 15226
rect 15844 15080 15896 15086
rect 15844 15022 15896 15028
rect 14956 14980 15252 15000
rect 15012 14978 15036 14980
rect 15092 14978 15116 14980
rect 15172 14978 15196 14980
rect 15034 14926 15036 14978
rect 15098 14926 15110 14978
rect 15172 14926 15174 14978
rect 15012 14924 15036 14926
rect 15092 14924 15116 14926
rect 15172 14924 15196 14926
rect 14956 14904 15252 14924
rect 14648 14808 14700 14814
rect 14648 14750 14700 14756
rect 15856 14746 15884 15022
rect 15844 14740 15896 14746
rect 15844 14682 15896 14688
rect 15476 14536 15528 14542
rect 15476 14478 15528 14484
rect 14464 14196 14516 14202
rect 14464 14138 14516 14144
rect 14476 13726 14504 14138
rect 15384 13992 15436 13998
rect 15384 13934 15436 13940
rect 14956 13892 15252 13912
rect 15012 13890 15036 13892
rect 15092 13890 15116 13892
rect 15172 13890 15196 13892
rect 15034 13838 15036 13890
rect 15098 13838 15110 13890
rect 15172 13838 15174 13890
rect 15012 13836 15036 13838
rect 15092 13836 15116 13838
rect 15172 13836 15196 13838
rect 14956 13816 15252 13836
rect 14464 13720 14516 13726
rect 14370 13688 14426 13697
rect 14464 13662 14516 13668
rect 14370 13623 14426 13632
rect 15396 13590 15424 13934
rect 13636 13584 13688 13590
rect 13636 13526 13688 13532
rect 15384 13584 15436 13590
rect 15384 13526 15436 13532
rect 12900 13244 12952 13250
rect 12900 13186 12952 13192
rect 13358 13144 13414 13153
rect 13268 13108 13320 13114
rect 13358 13079 13414 13088
rect 13268 13050 13320 13056
rect 2042 13008 2098 13017
rect 2042 12943 2098 12952
rect 2870 13008 2926 13017
rect 2870 12943 2926 12952
rect 12070 13008 12126 13017
rect 12070 12943 12126 12952
rect 2056 12706 2084 12943
rect 1492 12700 1544 12706
rect 1492 12642 1544 12648
rect 2044 12700 2096 12706
rect 2044 12642 2096 12648
rect 2884 4449 2912 12943
rect 5622 12804 5918 12824
rect 5678 12802 5702 12804
rect 5758 12802 5782 12804
rect 5838 12802 5862 12804
rect 5700 12750 5702 12802
rect 5764 12750 5776 12802
rect 5838 12750 5840 12802
rect 5678 12748 5702 12750
rect 5758 12748 5782 12750
rect 5838 12748 5862 12750
rect 5622 12728 5918 12748
rect 13280 12706 13308 13050
rect 13372 13046 13400 13079
rect 13648 13046 13676 13526
rect 15396 13182 15424 13526
rect 15488 13250 15516 14478
rect 15856 13776 15884 14682
rect 16212 14604 16264 14610
rect 16212 14546 16264 14552
rect 16224 14338 16252 14546
rect 16212 14332 16264 14338
rect 16212 14274 16264 14280
rect 15936 13788 15988 13794
rect 15856 13748 15936 13776
rect 15936 13730 15988 13736
rect 15476 13244 15528 13250
rect 15476 13186 15528 13192
rect 15384 13176 15436 13182
rect 15384 13118 15436 13124
rect 15844 13108 15896 13114
rect 15844 13050 15896 13056
rect 13360 13040 13412 13046
rect 13360 12982 13412 12988
rect 13636 13040 13688 13046
rect 13636 12982 13688 12988
rect 13268 12700 13320 12706
rect 13268 12642 13320 12648
rect 10289 12260 10585 12280
rect 10345 12258 10369 12260
rect 10425 12258 10449 12260
rect 10505 12258 10529 12260
rect 10367 12206 10369 12258
rect 10431 12206 10443 12258
rect 10505 12206 10507 12258
rect 10345 12204 10369 12206
rect 10425 12204 10449 12206
rect 10505 12204 10529 12206
rect 10289 12184 10585 12204
rect 5622 11716 5918 11736
rect 5678 11714 5702 11716
rect 5758 11714 5782 11716
rect 5838 11714 5862 11716
rect 5700 11662 5702 11714
rect 5764 11662 5776 11714
rect 5838 11662 5840 11714
rect 5678 11660 5702 11662
rect 5758 11660 5782 11662
rect 5838 11660 5862 11662
rect 5622 11640 5918 11660
rect 10289 11172 10585 11192
rect 10345 11170 10369 11172
rect 10425 11170 10449 11172
rect 10505 11170 10529 11172
rect 10367 11118 10369 11170
rect 10431 11118 10443 11170
rect 10505 11118 10507 11170
rect 10345 11116 10369 11118
rect 10425 11116 10449 11118
rect 10505 11116 10529 11118
rect 10289 11096 10585 11116
rect 5622 10628 5918 10648
rect 5678 10626 5702 10628
rect 5758 10626 5782 10628
rect 5838 10626 5862 10628
rect 5700 10574 5702 10626
rect 5764 10574 5776 10626
rect 5838 10574 5840 10626
rect 5678 10572 5702 10574
rect 5758 10572 5782 10574
rect 5838 10572 5862 10574
rect 5622 10552 5918 10572
rect 10289 10084 10585 10104
rect 10345 10082 10369 10084
rect 10425 10082 10449 10084
rect 10505 10082 10529 10084
rect 10367 10030 10369 10082
rect 10431 10030 10443 10082
rect 10505 10030 10507 10082
rect 10345 10028 10369 10030
rect 10425 10028 10449 10030
rect 10505 10028 10529 10030
rect 10289 10008 10585 10028
rect 5622 9540 5918 9560
rect 5678 9538 5702 9540
rect 5758 9538 5782 9540
rect 5838 9538 5862 9540
rect 5700 9486 5702 9538
rect 5764 9486 5776 9538
rect 5838 9486 5840 9538
rect 5678 9484 5702 9486
rect 5758 9484 5782 9486
rect 5838 9484 5862 9486
rect 5622 9464 5918 9484
rect 10289 8996 10585 9016
rect 10345 8994 10369 8996
rect 10425 8994 10449 8996
rect 10505 8994 10529 8996
rect 10367 8942 10369 8994
rect 10431 8942 10443 8994
rect 10505 8942 10507 8994
rect 10345 8940 10369 8942
rect 10425 8940 10449 8942
rect 10505 8940 10529 8942
rect 10289 8920 10585 8940
rect 5622 8452 5918 8472
rect 5678 8450 5702 8452
rect 5758 8450 5782 8452
rect 5838 8450 5862 8452
rect 5700 8398 5702 8450
rect 5764 8398 5776 8450
rect 5838 8398 5840 8450
rect 5678 8396 5702 8398
rect 5758 8396 5782 8398
rect 5838 8396 5862 8398
rect 5622 8376 5918 8396
rect 10289 7908 10585 7928
rect 10345 7906 10369 7908
rect 10425 7906 10449 7908
rect 10505 7906 10529 7908
rect 10367 7854 10369 7906
rect 10431 7854 10443 7906
rect 10505 7854 10507 7906
rect 10345 7852 10369 7854
rect 10425 7852 10449 7854
rect 10505 7852 10529 7854
rect 10289 7832 10585 7852
rect 5622 7364 5918 7384
rect 5678 7362 5702 7364
rect 5758 7362 5782 7364
rect 5838 7362 5862 7364
rect 5700 7310 5702 7362
rect 5764 7310 5776 7362
rect 5838 7310 5840 7362
rect 5678 7308 5702 7310
rect 5758 7308 5782 7310
rect 5838 7308 5862 7310
rect 5622 7288 5918 7308
rect 10289 6820 10585 6840
rect 10345 6818 10369 6820
rect 10425 6818 10449 6820
rect 10505 6818 10529 6820
rect 10367 6766 10369 6818
rect 10431 6766 10443 6818
rect 10505 6766 10507 6818
rect 10345 6764 10369 6766
rect 10425 6764 10449 6766
rect 10505 6764 10529 6766
rect 10289 6744 10585 6764
rect 5622 6276 5918 6296
rect 5678 6274 5702 6276
rect 5758 6274 5782 6276
rect 5838 6274 5862 6276
rect 5700 6222 5702 6274
rect 5764 6222 5776 6274
rect 5838 6222 5840 6274
rect 5678 6220 5702 6222
rect 5758 6220 5782 6222
rect 5838 6220 5862 6222
rect 5622 6200 5918 6220
rect 10289 5732 10585 5752
rect 10345 5730 10369 5732
rect 10425 5730 10449 5732
rect 10505 5730 10529 5732
rect 10367 5678 10369 5730
rect 10431 5678 10443 5730
rect 10505 5678 10507 5730
rect 10345 5676 10369 5678
rect 10425 5676 10449 5678
rect 10505 5676 10529 5678
rect 10289 5656 10585 5676
rect 5622 5188 5918 5208
rect 5678 5186 5702 5188
rect 5758 5186 5782 5188
rect 5838 5186 5862 5188
rect 5700 5134 5702 5186
rect 5764 5134 5776 5186
rect 5838 5134 5840 5186
rect 5678 5132 5702 5134
rect 5758 5132 5782 5134
rect 5838 5132 5862 5134
rect 5622 5112 5918 5132
rect 10289 4644 10585 4664
rect 10345 4642 10369 4644
rect 10425 4642 10449 4644
rect 10505 4642 10529 4644
rect 10367 4590 10369 4642
rect 10431 4590 10443 4642
rect 10505 4590 10507 4642
rect 10345 4588 10369 4590
rect 10425 4588 10449 4590
rect 10505 4588 10529 4590
rect 10289 4568 10585 4588
rect 2870 4440 2926 4449
rect 2870 4375 2926 4384
rect 5622 4100 5918 4120
rect 5678 4098 5702 4100
rect 5758 4098 5782 4100
rect 5838 4098 5862 4100
rect 5700 4046 5702 4098
rect 5764 4046 5776 4098
rect 5838 4046 5840 4098
rect 5678 4044 5702 4046
rect 5758 4044 5782 4046
rect 5838 4044 5862 4046
rect 5622 4024 5918 4044
rect 10289 3556 10585 3576
rect 10345 3554 10369 3556
rect 10425 3554 10449 3556
rect 10505 3554 10529 3556
rect 10367 3502 10369 3554
rect 10431 3502 10443 3554
rect 10505 3502 10507 3554
rect 10345 3500 10369 3502
rect 10425 3500 10449 3502
rect 10505 3500 10529 3502
rect 10289 3480 10585 3500
rect 5622 3012 5918 3032
rect 5678 3010 5702 3012
rect 5758 3010 5782 3012
rect 5838 3010 5862 3012
rect 5700 2958 5702 3010
rect 5764 2958 5776 3010
rect 5838 2958 5840 3010
rect 5678 2956 5702 2958
rect 5758 2956 5782 2958
rect 5838 2956 5862 2958
rect 5622 2936 5918 2956
rect 10289 2468 10585 2488
rect 10345 2466 10369 2468
rect 10425 2466 10449 2468
rect 10505 2466 10529 2468
rect 10367 2414 10369 2466
rect 10431 2414 10443 2466
rect 10505 2414 10507 2466
rect 10345 2412 10369 2414
rect 10425 2412 10449 2414
rect 10505 2412 10529 2414
rect 10289 2392 10585 2412
rect 5622 1924 5918 1944
rect 5678 1922 5702 1924
rect 5758 1922 5782 1924
rect 5838 1922 5862 1924
rect 5700 1870 5702 1922
rect 5764 1870 5776 1922
rect 5838 1870 5840 1922
rect 5678 1868 5702 1870
rect 5758 1868 5782 1870
rect 5838 1868 5862 1870
rect 5622 1848 5918 1868
rect 13280 1185 13308 12642
rect 13372 12502 13400 12982
rect 13648 12706 13676 12982
rect 14956 12804 15252 12824
rect 15012 12802 15036 12804
rect 15092 12802 15116 12804
rect 15172 12802 15196 12804
rect 15034 12750 15036 12802
rect 15098 12750 15110 12802
rect 15172 12750 15174 12802
rect 15012 12748 15036 12750
rect 15092 12748 15116 12750
rect 15172 12748 15196 12750
rect 14956 12728 15252 12748
rect 15856 12706 15884 13050
rect 15936 13040 15988 13046
rect 15936 12982 15988 12988
rect 16212 13040 16264 13046
rect 16212 12982 16264 12988
rect 13636 12700 13688 12706
rect 13636 12642 13688 12648
rect 15844 12700 15896 12706
rect 15844 12642 15896 12648
rect 13360 12496 13412 12502
rect 13358 12464 13360 12473
rect 13412 12464 13414 12473
rect 13358 12399 13414 12408
rect 14956 11716 15252 11736
rect 15012 11714 15036 11716
rect 15092 11714 15116 11716
rect 15172 11714 15196 11716
rect 15034 11662 15036 11714
rect 15098 11662 15110 11714
rect 15172 11662 15174 11714
rect 15012 11660 15036 11662
rect 15092 11660 15116 11662
rect 15172 11660 15196 11662
rect 14956 11640 15252 11660
rect 14956 10628 15252 10648
rect 15012 10626 15036 10628
rect 15092 10626 15116 10628
rect 15172 10626 15196 10628
rect 15034 10574 15036 10626
rect 15098 10574 15110 10626
rect 15172 10574 15174 10626
rect 15012 10572 15036 10574
rect 15092 10572 15116 10574
rect 15172 10572 15196 10574
rect 14956 10552 15252 10572
rect 14956 9540 15252 9560
rect 15012 9538 15036 9540
rect 15092 9538 15116 9540
rect 15172 9538 15196 9540
rect 15034 9486 15036 9538
rect 15098 9486 15110 9538
rect 15172 9486 15174 9538
rect 15012 9484 15036 9486
rect 15092 9484 15116 9486
rect 15172 9484 15196 9486
rect 14956 9464 15252 9484
rect 14956 8452 15252 8472
rect 15012 8450 15036 8452
rect 15092 8450 15116 8452
rect 15172 8450 15196 8452
rect 15034 8398 15036 8450
rect 15098 8398 15110 8450
rect 15172 8398 15174 8450
rect 15012 8396 15036 8398
rect 15092 8396 15116 8398
rect 15172 8396 15196 8398
rect 14956 8376 15252 8396
rect 14956 7364 15252 7384
rect 15012 7362 15036 7364
rect 15092 7362 15116 7364
rect 15172 7362 15196 7364
rect 15034 7310 15036 7362
rect 15098 7310 15110 7362
rect 15172 7310 15174 7362
rect 15012 7308 15036 7310
rect 15092 7308 15116 7310
rect 15172 7308 15196 7310
rect 14956 7288 15252 7308
rect 14956 6276 15252 6296
rect 15012 6274 15036 6276
rect 15092 6274 15116 6276
rect 15172 6274 15196 6276
rect 15034 6222 15036 6274
rect 15098 6222 15110 6274
rect 15172 6222 15174 6274
rect 15012 6220 15036 6222
rect 15092 6220 15116 6222
rect 15172 6220 15196 6222
rect 14956 6200 15252 6220
rect 14956 5188 15252 5208
rect 15012 5186 15036 5188
rect 15092 5186 15116 5188
rect 15172 5186 15196 5188
rect 15034 5134 15036 5186
rect 15098 5134 15110 5186
rect 15172 5134 15174 5186
rect 15012 5132 15036 5134
rect 15092 5132 15116 5134
rect 15172 5132 15196 5134
rect 14956 5112 15252 5132
rect 14956 4100 15252 4120
rect 15012 4098 15036 4100
rect 15092 4098 15116 4100
rect 15172 4098 15196 4100
rect 15034 4046 15036 4098
rect 15098 4046 15110 4098
rect 15172 4046 15174 4098
rect 15012 4044 15036 4046
rect 15092 4044 15116 4046
rect 15172 4044 15196 4046
rect 14956 4024 15252 4044
rect 14956 3012 15252 3032
rect 15012 3010 15036 3012
rect 15092 3010 15116 3012
rect 15172 3010 15196 3012
rect 15034 2958 15036 3010
rect 15098 2958 15110 3010
rect 15172 2958 15174 3010
rect 15012 2956 15036 2958
rect 15092 2956 15116 2958
rect 15172 2956 15196 2958
rect 14956 2936 15252 2956
rect 14956 1924 15252 1944
rect 15012 1922 15036 1924
rect 15092 1922 15116 1924
rect 15172 1922 15196 1924
rect 15034 1870 15036 1922
rect 15098 1870 15110 1922
rect 15172 1870 15174 1922
rect 15012 1868 15036 1870
rect 15092 1868 15116 1870
rect 15172 1868 15196 1870
rect 14956 1848 15252 1868
rect 15856 1321 15884 12642
rect 15948 12502 15976 12982
rect 16224 12706 16252 12982
rect 16212 12700 16264 12706
rect 16212 12642 16264 12648
rect 15936 12496 15988 12502
rect 15934 12464 15936 12473
rect 15988 12464 15990 12473
rect 15934 12399 15990 12408
rect 16500 8694 16528 24474
rect 16488 8688 16540 8694
rect 16488 8630 16540 8636
rect 16592 2930 16620 27240
rect 17328 24130 17356 27240
rect 17972 24538 18000 27240
rect 18708 27138 18736 27240
rect 18708 27110 18828 27138
rect 17960 24532 18012 24538
rect 17960 24474 18012 24480
rect 17316 24124 17368 24130
rect 17316 24066 17368 24072
rect 17224 23988 17276 23994
rect 17224 23930 17276 23936
rect 17236 23790 17264 23930
rect 17866 23888 17922 23897
rect 17866 23823 17922 23832
rect 16764 23784 16816 23790
rect 16764 23726 16816 23732
rect 17224 23784 17276 23790
rect 17224 23726 17276 23732
rect 16776 23382 16804 23726
rect 16764 23376 16816 23382
rect 16764 23318 16816 23324
rect 16776 22770 16804 23318
rect 16764 22764 16816 22770
rect 16764 22706 16816 22712
rect 16856 22696 16908 22702
rect 16856 22638 16908 22644
rect 16868 22294 16896 22638
rect 16856 22288 16908 22294
rect 16854 22256 16856 22265
rect 16908 22256 16910 22265
rect 16854 22191 16910 22200
rect 16764 20724 16816 20730
rect 16764 20666 16816 20672
rect 16672 20520 16724 20526
rect 16672 20462 16724 20468
rect 16684 19030 16712 20462
rect 16776 19817 16804 20666
rect 16856 20520 16908 20526
rect 16856 20462 16908 20468
rect 16762 19808 16818 19817
rect 16868 19778 16896 20462
rect 16762 19743 16818 19752
rect 16856 19772 16908 19778
rect 16776 19409 16804 19743
rect 16856 19714 16908 19720
rect 16762 19400 16818 19409
rect 16762 19335 16818 19344
rect 16672 19024 16724 19030
rect 16672 18966 16724 18972
rect 16868 16854 16896 19714
rect 16948 17800 17000 17806
rect 16948 17742 17000 17748
rect 16960 16922 16988 17742
rect 16948 16916 17000 16922
rect 16948 16858 17000 16864
rect 16856 16848 16908 16854
rect 16856 16790 16908 16796
rect 16868 16514 16896 16790
rect 16960 16718 16988 16858
rect 16948 16712 17000 16718
rect 16948 16654 17000 16660
rect 16856 16508 16908 16514
rect 16856 16450 16908 16456
rect 16960 15970 16988 16654
rect 16948 15964 17000 15970
rect 16948 15906 17000 15912
rect 17132 15692 17184 15698
rect 17132 15634 17184 15640
rect 17144 15426 17172 15634
rect 17132 15420 17184 15426
rect 17132 15362 17184 15368
rect 17236 14882 17264 23726
rect 17880 23586 17908 23823
rect 17868 23580 17920 23586
rect 17868 23522 17920 23528
rect 17880 23194 17908 23522
rect 17880 23166 18000 23194
rect 17500 22900 17552 22906
rect 17500 22842 17552 22848
rect 17512 22498 17540 22842
rect 17972 22838 18000 23166
rect 18236 22900 18288 22906
rect 18236 22842 18288 22848
rect 17960 22832 18012 22838
rect 17960 22774 18012 22780
rect 17684 22764 17736 22770
rect 17684 22706 17736 22712
rect 17696 22498 17724 22706
rect 18052 22696 18104 22702
rect 18052 22638 18104 22644
rect 17500 22492 17552 22498
rect 17500 22434 17552 22440
rect 17684 22492 17736 22498
rect 17684 22434 17736 22440
rect 17316 19432 17368 19438
rect 17316 19374 17368 19380
rect 17328 19098 17356 19374
rect 17316 19092 17368 19098
rect 17316 19034 17368 19040
rect 17328 18894 17356 19034
rect 17512 18962 17540 22434
rect 17696 21886 17724 22434
rect 17684 21880 17736 21886
rect 17684 21822 17736 21828
rect 18064 21818 18092 22638
rect 18248 22158 18276 22842
rect 18604 22832 18656 22838
rect 18604 22774 18656 22780
rect 18616 22498 18644 22774
rect 18604 22492 18656 22498
rect 18604 22434 18656 22440
rect 18510 22392 18566 22401
rect 18510 22327 18566 22336
rect 18236 22152 18288 22158
rect 18236 22094 18288 22100
rect 18248 21954 18276 22094
rect 18236 21948 18288 21954
rect 18236 21890 18288 21896
rect 18234 21848 18290 21857
rect 18052 21812 18104 21818
rect 18234 21783 18290 21792
rect 18052 21754 18104 21760
rect 18064 21410 18092 21754
rect 18248 21682 18276 21783
rect 18236 21676 18288 21682
rect 18236 21618 18288 21624
rect 18142 21440 18198 21449
rect 18052 21404 18104 21410
rect 18142 21375 18144 21384
rect 18052 21346 18104 21352
rect 18196 21375 18198 21384
rect 18144 21346 18196 21352
rect 17776 21064 17828 21070
rect 17776 21006 17828 21012
rect 17788 20662 17816 21006
rect 18524 20866 18552 22327
rect 18512 20860 18564 20866
rect 18512 20802 18564 20808
rect 18420 20724 18472 20730
rect 18420 20666 18472 20672
rect 17776 20656 17828 20662
rect 17776 20598 17828 20604
rect 17788 19982 17816 20598
rect 18432 20186 18460 20666
rect 18524 20322 18552 20802
rect 18512 20316 18564 20322
rect 18512 20258 18564 20264
rect 18420 20180 18472 20186
rect 18420 20122 18472 20128
rect 17776 19976 17828 19982
rect 17776 19918 17828 19924
rect 18696 19976 18748 19982
rect 18696 19918 18748 19924
rect 17788 19778 17816 19918
rect 18708 19778 18736 19918
rect 17776 19772 17828 19778
rect 17776 19714 17828 19720
rect 18696 19772 18748 19778
rect 18696 19714 18748 19720
rect 17960 19568 18012 19574
rect 17880 19528 17960 19556
rect 17880 19030 17908 19528
rect 17960 19510 18012 19516
rect 18052 19432 18104 19438
rect 18052 19374 18104 19380
rect 17868 19024 17920 19030
rect 17868 18966 17920 18972
rect 17500 18956 17552 18962
rect 17500 18898 17552 18904
rect 17316 18888 17368 18894
rect 17316 18830 17368 18836
rect 17592 18888 17644 18894
rect 17592 18830 17644 18836
rect 17684 18888 17736 18894
rect 17684 18830 17736 18836
rect 17328 17874 17356 18830
rect 17604 18622 17632 18830
rect 17696 18690 17724 18830
rect 18064 18690 18092 19374
rect 18800 19035 18828 27110
rect 18880 24532 18932 24538
rect 18880 24474 18932 24480
rect 18786 19026 18842 19035
rect 18326 18992 18382 19001
rect 18786 18961 18842 18970
rect 18326 18927 18382 18936
rect 18144 18888 18196 18894
rect 18144 18830 18196 18836
rect 17684 18684 17736 18690
rect 17684 18626 17736 18632
rect 18052 18684 18104 18690
rect 18052 18626 18104 18632
rect 17592 18616 17644 18622
rect 17592 18558 17644 18564
rect 18052 18344 18104 18350
rect 18156 18321 18184 18830
rect 18236 18480 18288 18486
rect 18236 18422 18288 18428
rect 18052 18286 18104 18292
rect 18142 18312 18198 18321
rect 17316 17868 17368 17874
rect 17316 17810 17368 17816
rect 17328 17262 17356 17810
rect 17316 17256 17368 17262
rect 17316 17198 17368 17204
rect 17328 17058 17356 17198
rect 17316 17052 17368 17058
rect 17316 16994 17368 17000
rect 17960 16508 18012 16514
rect 17960 16450 18012 16456
rect 17972 15970 18000 16450
rect 17960 15964 18012 15970
rect 17960 15906 18012 15912
rect 17684 15760 17736 15766
rect 17684 15702 17736 15708
rect 17224 14876 17276 14882
rect 17224 14818 17276 14824
rect 17592 14536 17644 14542
rect 17592 14478 17644 14484
rect 17604 14338 17632 14478
rect 17592 14332 17644 14338
rect 17592 14274 17644 14280
rect 17696 13726 17724 15702
rect 18064 14678 18092 18286
rect 18142 18247 18198 18256
rect 18248 17806 18276 18422
rect 18236 17800 18288 17806
rect 18236 17742 18288 17748
rect 18248 17534 18276 17742
rect 18236 17528 18288 17534
rect 18234 17496 18236 17505
rect 18288 17496 18290 17505
rect 18234 17431 18290 17440
rect 18052 14672 18104 14678
rect 18052 14614 18104 14620
rect 18236 14536 18288 14542
rect 18236 14478 18288 14484
rect 18052 14196 18104 14202
rect 18052 14138 18104 14144
rect 18064 13794 18092 14138
rect 18052 13788 18104 13794
rect 18052 13730 18104 13736
rect 17684 13720 17736 13726
rect 17684 13662 17736 13668
rect 17696 13590 17724 13662
rect 17684 13584 17736 13590
rect 17684 13526 17736 13532
rect 17868 13584 17920 13590
rect 17868 13526 17920 13532
rect 17880 13250 17908 13526
rect 18064 13250 18092 13730
rect 17868 13244 17920 13250
rect 17868 13186 17920 13192
rect 18052 13244 18104 13250
rect 18052 13186 18104 13192
rect 18248 13017 18276 14478
rect 18234 13008 18290 13017
rect 18234 12943 18290 12952
rect 18340 12858 18368 18927
rect 18604 18616 18656 18622
rect 18604 18558 18656 18564
rect 18616 17602 18644 18558
rect 18604 17596 18656 17602
rect 18604 17538 18656 17544
rect 18512 14128 18564 14134
rect 18512 14070 18564 14076
rect 18604 14128 18656 14134
rect 18604 14070 18656 14076
rect 18524 13250 18552 14070
rect 18512 13244 18564 13250
rect 18512 13186 18564 13192
rect 18616 13182 18644 14070
rect 18696 13244 18748 13250
rect 18696 13186 18748 13192
rect 18604 13176 18656 13182
rect 18604 13118 18656 13124
rect 18248 12830 18368 12858
rect 18052 12700 18104 12706
rect 18052 12642 18104 12648
rect 18064 12502 18092 12642
rect 18052 12496 18104 12502
rect 18052 12438 18104 12444
rect 18248 9442 18276 12830
rect 18510 12464 18566 12473
rect 18510 12399 18566 12408
rect 18328 12020 18380 12026
rect 18328 11962 18380 11968
rect 18340 11278 18368 11962
rect 18524 11958 18552 12399
rect 18708 12162 18736 13186
rect 18892 12337 18920 24474
rect 19352 24062 19380 27240
rect 19984 26300 20036 26306
rect 19984 26242 20036 26248
rect 19622 25316 19918 25336
rect 19678 25314 19702 25316
rect 19758 25314 19782 25316
rect 19838 25314 19862 25316
rect 19700 25262 19702 25314
rect 19764 25262 19776 25314
rect 19838 25262 19840 25314
rect 19678 25260 19702 25262
rect 19758 25260 19782 25262
rect 19838 25260 19862 25262
rect 19622 25240 19918 25260
rect 19622 24228 19918 24248
rect 19678 24226 19702 24228
rect 19758 24226 19782 24228
rect 19838 24226 19862 24228
rect 19700 24174 19702 24226
rect 19764 24174 19776 24226
rect 19838 24174 19840 24226
rect 19678 24172 19702 24174
rect 19758 24172 19782 24174
rect 19838 24172 19862 24174
rect 19622 24152 19918 24172
rect 19340 24056 19392 24062
rect 19340 23998 19392 24004
rect 19892 23988 19944 23994
rect 19892 23930 19944 23936
rect 19616 23920 19668 23926
rect 19904 23897 19932 23930
rect 19890 23888 19946 23897
rect 19616 23862 19668 23868
rect 19628 23518 19656 23862
rect 19812 23846 19890 23874
rect 19812 23586 19840 23846
rect 19890 23823 19946 23832
rect 19892 23784 19944 23790
rect 19892 23726 19944 23732
rect 19800 23580 19852 23586
rect 19800 23522 19852 23528
rect 19616 23512 19668 23518
rect 19616 23454 19668 23460
rect 19904 23450 19932 23726
rect 19892 23444 19944 23450
rect 19892 23386 19944 23392
rect 19432 23376 19484 23382
rect 19062 23344 19118 23353
rect 19432 23318 19484 23324
rect 19062 23279 19064 23288
rect 19116 23279 19118 23288
rect 19064 23250 19116 23256
rect 19340 23240 19392 23246
rect 19340 23182 19392 23188
rect 18972 23036 19024 23042
rect 18972 22978 19024 22984
rect 18984 22498 19012 22978
rect 18972 22492 19024 22498
rect 18972 22434 19024 22440
rect 19352 21750 19380 23182
rect 19444 23042 19472 23318
rect 19904 23228 19932 23386
rect 19996 23382 20024 26242
rect 19984 23376 20036 23382
rect 19984 23318 20036 23324
rect 19904 23200 20024 23228
rect 19622 23140 19918 23160
rect 19678 23138 19702 23140
rect 19758 23138 19782 23140
rect 19838 23138 19862 23140
rect 19700 23086 19702 23138
rect 19764 23086 19776 23138
rect 19838 23086 19840 23138
rect 19678 23084 19702 23086
rect 19758 23084 19782 23086
rect 19838 23084 19862 23086
rect 19622 23064 19918 23084
rect 19432 23036 19484 23042
rect 19432 22978 19484 22984
rect 19996 22974 20024 23200
rect 19984 22968 20036 22974
rect 19984 22910 20036 22916
rect 19708 22900 19760 22906
rect 19708 22842 19760 22848
rect 19720 22498 19748 22842
rect 19996 22498 20024 22910
rect 19432 22492 19484 22498
rect 19432 22434 19484 22440
rect 19708 22492 19760 22498
rect 19708 22434 19760 22440
rect 19984 22492 20036 22498
rect 19984 22434 20036 22440
rect 19340 21744 19392 21750
rect 19340 21686 19392 21692
rect 19444 21449 19472 22434
rect 19622 22052 19918 22072
rect 19678 22050 19702 22052
rect 19758 22050 19782 22052
rect 19838 22050 19862 22052
rect 19700 21998 19702 22050
rect 19764 21998 19776 22050
rect 19838 21998 19840 22050
rect 19678 21996 19702 21998
rect 19758 21996 19782 21998
rect 19838 21996 19862 21998
rect 19622 21976 19918 21996
rect 19524 21744 19576 21750
rect 19524 21686 19576 21692
rect 19430 21440 19486 21449
rect 19430 21375 19486 21384
rect 19248 20520 19300 20526
rect 19248 20462 19300 20468
rect 19062 20216 19118 20225
rect 19260 20186 19288 20462
rect 19062 20151 19118 20160
rect 19248 20180 19300 20186
rect 19076 20118 19104 20151
rect 19248 20122 19300 20128
rect 19064 20112 19116 20118
rect 19064 20054 19116 20060
rect 19076 19710 19104 20054
rect 19064 19704 19116 19710
rect 19064 19646 19116 19652
rect 19444 19114 19472 21375
rect 19536 20866 19564 21686
rect 19622 20964 19918 20984
rect 19678 20962 19702 20964
rect 19758 20962 19782 20964
rect 19838 20962 19862 20964
rect 19700 20910 19702 20962
rect 19764 20910 19776 20962
rect 19838 20910 19840 20962
rect 19678 20908 19702 20910
rect 19758 20908 19782 20910
rect 19838 20908 19862 20910
rect 19622 20888 19918 20908
rect 19524 20860 19576 20866
rect 19524 20802 19576 20808
rect 19984 20724 20036 20730
rect 19984 20666 20036 20672
rect 19798 20352 19854 20361
rect 19996 20322 20024 20666
rect 19798 20287 19800 20296
rect 19852 20287 19854 20296
rect 19984 20316 20036 20322
rect 19800 20258 19852 20264
rect 19984 20258 20036 20264
rect 19622 19876 19918 19896
rect 19678 19874 19702 19876
rect 19758 19874 19782 19876
rect 19838 19874 19862 19876
rect 19700 19822 19702 19874
rect 19764 19822 19776 19874
rect 19838 19822 19840 19874
rect 19678 19820 19702 19822
rect 19758 19820 19782 19822
rect 19838 19820 19862 19822
rect 19622 19800 19918 19820
rect 19996 19778 20024 20258
rect 19984 19772 20036 19778
rect 19984 19714 20036 19720
rect 19444 19086 19840 19114
rect 19524 19024 19576 19030
rect 19524 18966 19576 18972
rect 18972 18888 19024 18894
rect 18972 18830 19024 18836
rect 19248 18888 19300 18894
rect 19248 18830 19300 18836
rect 19340 18888 19392 18894
rect 19340 18830 19392 18836
rect 18984 18593 19012 18830
rect 19064 18684 19116 18690
rect 19064 18626 19116 18632
rect 18970 18584 19026 18593
rect 18970 18519 19026 18528
rect 19076 18146 19104 18626
rect 19064 18140 19116 18146
rect 19064 18082 19116 18088
rect 19260 17913 19288 18830
rect 19352 18729 19380 18830
rect 19338 18720 19394 18729
rect 19338 18655 19340 18664
rect 19392 18655 19394 18664
rect 19340 18626 19392 18632
rect 19536 18418 19564 18966
rect 19812 18962 19840 19086
rect 19800 18956 19852 18962
rect 19800 18898 19852 18904
rect 19622 18788 19918 18808
rect 19678 18786 19702 18788
rect 19758 18786 19782 18788
rect 19838 18786 19862 18788
rect 19700 18734 19702 18786
rect 19764 18734 19776 18786
rect 19838 18734 19840 18786
rect 19678 18732 19702 18734
rect 19758 18732 19782 18734
rect 19838 18732 19862 18734
rect 19622 18712 19918 18732
rect 19524 18412 19576 18418
rect 19524 18354 19576 18360
rect 20088 18298 20116 27240
rect 20732 24470 20760 27240
rect 21376 24554 21404 27240
rect 21192 24526 21404 24554
rect 21732 24600 21784 24606
rect 21732 24542 21784 24548
rect 20720 24464 20772 24470
rect 20720 24406 20772 24412
rect 20444 24056 20496 24062
rect 20444 23998 20496 24004
rect 20168 23512 20220 23518
rect 20168 23454 20220 23460
rect 20180 22906 20208 23454
rect 20352 23376 20404 23382
rect 20352 23318 20404 23324
rect 20168 22900 20220 22906
rect 20168 22842 20220 22848
rect 20168 22152 20220 22158
rect 20168 22094 20220 22100
rect 20180 21954 20208 22094
rect 20168 21948 20220 21954
rect 20168 21890 20220 21896
rect 20180 21410 20208 21890
rect 20168 21404 20220 21410
rect 20168 21346 20220 21352
rect 20168 21064 20220 21070
rect 20168 21006 20220 21012
rect 20180 20662 20208 21006
rect 20168 20656 20220 20662
rect 20168 20598 20220 20604
rect 20180 20322 20208 20598
rect 20260 20588 20312 20594
rect 20260 20530 20312 20536
rect 20168 20316 20220 20322
rect 20168 20258 20220 20264
rect 20272 19778 20300 20530
rect 20260 19772 20312 19778
rect 20260 19714 20312 19720
rect 20168 18888 20220 18894
rect 20166 18856 20168 18865
rect 20220 18856 20222 18865
rect 20166 18791 20222 18800
rect 20168 18412 20220 18418
rect 20168 18354 20220 18360
rect 19996 18270 20116 18298
rect 19246 17904 19302 17913
rect 19246 17839 19302 17848
rect 19622 17700 19918 17720
rect 19678 17698 19702 17700
rect 19758 17698 19782 17700
rect 19838 17698 19862 17700
rect 19700 17646 19702 17698
rect 19764 17646 19776 17698
rect 19838 17646 19840 17698
rect 19678 17644 19702 17646
rect 19758 17644 19782 17646
rect 19838 17644 19862 17646
rect 19622 17624 19918 17644
rect 19156 17392 19208 17398
rect 19156 17334 19208 17340
rect 19168 17058 19196 17334
rect 19156 17052 19208 17058
rect 19156 16994 19208 17000
rect 19432 16712 19484 16718
rect 19432 16654 19484 16660
rect 19444 16514 19472 16654
rect 19622 16612 19918 16632
rect 19678 16610 19702 16612
rect 19758 16610 19782 16612
rect 19838 16610 19862 16612
rect 19700 16558 19702 16610
rect 19764 16558 19776 16610
rect 19838 16558 19840 16610
rect 19678 16556 19702 16558
rect 19758 16556 19782 16558
rect 19838 16556 19862 16558
rect 19622 16536 19918 16556
rect 19432 16508 19484 16514
rect 19432 16450 19484 16456
rect 19156 15760 19208 15766
rect 19156 15702 19208 15708
rect 19168 15290 19196 15702
rect 19444 15290 19472 16450
rect 19616 16304 19668 16310
rect 19616 16246 19668 16252
rect 19628 15766 19656 16246
rect 19616 15760 19668 15766
rect 19616 15702 19668 15708
rect 19622 15524 19918 15544
rect 19678 15522 19702 15524
rect 19758 15522 19782 15524
rect 19838 15522 19862 15524
rect 19700 15470 19702 15522
rect 19764 15470 19776 15522
rect 19838 15470 19840 15522
rect 19678 15468 19702 15470
rect 19758 15468 19782 15470
rect 19838 15468 19862 15470
rect 19622 15448 19918 15468
rect 19156 15284 19208 15290
rect 19156 15226 19208 15232
rect 19432 15284 19484 15290
rect 19432 15226 19484 15232
rect 19168 14882 19196 15226
rect 19444 14882 19472 15226
rect 19156 14876 19208 14882
rect 19156 14818 19208 14824
rect 19432 14876 19484 14882
rect 19432 14818 19484 14824
rect 19168 13572 19196 14818
rect 19622 14436 19918 14456
rect 19678 14434 19702 14436
rect 19758 14434 19782 14436
rect 19838 14434 19862 14436
rect 19700 14382 19702 14434
rect 19764 14382 19776 14434
rect 19838 14382 19840 14434
rect 19678 14380 19702 14382
rect 19758 14380 19782 14382
rect 19838 14380 19862 14382
rect 19622 14360 19918 14380
rect 19168 13544 19288 13572
rect 19156 13448 19208 13454
rect 19156 13390 19208 13396
rect 19168 12502 19196 13390
rect 19260 13046 19288 13544
rect 19622 13348 19918 13368
rect 19678 13346 19702 13348
rect 19758 13346 19782 13348
rect 19838 13346 19862 13348
rect 19700 13294 19702 13346
rect 19764 13294 19776 13346
rect 19838 13294 19840 13346
rect 19678 13292 19702 13294
rect 19758 13292 19782 13294
rect 19838 13292 19862 13294
rect 19622 13272 19918 13292
rect 19432 13176 19484 13182
rect 19432 13118 19484 13124
rect 19248 13040 19300 13046
rect 19248 12982 19300 12988
rect 19260 12706 19288 12982
rect 19444 12706 19472 13118
rect 19248 12700 19300 12706
rect 19248 12642 19300 12648
rect 19432 12700 19484 12706
rect 19432 12642 19484 12648
rect 19156 12496 19208 12502
rect 19156 12438 19208 12444
rect 18878 12328 18934 12337
rect 18878 12263 18934 12272
rect 18696 12156 18748 12162
rect 18696 12098 18748 12104
rect 18878 12056 18934 12065
rect 18878 11991 18934 12000
rect 18512 11952 18564 11958
rect 18512 11894 18564 11900
rect 18524 11618 18552 11894
rect 18512 11612 18564 11618
rect 18512 11554 18564 11560
rect 18328 11272 18380 11278
rect 18328 11214 18380 11220
rect 18236 9436 18288 9442
rect 18236 9378 18288 9384
rect 16672 8688 16724 8694
rect 16672 8630 16724 8636
rect 16500 2914 16620 2930
rect 16488 2908 16620 2914
rect 16540 2902 16620 2908
rect 16488 2850 16540 2856
rect 16684 2137 16712 8630
rect 18340 5401 18368 11214
rect 18326 5392 18382 5401
rect 18326 5327 18382 5336
rect 18892 3769 18920 11991
rect 19168 11958 19196 12438
rect 19444 12162 19472 12642
rect 19622 12260 19918 12280
rect 19678 12258 19702 12260
rect 19758 12258 19782 12260
rect 19838 12258 19862 12260
rect 19700 12206 19702 12258
rect 19764 12206 19776 12258
rect 19838 12206 19840 12258
rect 19678 12204 19702 12206
rect 19758 12204 19782 12206
rect 19838 12204 19862 12206
rect 19622 12184 19918 12204
rect 19432 12156 19484 12162
rect 19432 12098 19484 12104
rect 19156 11952 19208 11958
rect 19156 11894 19208 11900
rect 19168 11618 19196 11894
rect 19156 11612 19208 11618
rect 19156 11554 19208 11560
rect 19622 11172 19918 11192
rect 19678 11170 19702 11172
rect 19758 11170 19782 11172
rect 19838 11170 19862 11172
rect 19700 11118 19702 11170
rect 19764 11118 19776 11170
rect 19838 11118 19840 11170
rect 19678 11116 19702 11118
rect 19758 11116 19782 11118
rect 19838 11116 19862 11118
rect 19622 11096 19918 11116
rect 19622 10084 19918 10104
rect 19678 10082 19702 10084
rect 19758 10082 19782 10084
rect 19838 10082 19862 10084
rect 19700 10030 19702 10082
rect 19764 10030 19776 10082
rect 19838 10030 19840 10082
rect 19678 10028 19702 10030
rect 19758 10028 19782 10030
rect 19838 10028 19862 10030
rect 19622 10008 19918 10028
rect 18972 9436 19024 9442
rect 18972 9378 19024 9384
rect 18984 9322 19012 9378
rect 18984 9294 19104 9322
rect 19076 4857 19104 9294
rect 19622 8996 19918 9016
rect 19678 8994 19702 8996
rect 19758 8994 19782 8996
rect 19838 8994 19862 8996
rect 19700 8942 19702 8994
rect 19764 8942 19776 8994
rect 19838 8942 19840 8994
rect 19678 8940 19702 8942
rect 19758 8940 19782 8942
rect 19838 8940 19862 8942
rect 19622 8920 19918 8940
rect 19622 7908 19918 7928
rect 19678 7906 19702 7908
rect 19758 7906 19782 7908
rect 19838 7906 19862 7908
rect 19700 7854 19702 7906
rect 19764 7854 19776 7906
rect 19838 7854 19840 7906
rect 19678 7852 19702 7854
rect 19758 7852 19782 7854
rect 19838 7852 19862 7854
rect 19622 7832 19918 7852
rect 19622 6820 19918 6840
rect 19678 6818 19702 6820
rect 19758 6818 19782 6820
rect 19838 6818 19862 6820
rect 19700 6766 19702 6818
rect 19764 6766 19776 6818
rect 19838 6766 19840 6818
rect 19678 6764 19702 6766
rect 19758 6764 19782 6766
rect 19838 6764 19862 6766
rect 19622 6744 19918 6764
rect 19996 6178 20024 18270
rect 20180 18146 20208 18354
rect 20168 18140 20220 18146
rect 20088 18100 20168 18128
rect 20088 16922 20116 18100
rect 20168 18082 20220 18088
rect 20364 17534 20392 23318
rect 20352 17528 20404 17534
rect 20352 17470 20404 17476
rect 20168 17460 20220 17466
rect 20168 17402 20220 17408
rect 20180 17058 20208 17402
rect 20260 17392 20312 17398
rect 20260 17334 20312 17340
rect 20352 17392 20404 17398
rect 20352 17334 20404 17340
rect 20272 17058 20300 17334
rect 20168 17052 20220 17058
rect 20168 16994 20220 17000
rect 20260 17052 20312 17058
rect 20260 16994 20312 17000
rect 20076 16916 20128 16922
rect 20076 16858 20128 16864
rect 20088 16446 20116 16858
rect 20076 16440 20128 16446
rect 20076 16382 20128 16388
rect 20088 15970 20116 16382
rect 20076 15964 20128 15970
rect 20076 15906 20128 15912
rect 20180 15834 20208 16994
rect 20364 16514 20392 17334
rect 20352 16508 20404 16514
rect 20352 16450 20404 16456
rect 20168 15828 20220 15834
rect 20168 15770 20220 15776
rect 20352 6580 20404 6586
rect 20352 6522 20404 6528
rect 20364 6489 20392 6522
rect 20350 6480 20406 6489
rect 20350 6415 20406 6424
rect 20364 6178 20392 6415
rect 19984 6172 20036 6178
rect 19984 6114 20036 6120
rect 20352 6172 20404 6178
rect 20352 6114 20404 6120
rect 20076 5832 20128 5838
rect 20074 5800 20076 5809
rect 20128 5800 20130 5809
rect 19622 5732 19918 5752
rect 20074 5735 20130 5744
rect 19678 5730 19702 5732
rect 19758 5730 19782 5732
rect 19838 5730 19862 5732
rect 19700 5678 19702 5730
rect 19764 5678 19776 5730
rect 19838 5678 19840 5730
rect 19678 5676 19702 5678
rect 19758 5676 19782 5678
rect 19838 5676 19862 5678
rect 19622 5656 19918 5676
rect 20456 5129 20484 23998
rect 20536 22696 20588 22702
rect 20536 22638 20588 22644
rect 20548 22265 20576 22638
rect 20628 22288 20680 22294
rect 20534 22256 20590 22265
rect 20628 22230 20680 22236
rect 20534 22191 20590 22200
rect 20548 21750 20576 22191
rect 20536 21744 20588 21750
rect 20536 21686 20588 21692
rect 20640 21682 20668 22230
rect 20628 21676 20680 21682
rect 20628 21618 20680 21624
rect 20718 21440 20774 21449
rect 20718 21375 20720 21384
rect 20772 21375 20774 21384
rect 20720 21346 20772 21352
rect 20720 20520 20772 20526
rect 20720 20462 20772 20468
rect 20732 20118 20760 20462
rect 20720 20112 20772 20118
rect 20720 20054 20772 20060
rect 21088 19976 21140 19982
rect 21088 19918 21140 19924
rect 20904 19568 20956 19574
rect 20904 19510 20956 19516
rect 20916 19030 20944 19510
rect 20996 19432 21048 19438
rect 20996 19374 21048 19380
rect 21008 19030 21036 19374
rect 20904 19024 20956 19030
rect 20904 18966 20956 18972
rect 20996 19024 21048 19030
rect 20996 18966 21048 18972
rect 20536 18480 20588 18486
rect 20534 18448 20536 18457
rect 20588 18448 20590 18457
rect 20534 18383 20590 18392
rect 20548 17806 20576 18383
rect 20720 18344 20772 18350
rect 20720 18286 20772 18292
rect 20536 17800 20588 17806
rect 20534 17768 20536 17777
rect 20588 17768 20590 17777
rect 20534 17703 20590 17712
rect 20732 17602 20760 18286
rect 21008 18146 21036 18966
rect 20996 18140 21048 18146
rect 20996 18082 21048 18088
rect 20720 17596 20772 17602
rect 20720 17538 20772 17544
rect 20904 17528 20956 17534
rect 20904 17470 20956 17476
rect 20916 16854 20944 17470
rect 20996 17324 21048 17330
rect 20996 17266 21048 17272
rect 20720 16848 20772 16854
rect 20718 16816 20720 16825
rect 20904 16848 20956 16854
rect 20772 16816 20774 16825
rect 20904 16790 20956 16796
rect 20718 16751 20774 16760
rect 21008 15630 21036 17266
rect 21100 16417 21128 19918
rect 21086 16408 21142 16417
rect 21086 16343 21142 16352
rect 20628 15624 20680 15630
rect 20628 15566 20680 15572
rect 20996 15624 21048 15630
rect 20996 15566 21048 15572
rect 20640 15426 20668 15566
rect 20628 15420 20680 15426
rect 20628 15362 20680 15368
rect 20996 14672 21048 14678
rect 20996 14614 21048 14620
rect 21008 14338 21036 14614
rect 20996 14332 21048 14338
rect 20996 14274 21048 14280
rect 20812 12904 20864 12910
rect 20812 12846 20864 12852
rect 20824 12502 20852 12846
rect 20812 12496 20864 12502
rect 20812 12438 20864 12444
rect 20824 12162 20852 12438
rect 20812 12156 20864 12162
rect 20812 12098 20864 12104
rect 21192 7266 21220 24526
rect 21272 24464 21324 24470
rect 21272 24406 21324 24412
rect 21180 7260 21232 7266
rect 21180 7202 21232 7208
rect 21284 6450 21312 24406
rect 21548 23240 21600 23246
rect 21548 23182 21600 23188
rect 21364 21744 21416 21750
rect 21364 21686 21416 21692
rect 21376 20905 21404 21686
rect 21362 20896 21418 20905
rect 21362 20831 21364 20840
rect 21416 20831 21418 20840
rect 21364 20802 21416 20808
rect 21364 19636 21416 19642
rect 21364 19578 21416 19584
rect 21376 18962 21404 19578
rect 21364 18956 21416 18962
rect 21364 18898 21416 18904
rect 21376 18690 21404 18898
rect 21364 18684 21416 18690
rect 21364 18626 21416 18632
rect 21364 17256 21416 17262
rect 21364 17198 21416 17204
rect 21376 15834 21404 17198
rect 21364 15828 21416 15834
rect 21364 15770 21416 15776
rect 21376 15426 21404 15770
rect 21364 15420 21416 15426
rect 21364 15362 21416 15368
rect 21560 14882 21588 23182
rect 21744 21954 21772 24542
rect 22008 22696 22060 22702
rect 22008 22638 22060 22644
rect 22020 22294 22048 22638
rect 22008 22288 22060 22294
rect 22008 22230 22060 22236
rect 21732 21948 21784 21954
rect 21732 21890 21784 21896
rect 21744 20866 21772 21890
rect 22020 21750 22048 22230
rect 22008 21744 22060 21750
rect 22008 21686 22060 21692
rect 22020 21410 22048 21686
rect 22008 21404 22060 21410
rect 22008 21346 22060 21352
rect 22020 20866 22048 21346
rect 21732 20860 21784 20866
rect 21732 20802 21784 20808
rect 22008 20860 22060 20866
rect 22008 20802 22060 20808
rect 21744 18622 21772 20802
rect 22112 19234 22140 27240
rect 22756 23586 22784 27240
rect 23202 24432 23258 24441
rect 23202 24367 23204 24376
rect 23256 24367 23258 24376
rect 23204 24338 23256 24344
rect 23296 23988 23348 23994
rect 23296 23930 23348 23936
rect 23308 23586 23336 23930
rect 22744 23580 22796 23586
rect 22744 23522 22796 23528
rect 23296 23580 23348 23586
rect 23296 23522 23348 23528
rect 23202 23480 23258 23489
rect 23202 23415 23258 23424
rect 22652 22900 22704 22906
rect 22652 22842 22704 22848
rect 22664 21954 22692 22842
rect 22744 22696 22796 22702
rect 22744 22638 22796 22644
rect 22756 22401 22784 22638
rect 22742 22392 22798 22401
rect 22742 22327 22798 22336
rect 22652 21948 22704 21954
rect 22652 21890 22704 21896
rect 22652 20180 22704 20186
rect 22652 20122 22704 20128
rect 22560 19432 22612 19438
rect 22664 19409 22692 20122
rect 22560 19374 22612 19380
rect 22650 19400 22706 19409
rect 22100 19228 22152 19234
rect 22100 19170 22152 19176
rect 22284 18888 22336 18894
rect 22284 18830 22336 18836
rect 21732 18616 21784 18622
rect 21732 18558 21784 18564
rect 21744 18185 21772 18558
rect 22296 18486 22324 18830
rect 22572 18486 22600 19374
rect 22650 19335 22706 19344
rect 23216 18865 23244 23415
rect 23492 22922 23520 27240
rect 23754 26336 23810 26345
rect 23754 26271 23810 26280
rect 23768 24470 23796 26271
rect 23940 24872 23992 24878
rect 23940 24814 23992 24820
rect 23952 24538 23980 24814
rect 23940 24532 23992 24538
rect 23940 24474 23992 24480
rect 23756 24464 23808 24470
rect 23756 24406 23808 24412
rect 23572 24328 23624 24334
rect 23572 24270 23624 24276
rect 23584 23926 23612 24270
rect 23768 24130 23796 24406
rect 23756 24124 23808 24130
rect 23676 24084 23756 24112
rect 23572 23920 23624 23926
rect 23572 23862 23624 23868
rect 23584 23042 23612 23862
rect 23676 23586 23704 24084
rect 23756 24066 23808 24072
rect 23848 24124 23900 24130
rect 23848 24066 23900 24072
rect 23756 23852 23808 23858
rect 23756 23794 23808 23800
rect 23664 23580 23716 23586
rect 23664 23522 23716 23528
rect 23664 23240 23716 23246
rect 23664 23182 23716 23188
rect 23572 23036 23624 23042
rect 23572 22978 23624 22984
rect 23492 22894 23612 22922
rect 23480 21744 23532 21750
rect 23480 21686 23532 21692
rect 23492 21614 23520 21686
rect 23480 21608 23532 21614
rect 23480 21550 23532 21556
rect 23492 21410 23520 21550
rect 23480 21404 23532 21410
rect 23480 21346 23532 21352
rect 23478 20080 23534 20089
rect 23478 20015 23480 20024
rect 23532 20015 23534 20024
rect 23480 19986 23532 19992
rect 23388 19976 23440 19982
rect 23584 19930 23612 22894
rect 23676 22838 23704 23182
rect 23768 22906 23796 23794
rect 23756 22900 23808 22906
rect 23756 22842 23808 22848
rect 23664 22832 23716 22838
rect 23664 22774 23716 22780
rect 23676 22294 23704 22774
rect 23664 22288 23716 22294
rect 23664 22230 23716 22236
rect 23860 22106 23888 24066
rect 23952 23772 23980 24474
rect 24032 23784 24084 23790
rect 23952 23744 24032 23772
rect 24032 23726 24084 23732
rect 23940 23580 23992 23586
rect 23940 23522 23992 23528
rect 23952 22106 23980 23522
rect 24044 23314 24072 23726
rect 24032 23308 24084 23314
rect 24032 23250 24084 23256
rect 23676 22078 23888 22106
rect 23943 22078 23980 22106
rect 23676 21732 23704 22078
rect 23943 21936 23971 22078
rect 23943 21908 23980 21936
rect 23676 21704 23796 21732
rect 23664 21608 23716 21614
rect 23664 21550 23716 21556
rect 23676 21206 23704 21550
rect 23664 21200 23716 21206
rect 23664 21142 23716 21148
rect 23388 19918 23440 19924
rect 23296 19228 23348 19234
rect 23296 19170 23348 19176
rect 23202 18856 23258 18865
rect 23202 18791 23258 18800
rect 22284 18480 22336 18486
rect 22284 18422 22336 18428
rect 22560 18480 22612 18486
rect 22560 18422 22612 18428
rect 22008 18344 22060 18350
rect 22008 18286 22060 18292
rect 21730 18176 21786 18185
rect 21730 18111 21786 18120
rect 21744 18078 21772 18111
rect 21732 18072 21784 18078
rect 21732 18014 21784 18020
rect 21822 17904 21878 17913
rect 21822 17839 21878 17848
rect 21836 17534 21864 17839
rect 21916 17596 21968 17602
rect 21916 17538 21968 17544
rect 21824 17528 21876 17534
rect 21824 17470 21876 17476
rect 21732 17392 21784 17398
rect 21732 17334 21784 17340
rect 21640 16848 21692 16854
rect 21640 16790 21692 16796
rect 21652 16553 21680 16790
rect 21744 16718 21772 17334
rect 21732 16712 21784 16718
rect 21732 16654 21784 16660
rect 21638 16544 21694 16553
rect 21744 16514 21772 16654
rect 21638 16479 21694 16488
rect 21732 16508 21784 16514
rect 21732 16450 21784 16456
rect 21836 16446 21864 17470
rect 21928 16514 21956 17538
rect 21916 16508 21968 16514
rect 21916 16450 21968 16456
rect 21824 16440 21876 16446
rect 21824 16382 21876 16388
rect 21548 14876 21600 14882
rect 21548 14818 21600 14824
rect 21364 14196 21416 14202
rect 21364 14138 21416 14144
rect 21376 13794 21404 14138
rect 21456 14128 21508 14134
rect 21456 14070 21508 14076
rect 21640 14128 21692 14134
rect 21640 14070 21692 14076
rect 21364 13788 21416 13794
rect 21364 13730 21416 13736
rect 21468 13590 21496 14070
rect 21456 13584 21508 13590
rect 21456 13526 21508 13532
rect 21468 13250 21496 13526
rect 21652 13522 21680 14070
rect 21640 13516 21692 13522
rect 21640 13458 21692 13464
rect 21456 13244 21508 13250
rect 21456 13186 21508 13192
rect 22020 12042 22048 18286
rect 23216 17942 23244 18791
rect 22468 17936 22520 17942
rect 22190 17904 22246 17913
rect 22468 17878 22520 17884
rect 23204 17936 23256 17942
rect 23204 17878 23256 17884
rect 22190 17839 22192 17848
rect 22244 17839 22246 17848
rect 22192 17810 22244 17816
rect 22480 17602 22508 17878
rect 22744 17800 22796 17806
rect 22744 17742 22796 17748
rect 22756 17602 22784 17742
rect 22468 17596 22520 17602
rect 22468 17538 22520 17544
rect 22744 17596 22796 17602
rect 22744 17538 22796 17544
rect 22756 16786 22784 17538
rect 23204 16916 23256 16922
rect 23204 16858 23256 16864
rect 22744 16780 22796 16786
rect 22744 16722 22796 16728
rect 23216 16718 23244 16858
rect 23204 16712 23256 16718
rect 23204 16654 23256 16660
rect 22100 16304 22152 16310
rect 22100 16246 22152 16252
rect 22112 15970 22140 16246
rect 23020 16236 23072 16242
rect 23020 16178 23072 16184
rect 22100 15964 22152 15970
rect 22100 15906 22152 15912
rect 22100 15624 22152 15630
rect 22100 15566 22152 15572
rect 22112 14202 22140 15566
rect 23032 15426 23060 16178
rect 23216 16174 23244 16654
rect 23204 16168 23256 16174
rect 23204 16110 23256 16116
rect 23112 15828 23164 15834
rect 23112 15770 23164 15776
rect 23020 15420 23072 15426
rect 23020 15362 23072 15368
rect 22926 14640 22982 14649
rect 22926 14575 22928 14584
rect 22980 14575 22982 14584
rect 22928 14546 22980 14552
rect 23032 14270 23060 15362
rect 23020 14264 23072 14270
rect 23020 14206 23072 14212
rect 23124 14202 23152 15770
rect 23216 15698 23244 16110
rect 23204 15692 23256 15698
rect 23204 15634 23256 15640
rect 22100 14196 22152 14202
rect 22100 14138 22152 14144
rect 22928 14196 22980 14202
rect 22928 14138 22980 14144
rect 23112 14196 23164 14202
rect 23112 14138 23164 14144
rect 22376 14060 22428 14066
rect 22376 14002 22428 14008
rect 22388 13522 22416 14002
rect 22376 13516 22428 13522
rect 22376 13458 22428 13464
rect 22192 13108 22244 13114
rect 22192 13050 22244 13056
rect 22020 12026 22140 12042
rect 22020 12020 22152 12026
rect 22020 12014 22100 12020
rect 22100 11962 22152 11968
rect 22008 11952 22060 11958
rect 22204 11906 22232 13050
rect 22284 12972 22336 12978
rect 22284 12914 22336 12920
rect 22296 12473 22324 12914
rect 22388 12706 22416 13458
rect 22940 13250 22968 14138
rect 23124 13794 23152 14138
rect 23112 13788 23164 13794
rect 23112 13730 23164 13736
rect 22928 13244 22980 13250
rect 22928 13186 22980 13192
rect 22468 13040 22520 13046
rect 22468 12982 22520 12988
rect 22376 12700 22428 12706
rect 22376 12642 22428 12648
rect 22480 12502 22508 12982
rect 22468 12496 22520 12502
rect 22282 12464 22338 12473
rect 22468 12438 22520 12444
rect 22282 12399 22338 12408
rect 22296 12162 22324 12399
rect 22284 12156 22336 12162
rect 22284 12098 22336 12104
rect 22560 12020 22612 12026
rect 22560 11962 22612 11968
rect 22060 11900 22232 11906
rect 22008 11894 22232 11900
rect 22020 11878 22232 11894
rect 22020 11793 22048 11878
rect 22006 11784 22062 11793
rect 22006 11719 22062 11728
rect 22572 11618 22600 11962
rect 22560 11612 22612 11618
rect 22560 11554 22612 11560
rect 23308 7826 23336 19170
rect 23400 18554 23428 19918
rect 23492 19902 23612 19930
rect 23664 19976 23716 19982
rect 23664 19918 23716 19924
rect 23492 18570 23520 19902
rect 23572 19568 23624 19574
rect 23572 19510 23624 19516
rect 23584 19234 23612 19510
rect 23572 19228 23624 19234
rect 23572 19170 23624 19176
rect 23676 19098 23704 19918
rect 23664 19092 23716 19098
rect 23664 19034 23716 19040
rect 23572 18888 23624 18894
rect 23572 18830 23624 18836
rect 23584 18690 23612 18830
rect 23572 18684 23624 18690
rect 23572 18626 23624 18632
rect 23664 18684 23716 18690
rect 23664 18626 23716 18632
rect 23388 18548 23440 18554
rect 23492 18542 23612 18570
rect 23388 18490 23440 18496
rect 23480 18072 23532 18078
rect 23480 18014 23532 18020
rect 23388 17596 23440 17602
rect 23492 17584 23520 18014
rect 23440 17556 23520 17584
rect 23388 17538 23440 17544
rect 23400 16854 23428 17538
rect 23480 17052 23532 17058
rect 23480 16994 23532 17000
rect 23388 16848 23440 16854
rect 23388 16790 23440 16796
rect 23492 16496 23520 16994
rect 23400 16468 23520 16496
rect 23400 15970 23428 16468
rect 23480 16372 23532 16378
rect 23480 16314 23532 16320
rect 23388 15964 23440 15970
rect 23388 15906 23440 15912
rect 23492 15358 23520 16314
rect 23480 15352 23532 15358
rect 23480 15294 23532 15300
rect 23584 15057 23612 18542
rect 23676 18457 23704 18626
rect 23662 18448 23718 18457
rect 23662 18383 23718 18392
rect 23676 17942 23704 18383
rect 23664 17936 23716 17942
rect 23664 17878 23716 17884
rect 23662 16816 23718 16825
rect 23662 16751 23718 16760
rect 23676 16514 23704 16751
rect 23664 16508 23716 16514
rect 23664 16450 23716 16456
rect 23664 16168 23716 16174
rect 23664 16110 23716 16116
rect 23676 15426 23704 16110
rect 23664 15420 23716 15426
rect 23664 15362 23716 15368
rect 23570 15048 23626 15057
rect 23570 14983 23626 14992
rect 23676 14898 23704 15362
rect 23584 14882 23704 14898
rect 23572 14876 23704 14882
rect 23624 14870 23704 14876
rect 23572 14818 23624 14824
rect 23664 14740 23716 14746
rect 23664 14682 23716 14688
rect 23572 14264 23624 14270
rect 23572 14206 23624 14212
rect 23480 13992 23532 13998
rect 23480 13934 23532 13940
rect 23492 12502 23520 13934
rect 23584 13726 23612 14206
rect 23572 13720 23624 13726
rect 23572 13662 23624 13668
rect 23676 13538 23704 14682
rect 23768 14678 23796 21704
rect 23952 20866 23980 21908
rect 24032 21676 24084 21682
rect 24032 21618 24084 21624
rect 24044 21410 24072 21618
rect 24032 21404 24084 21410
rect 24032 21346 24084 21352
rect 23940 20860 23992 20866
rect 23860 20820 23940 20848
rect 23860 20225 23888 20820
rect 23940 20802 23992 20808
rect 24032 20656 24084 20662
rect 24032 20598 24084 20604
rect 23940 20520 23992 20526
rect 23940 20462 23992 20468
rect 23846 20216 23902 20225
rect 23846 20151 23902 20160
rect 23952 19030 23980 20462
rect 24044 20361 24072 20598
rect 24030 20352 24086 20361
rect 24030 20287 24032 20296
rect 24084 20287 24086 20296
rect 24032 20258 24084 20264
rect 24032 19636 24084 19642
rect 24032 19578 24084 19584
rect 24044 19234 24072 19578
rect 24032 19228 24084 19234
rect 24032 19170 24084 19176
rect 23940 19024 23992 19030
rect 23940 18966 23992 18972
rect 23952 18622 23980 18966
rect 23940 18616 23992 18622
rect 23940 18558 23992 18564
rect 23938 18176 23994 18185
rect 23938 18111 23994 18120
rect 23848 17936 23900 17942
rect 23848 17878 23900 17884
rect 23860 17777 23888 17878
rect 23952 17806 23980 18111
rect 23940 17800 23992 17806
rect 23846 17768 23902 17777
rect 23940 17742 23992 17748
rect 23846 17703 23902 17712
rect 23952 17602 23980 17742
rect 23940 17596 23992 17602
rect 23940 17538 23992 17544
rect 24032 17392 24084 17398
rect 24032 17334 24084 17340
rect 24044 17058 24072 17334
rect 24032 17052 24084 17058
rect 24032 16994 24084 17000
rect 23848 16780 23900 16786
rect 23848 16722 23900 16728
rect 23756 14672 23808 14678
rect 23756 14614 23808 14620
rect 23756 14536 23808 14542
rect 23756 14478 23808 14484
rect 23584 13510 23704 13538
rect 23480 12496 23532 12502
rect 23480 12438 23532 12444
rect 23480 12360 23532 12366
rect 23480 12302 23532 12308
rect 23492 12162 23520 12302
rect 23480 12156 23532 12162
rect 23480 12098 23532 12104
rect 23308 7810 23520 7826
rect 23308 7804 23532 7810
rect 23308 7798 23480 7804
rect 23480 7746 23532 7752
rect 21640 6920 21692 6926
rect 21638 6888 21640 6897
rect 21692 6888 21694 6897
rect 21638 6823 21694 6832
rect 21272 6444 21324 6450
rect 21272 6386 21324 6392
rect 20442 5120 20498 5129
rect 20442 5055 20498 5064
rect 23478 5120 23534 5129
rect 23478 5055 23480 5064
rect 23532 5055 23534 5064
rect 23480 5026 23532 5032
rect 19062 4848 19118 4857
rect 19062 4783 19118 4792
rect 19622 4644 19918 4664
rect 19678 4642 19702 4644
rect 19758 4642 19782 4644
rect 19838 4642 19862 4644
rect 19700 4590 19702 4642
rect 19764 4590 19776 4642
rect 19838 4590 19840 4642
rect 19678 4588 19702 4590
rect 19758 4588 19782 4590
rect 19838 4588 19862 4590
rect 19622 4568 19918 4588
rect 18878 3760 18934 3769
rect 18878 3695 18934 3704
rect 19622 3556 19918 3576
rect 19678 3554 19702 3556
rect 19758 3554 19782 3556
rect 19838 3554 19862 3556
rect 19700 3502 19702 3554
rect 19764 3502 19776 3554
rect 19838 3502 19840 3554
rect 19678 3500 19702 3502
rect 19758 3500 19782 3502
rect 19838 3500 19862 3502
rect 19622 3480 19918 3500
rect 16762 2808 16818 2817
rect 16762 2743 16764 2752
rect 16816 2743 16818 2752
rect 16764 2714 16816 2720
rect 19622 2468 19918 2488
rect 19678 2466 19702 2468
rect 19758 2466 19782 2468
rect 19838 2466 19862 2468
rect 19700 2414 19702 2466
rect 19764 2414 19776 2466
rect 19838 2414 19840 2466
rect 19678 2412 19702 2414
rect 19758 2412 19782 2414
rect 19838 2412 19862 2414
rect 19622 2392 19918 2412
rect 16670 2128 16726 2137
rect 16670 2063 16726 2072
rect 15842 1312 15898 1321
rect 15842 1247 15898 1256
rect 13266 1176 13322 1185
rect 13266 1111 13322 1120
rect 23584 97 23612 13510
rect 23662 13144 23718 13153
rect 23662 13079 23718 13088
rect 23676 12706 23704 13079
rect 23664 12700 23716 12706
rect 23664 12642 23716 12648
rect 23662 11784 23718 11793
rect 23662 11719 23718 11728
rect 23676 7985 23704 11719
rect 23768 11074 23796 14478
rect 23860 11550 23888 16722
rect 24136 16700 24164 27240
rect 24780 27002 24808 27240
rect 24228 26974 24808 27002
rect 24228 24130 24256 26974
rect 24766 26880 24822 26889
rect 24766 26815 24822 26824
rect 24780 26306 24808 26815
rect 24768 26300 24820 26306
rect 24768 26242 24820 26248
rect 24766 25792 24822 25801
rect 24766 25727 24822 25736
rect 24674 25112 24730 25121
rect 24674 25047 24730 25056
rect 24289 24772 24585 24792
rect 24345 24770 24369 24772
rect 24425 24770 24449 24772
rect 24505 24770 24529 24772
rect 24367 24718 24369 24770
rect 24431 24718 24443 24770
rect 24505 24718 24507 24770
rect 24345 24716 24369 24718
rect 24425 24716 24449 24718
rect 24505 24716 24529 24718
rect 24289 24696 24585 24716
rect 24216 24124 24268 24130
rect 24216 24066 24268 24072
rect 24688 24010 24716 25047
rect 24780 24606 24808 25727
rect 24768 24600 24820 24606
rect 24768 24542 24820 24548
rect 24950 24568 25006 24577
rect 24950 24503 25006 24512
rect 24964 24470 24992 24503
rect 24952 24464 25004 24470
rect 24952 24406 25004 24412
rect 25136 24328 25188 24334
rect 25136 24270 25188 24276
rect 24688 23982 24808 24010
rect 24676 23920 24728 23926
rect 24674 23888 24676 23897
rect 24728 23888 24730 23897
rect 24674 23823 24730 23832
rect 24289 23684 24585 23704
rect 24345 23682 24369 23684
rect 24425 23682 24449 23684
rect 24505 23682 24529 23684
rect 24367 23630 24369 23682
rect 24431 23630 24443 23682
rect 24505 23630 24507 23682
rect 24345 23628 24369 23630
rect 24425 23628 24449 23630
rect 24505 23628 24529 23630
rect 24289 23608 24585 23628
rect 24688 23586 24716 23823
rect 24676 23580 24728 23586
rect 24676 23522 24728 23528
rect 24780 23466 24808 23982
rect 24688 23438 24808 23466
rect 24216 22900 24268 22906
rect 24216 22842 24268 22848
rect 24228 22158 24256 22842
rect 24289 22596 24585 22616
rect 24345 22594 24369 22596
rect 24425 22594 24449 22596
rect 24505 22594 24529 22596
rect 24367 22542 24369 22594
rect 24431 22542 24443 22594
rect 24505 22542 24507 22594
rect 24345 22540 24369 22542
rect 24425 22540 24449 22542
rect 24505 22540 24529 22542
rect 24289 22520 24585 22540
rect 24584 22288 24636 22294
rect 24688 22276 24716 23438
rect 25044 23308 25096 23314
rect 25044 23250 25096 23256
rect 25056 23042 25084 23250
rect 25044 23036 25096 23042
rect 25044 22978 25096 22984
rect 25148 22945 25176 24270
rect 25516 24146 25544 27240
rect 25686 24568 25742 24577
rect 25686 24503 25742 24512
rect 25516 24118 25636 24146
rect 25502 24024 25558 24033
rect 25502 23959 25558 23968
rect 25134 22936 25190 22945
rect 25134 22871 25190 22880
rect 25228 22492 25280 22498
rect 25228 22434 25280 22440
rect 25042 22392 25098 22401
rect 25042 22327 25098 22336
rect 24688 22248 24808 22276
rect 24584 22230 24636 22236
rect 24216 22152 24268 22158
rect 24216 22094 24268 22100
rect 24228 21750 24256 22094
rect 24596 21857 24624 22230
rect 24676 22152 24728 22158
rect 24676 22094 24728 22100
rect 24582 21848 24638 21857
rect 24582 21783 24638 21792
rect 24216 21744 24268 21750
rect 24216 21686 24268 21692
rect 24228 21410 24256 21686
rect 24289 21508 24585 21528
rect 24345 21506 24369 21508
rect 24425 21506 24449 21508
rect 24505 21506 24529 21508
rect 24367 21454 24369 21506
rect 24431 21454 24443 21506
rect 24505 21454 24507 21506
rect 24345 21452 24369 21454
rect 24425 21452 24449 21454
rect 24505 21452 24529 21454
rect 24289 21432 24585 21452
rect 24216 21404 24268 21410
rect 24216 21346 24268 21352
rect 24688 21274 24716 22094
rect 24780 21936 24808 22248
rect 24780 21908 24992 21936
rect 24766 21712 24822 21721
rect 24766 21647 24822 21656
rect 24216 21268 24268 21274
rect 24216 21210 24268 21216
rect 24676 21268 24728 21274
rect 24676 21210 24728 21216
rect 24228 18457 24256 21210
rect 24780 21177 24808 21647
rect 24860 21608 24912 21614
rect 24860 21550 24912 21556
rect 24766 21168 24822 21177
rect 24766 21103 24822 21112
rect 24676 21064 24728 21070
rect 24872 21018 24900 21550
rect 24676 21006 24728 21012
rect 24289 20420 24585 20440
rect 24345 20418 24369 20420
rect 24425 20418 24449 20420
rect 24505 20418 24529 20420
rect 24367 20366 24369 20418
rect 24431 20366 24443 20418
rect 24505 20366 24507 20418
rect 24345 20364 24369 20366
rect 24425 20364 24449 20366
rect 24505 20364 24529 20366
rect 24289 20344 24585 20364
rect 24308 20180 24360 20186
rect 24308 20122 24360 20128
rect 24320 19642 24348 20122
rect 24308 19636 24360 19642
rect 24308 19578 24360 19584
rect 24289 19332 24585 19352
rect 24345 19330 24369 19332
rect 24425 19330 24449 19332
rect 24505 19330 24529 19332
rect 24367 19278 24369 19330
rect 24431 19278 24443 19330
rect 24505 19278 24507 19330
rect 24345 19276 24369 19278
rect 24425 19276 24449 19278
rect 24505 19276 24529 19278
rect 24289 19256 24585 19276
rect 24492 19160 24544 19166
rect 24492 19102 24544 19108
rect 24308 19092 24360 19098
rect 24308 19034 24360 19040
rect 24320 18962 24348 19034
rect 24308 18956 24360 18962
rect 24308 18898 24360 18904
rect 24320 18486 24348 18898
rect 24504 18690 24532 19102
rect 24492 18684 24544 18690
rect 24492 18626 24544 18632
rect 24308 18480 24360 18486
rect 24214 18448 24270 18457
rect 24308 18422 24360 18428
rect 24214 18383 24270 18392
rect 24216 18344 24268 18350
rect 24216 18286 24268 18292
rect 24228 18010 24256 18286
rect 24289 18244 24585 18264
rect 24345 18242 24369 18244
rect 24425 18242 24449 18244
rect 24505 18242 24529 18244
rect 24367 18190 24369 18242
rect 24431 18190 24443 18242
rect 24505 18190 24507 18242
rect 24345 18188 24369 18190
rect 24425 18188 24449 18190
rect 24505 18188 24529 18190
rect 24289 18168 24585 18188
rect 24216 18004 24268 18010
rect 24216 17946 24268 17952
rect 24044 16672 24164 16700
rect 23938 16544 23994 16553
rect 23938 16479 23994 16488
rect 23952 16378 23980 16479
rect 23940 16372 23992 16378
rect 23940 16314 23992 16320
rect 24044 16258 24072 16672
rect 24228 16666 24256 17946
rect 24289 17156 24585 17176
rect 24345 17154 24369 17156
rect 24425 17154 24449 17156
rect 24505 17154 24529 17156
rect 24367 17102 24369 17154
rect 24431 17102 24443 17154
rect 24505 17102 24507 17154
rect 24345 17100 24369 17102
rect 24425 17100 24449 17102
rect 24505 17100 24529 17102
rect 24289 17080 24585 17100
rect 24584 16712 24636 16718
rect 24228 16638 24348 16666
rect 24584 16654 24636 16660
rect 24214 16544 24270 16553
rect 24214 16479 24270 16488
rect 24124 16440 24176 16446
rect 24124 16382 24176 16388
rect 23952 16230 24072 16258
rect 23848 11544 23900 11550
rect 23848 11486 23900 11492
rect 23756 11068 23808 11074
rect 23756 11010 23808 11016
rect 23952 9374 23980 16230
rect 24032 15352 24084 15358
rect 24032 15294 24084 15300
rect 24044 14814 24072 15294
rect 24136 15154 24164 16382
rect 24124 15148 24176 15154
rect 24124 15090 24176 15096
rect 24122 15048 24178 15057
rect 24122 14983 24178 14992
rect 24032 14808 24084 14814
rect 24032 14750 24084 14756
rect 24032 14672 24084 14678
rect 24032 14614 24084 14620
rect 24044 9986 24072 14614
rect 24032 9980 24084 9986
rect 24032 9922 24084 9928
rect 23940 9368 23992 9374
rect 23940 9310 23992 9316
rect 24136 8898 24164 14983
rect 24228 14814 24256 16479
rect 24320 16310 24348 16638
rect 24596 16446 24624 16654
rect 24584 16440 24636 16446
rect 24584 16382 24636 16388
rect 24308 16304 24360 16310
rect 24308 16246 24360 16252
rect 24289 16068 24585 16088
rect 24345 16066 24369 16068
rect 24425 16066 24449 16068
rect 24505 16066 24529 16068
rect 24367 16014 24369 16066
rect 24431 16014 24443 16066
rect 24505 16014 24507 16066
rect 24345 16012 24369 16014
rect 24425 16012 24449 16014
rect 24505 16012 24529 16014
rect 24289 15992 24585 16012
rect 24308 15692 24360 15698
rect 24308 15634 24360 15640
rect 24320 15222 24348 15634
rect 24688 15426 24716 21006
rect 24780 20990 24900 21018
rect 24780 17777 24808 20990
rect 24964 20730 24992 21908
rect 24952 20724 25004 20730
rect 24952 20666 25004 20672
rect 24860 20656 24912 20662
rect 24860 20598 24912 20604
rect 24872 19642 24900 20598
rect 24860 19636 24912 19642
rect 24860 19578 24912 19584
rect 25056 18554 25084 22327
rect 25240 21818 25268 22434
rect 25228 21812 25280 21818
rect 25228 21754 25280 21760
rect 25240 21410 25268 21754
rect 25228 21404 25280 21410
rect 25228 21346 25280 21352
rect 25136 20860 25188 20866
rect 25136 20802 25188 20808
rect 25148 20322 25176 20802
rect 25318 20760 25374 20769
rect 25318 20695 25320 20704
rect 25372 20695 25374 20704
rect 25320 20666 25372 20672
rect 25136 20316 25188 20322
rect 25136 20258 25188 20264
rect 25332 20118 25360 20666
rect 25320 20112 25372 20118
rect 25320 20054 25372 20060
rect 25516 20050 25544 23959
rect 25504 20044 25556 20050
rect 25504 19986 25556 19992
rect 25412 19976 25464 19982
rect 25412 19918 25464 19924
rect 25134 19672 25190 19681
rect 25134 19607 25190 19616
rect 25148 19030 25176 19607
rect 25424 19409 25452 19918
rect 25504 19432 25556 19438
rect 25410 19400 25466 19409
rect 25504 19374 25556 19380
rect 25410 19335 25466 19344
rect 25136 19024 25188 19030
rect 25136 18966 25188 18972
rect 25320 18888 25372 18894
rect 25318 18856 25320 18865
rect 25372 18856 25374 18865
rect 25318 18791 25374 18800
rect 24952 18548 25004 18554
rect 24952 18490 25004 18496
rect 25044 18548 25096 18554
rect 25044 18490 25096 18496
rect 24964 18146 24992 18490
rect 25056 18146 25084 18490
rect 25516 18486 25544 19374
rect 25504 18480 25556 18486
rect 25504 18422 25556 18428
rect 25412 18344 25464 18350
rect 25412 18286 25464 18292
rect 24952 18140 25004 18146
rect 24952 18082 25004 18088
rect 25044 18140 25096 18146
rect 25044 18082 25096 18088
rect 24766 17768 24822 17777
rect 24766 17703 24822 17712
rect 24768 17460 24820 17466
rect 24768 17402 24820 17408
rect 24780 16786 24808 17402
rect 25424 17233 25452 18286
rect 25516 18078 25544 18422
rect 25504 18072 25556 18078
rect 25504 18014 25556 18020
rect 25410 17224 25466 17233
rect 25410 17159 25466 17168
rect 25134 16952 25190 16961
rect 25134 16887 25190 16896
rect 25042 16816 25098 16825
rect 24768 16780 24820 16786
rect 25042 16751 25098 16760
rect 24768 16722 24820 16728
rect 24780 16514 24808 16722
rect 24768 16508 24820 16514
rect 24768 16450 24820 16456
rect 24780 15970 24808 16450
rect 24860 16372 24912 16378
rect 24860 16314 24912 16320
rect 24768 15964 24820 15970
rect 24768 15906 24820 15912
rect 24872 15902 24900 16314
rect 25056 15970 25084 16751
rect 25044 15964 25096 15970
rect 25044 15906 25096 15912
rect 24860 15896 24912 15902
rect 24860 15838 24912 15844
rect 24676 15420 24728 15426
rect 24676 15362 24728 15368
rect 24308 15216 24360 15222
rect 24308 15158 24360 15164
rect 24688 15034 24716 15362
rect 24768 15216 24820 15222
rect 24820 15164 24900 15170
rect 24768 15158 24900 15164
rect 24780 15142 24900 15158
rect 24688 15006 24808 15034
rect 24289 14980 24585 15000
rect 24345 14978 24369 14980
rect 24425 14978 24449 14980
rect 24505 14978 24529 14980
rect 24367 14926 24369 14978
rect 24431 14926 24443 14978
rect 24505 14926 24507 14978
rect 24345 14924 24369 14926
rect 24425 14924 24449 14926
rect 24505 14924 24529 14926
rect 24289 14904 24585 14924
rect 24674 14912 24730 14921
rect 24674 14847 24676 14856
rect 24728 14847 24730 14856
rect 24676 14818 24728 14824
rect 24216 14808 24268 14814
rect 24216 14750 24268 14756
rect 24780 14678 24808 15006
rect 24768 14672 24820 14678
rect 24768 14614 24820 14620
rect 24872 14542 24900 15142
rect 25056 14746 25084 15906
rect 25148 15290 25176 16887
rect 25412 16508 25464 16514
rect 25412 16450 25464 16456
rect 25226 16408 25282 16417
rect 25226 16343 25228 16352
rect 25280 16343 25282 16352
rect 25228 16314 25280 16320
rect 25240 15970 25268 16314
rect 25424 16009 25452 16450
rect 25410 16000 25466 16009
rect 25228 15964 25280 15970
rect 25410 15935 25466 15944
rect 25228 15906 25280 15912
rect 25410 15456 25466 15465
rect 25410 15391 25412 15400
rect 25464 15391 25466 15400
rect 25412 15362 25464 15368
rect 25136 15284 25188 15290
rect 25136 15226 25188 15232
rect 25148 14882 25176 15226
rect 25136 14876 25188 14882
rect 25136 14818 25188 14824
rect 25044 14740 25096 14746
rect 25044 14682 25096 14688
rect 24492 14536 24544 14542
rect 24492 14478 24544 14484
rect 24860 14536 24912 14542
rect 24860 14478 24912 14484
rect 24504 14338 24532 14478
rect 24858 14368 24914 14377
rect 24492 14332 24544 14338
rect 24858 14303 24914 14312
rect 24492 14274 24544 14280
rect 24289 13892 24585 13912
rect 24345 13890 24369 13892
rect 24425 13890 24449 13892
rect 24505 13890 24529 13892
rect 24367 13838 24369 13890
rect 24431 13838 24443 13890
rect 24505 13838 24507 13890
rect 24345 13836 24369 13838
rect 24425 13836 24449 13838
rect 24505 13836 24529 13838
rect 24289 13816 24585 13836
rect 24872 13794 24900 14303
rect 24860 13788 24912 13794
rect 24860 13730 24912 13736
rect 24582 13688 24638 13697
rect 24582 13623 24638 13632
rect 24766 13688 24822 13697
rect 24766 13623 24822 13632
rect 24596 13590 24624 13623
rect 24584 13584 24636 13590
rect 24584 13526 24636 13532
rect 24780 13250 24808 13623
rect 24768 13244 24820 13250
rect 24768 13186 24820 13192
rect 24584 13108 24636 13114
rect 24584 13050 24636 13056
rect 24596 13017 24624 13050
rect 24582 13008 24638 13017
rect 24638 12966 24716 12994
rect 24582 12943 24638 12952
rect 24289 12804 24585 12824
rect 24345 12802 24369 12804
rect 24425 12802 24449 12804
rect 24505 12802 24529 12804
rect 24367 12750 24369 12802
rect 24431 12750 24443 12802
rect 24505 12750 24507 12802
rect 24345 12748 24369 12750
rect 24425 12748 24449 12750
rect 24505 12748 24529 12750
rect 24289 12728 24585 12748
rect 24688 12706 24716 12966
rect 24676 12700 24728 12706
rect 24676 12642 24728 12648
rect 24768 12632 24820 12638
rect 24766 12600 24768 12609
rect 24820 12600 24822 12609
rect 24766 12535 24822 12544
rect 24768 12156 24820 12162
rect 24768 12098 24820 12104
rect 24780 12065 24808 12098
rect 24766 12056 24822 12065
rect 24676 12020 24728 12026
rect 24766 11991 24822 12000
rect 24676 11962 24728 11968
rect 24289 11716 24585 11736
rect 24345 11714 24369 11716
rect 24425 11714 24449 11716
rect 24505 11714 24529 11716
rect 24367 11662 24369 11714
rect 24431 11662 24443 11714
rect 24505 11662 24507 11714
rect 24345 11660 24369 11662
rect 24425 11660 24449 11662
rect 24505 11660 24529 11662
rect 24289 11640 24585 11660
rect 24688 11618 24716 11962
rect 24766 11648 24822 11657
rect 24676 11612 24728 11618
rect 24766 11583 24768 11592
rect 24676 11554 24728 11560
rect 24820 11583 24822 11592
rect 24768 11554 24820 11560
rect 25226 11512 25282 11521
rect 25226 11447 25228 11456
rect 25280 11447 25282 11456
rect 25228 11418 25280 11424
rect 24584 10932 24636 10938
rect 24584 10874 24636 10880
rect 24596 10841 24624 10874
rect 24582 10832 24638 10841
rect 24638 10790 24716 10818
rect 24582 10767 24638 10776
rect 24289 10628 24585 10648
rect 24345 10626 24369 10628
rect 24425 10626 24449 10628
rect 24505 10626 24529 10628
rect 24367 10574 24369 10626
rect 24431 10574 24443 10626
rect 24505 10574 24507 10626
rect 24345 10572 24369 10574
rect 24425 10572 24449 10574
rect 24505 10572 24529 10574
rect 24289 10552 24585 10572
rect 24688 10462 24716 10790
rect 25608 10569 25636 24118
rect 25700 17942 25728 24503
rect 25780 19976 25832 19982
rect 25780 19918 25832 19924
rect 25792 19642 25820 19918
rect 25780 19636 25832 19642
rect 25780 19578 25832 19584
rect 25688 17936 25740 17942
rect 25688 17878 25740 17884
rect 25792 17602 25820 19578
rect 25884 19166 25912 27359
rect 26146 27240 26202 27720
rect 26882 27240 26938 27720
rect 27526 27240 27582 27720
rect 25872 19160 25924 19166
rect 25872 19102 25924 19108
rect 25780 17596 25832 17602
rect 25780 17538 25832 17544
rect 26160 14610 26188 27240
rect 26240 16984 26292 16990
rect 26240 16926 26292 16932
rect 26148 14604 26200 14610
rect 26148 14546 26200 14552
rect 24766 10560 24822 10569
rect 24766 10495 24768 10504
rect 24820 10495 24822 10504
rect 25594 10560 25650 10569
rect 25594 10495 25650 10504
rect 24768 10466 24820 10472
rect 24676 10456 24728 10462
rect 24676 10398 24728 10404
rect 25226 10288 25282 10297
rect 25226 10223 25228 10232
rect 25280 10223 25282 10232
rect 25228 10194 25280 10200
rect 24584 9844 24636 9850
rect 24584 9786 24636 9792
rect 24596 9753 24624 9786
rect 24582 9744 24638 9753
rect 24638 9702 24716 9730
rect 24582 9679 24638 9688
rect 24289 9540 24585 9560
rect 24345 9538 24369 9540
rect 24425 9538 24449 9540
rect 24505 9538 24529 9540
rect 24367 9486 24369 9538
rect 24431 9486 24443 9538
rect 24505 9486 24507 9538
rect 24345 9484 24369 9486
rect 24425 9484 24449 9486
rect 24505 9484 24529 9486
rect 24289 9464 24585 9484
rect 24688 9442 24716 9702
rect 24676 9436 24728 9442
rect 24676 9378 24728 9384
rect 24398 9200 24454 9209
rect 24398 9135 24400 9144
rect 24452 9135 24454 9144
rect 24400 9106 24452 9112
rect 24124 8892 24176 8898
rect 24124 8834 24176 8840
rect 24400 8756 24452 8762
rect 24400 8698 24452 8704
rect 24412 8665 24440 8698
rect 24398 8656 24454 8665
rect 24398 8591 24454 8600
rect 24674 8656 24730 8665
rect 24674 8591 24730 8600
rect 24289 8452 24585 8472
rect 24345 8450 24369 8452
rect 24425 8450 24449 8452
rect 24505 8450 24529 8452
rect 24367 8398 24369 8450
rect 24431 8398 24443 8450
rect 24505 8398 24507 8450
rect 24345 8396 24369 8398
rect 24425 8396 24449 8398
rect 24505 8396 24529 8398
rect 24289 8376 24585 8396
rect 24688 8354 24716 8591
rect 24676 8348 24728 8354
rect 24676 8290 24728 8296
rect 23662 7976 23718 7985
rect 23662 7911 23718 7920
rect 24676 7668 24728 7674
rect 24676 7610 24728 7616
rect 24688 7441 24716 7610
rect 24674 7432 24730 7441
rect 24289 7364 24585 7384
rect 24674 7367 24730 7376
rect 24345 7362 24369 7364
rect 24425 7362 24449 7364
rect 24505 7362 24529 7364
rect 24367 7310 24369 7362
rect 24431 7310 24443 7362
rect 24505 7310 24507 7362
rect 24345 7308 24369 7310
rect 24425 7308 24449 7310
rect 24505 7308 24529 7310
rect 24289 7288 24585 7308
rect 24688 7266 24716 7367
rect 24676 7260 24728 7266
rect 24676 7202 24728 7208
rect 24289 6276 24585 6296
rect 24345 6274 24369 6276
rect 24425 6274 24449 6276
rect 24505 6274 24529 6276
rect 24367 6222 24369 6274
rect 24431 6222 24443 6274
rect 24505 6222 24507 6274
rect 24345 6220 24369 6222
rect 24425 6220 24449 6222
rect 24505 6220 24529 6222
rect 24289 6200 24585 6220
rect 23938 5392 23994 5401
rect 23938 5327 23994 5336
rect 23952 3497 23980 5327
rect 24289 5188 24585 5208
rect 24345 5186 24369 5188
rect 24425 5186 24449 5188
rect 24505 5186 24529 5188
rect 24367 5134 24369 5186
rect 24431 5134 24443 5186
rect 24505 5134 24507 5186
rect 24345 5132 24369 5134
rect 24425 5132 24449 5134
rect 24505 5132 24529 5134
rect 24289 5112 24585 5132
rect 25226 5120 25282 5129
rect 25226 5055 25228 5064
rect 25280 5055 25282 5064
rect 25228 5026 25280 5032
rect 25240 4886 25268 5026
rect 25228 4880 25280 4886
rect 24766 4848 24822 4857
rect 25228 4822 25280 4828
rect 24766 4783 24822 4792
rect 24582 4576 24638 4585
rect 24780 4546 24808 4783
rect 24582 4511 24638 4520
rect 24768 4540 24820 4546
rect 24596 4410 24624 4511
rect 24768 4482 24820 4488
rect 24584 4404 24636 4410
rect 24584 4346 24636 4352
rect 24596 4290 24624 4346
rect 24596 4262 24716 4290
rect 24289 4100 24585 4120
rect 24345 4098 24369 4100
rect 24425 4098 24449 4100
rect 24505 4098 24529 4100
rect 24367 4046 24369 4098
rect 24431 4046 24443 4098
rect 24505 4046 24507 4098
rect 24345 4044 24369 4046
rect 24425 4044 24449 4046
rect 24505 4044 24529 4046
rect 24289 4024 24585 4044
rect 24688 4002 24716 4262
rect 25226 4032 25282 4041
rect 24676 3996 24728 4002
rect 25226 3967 25282 3976
rect 24676 3938 24728 3944
rect 25240 3866 25268 3967
rect 25228 3860 25280 3866
rect 25228 3802 25280 3808
rect 24766 3760 24822 3769
rect 24766 3695 24822 3704
rect 24780 3662 24808 3695
rect 24768 3656 24820 3662
rect 24768 3598 24820 3604
rect 23938 3488 23994 3497
rect 23938 3423 23994 3432
rect 26252 3089 26280 16926
rect 26896 11657 26924 27240
rect 27540 16990 27568 27240
rect 27528 16984 27580 16990
rect 27528 16926 27580 16932
rect 26882 11648 26938 11657
rect 26882 11583 26938 11592
rect 24766 3080 24822 3089
rect 24289 3012 24585 3032
rect 24766 3015 24822 3024
rect 26238 3080 26294 3089
rect 26238 3015 26294 3024
rect 24345 3010 24369 3012
rect 24425 3010 24449 3012
rect 24505 3010 24529 3012
rect 24367 2958 24369 3010
rect 24431 2958 24443 3010
rect 24505 2958 24507 3010
rect 24345 2956 24369 2958
rect 24425 2956 24449 2958
rect 24505 2956 24529 2958
rect 24289 2936 24585 2956
rect 24780 2914 24808 3015
rect 24768 2908 24820 2914
rect 24768 2850 24820 2856
rect 24676 2704 24728 2710
rect 24676 2646 24728 2652
rect 24289 1924 24585 1944
rect 24345 1922 24369 1924
rect 24425 1922 24449 1924
rect 24505 1922 24529 1924
rect 24367 1870 24369 1922
rect 24431 1870 24443 1922
rect 24505 1870 24507 1922
rect 24345 1868 24369 1870
rect 24425 1868 24449 1870
rect 24505 1868 24529 1870
rect 24289 1848 24585 1868
rect 24688 641 24716 2646
rect 25228 2228 25280 2234
rect 25228 2170 25280 2176
rect 24766 2128 24822 2137
rect 24766 2063 24768 2072
rect 24820 2063 24822 2072
rect 24768 2034 24820 2040
rect 25240 2030 25268 2170
rect 25228 2024 25280 2030
rect 25228 1966 25280 1972
rect 25240 1729 25268 1966
rect 25226 1720 25282 1729
rect 25226 1655 25282 1664
rect 24674 632 24730 641
rect 24674 567 24730 576
rect 23570 88 23626 97
rect 23570 23 23626 32
<< via2 >>
rect 25870 27368 25926 27424
rect 938 20024 994 20080
rect 2318 21248 2374 21304
rect 1582 18528 1638 18584
rect 3698 20160 3754 20216
rect 5622 24770 5678 24772
rect 5702 24770 5758 24772
rect 5782 24770 5838 24772
rect 5862 24770 5918 24772
rect 5622 24718 5648 24770
rect 5648 24718 5678 24770
rect 5702 24718 5712 24770
rect 5712 24718 5758 24770
rect 5782 24718 5828 24770
rect 5828 24718 5838 24770
rect 5862 24718 5892 24770
rect 5892 24718 5918 24770
rect 5622 24716 5678 24718
rect 5702 24716 5758 24718
rect 5782 24716 5838 24718
rect 5862 24716 5918 24718
rect 6366 24376 6422 24432
rect 5998 23832 6054 23888
rect 5622 23682 5678 23684
rect 5702 23682 5758 23684
rect 5782 23682 5838 23684
rect 5862 23682 5918 23684
rect 5622 23630 5648 23682
rect 5648 23630 5678 23682
rect 5702 23630 5712 23682
rect 5712 23630 5758 23682
rect 5782 23630 5828 23682
rect 5828 23630 5838 23682
rect 5862 23630 5892 23682
rect 5892 23630 5918 23682
rect 5622 23628 5678 23630
rect 5702 23628 5758 23630
rect 5782 23628 5838 23630
rect 5862 23628 5918 23630
rect 7102 23288 7158 23344
rect 8390 22880 8446 22936
rect 7746 22744 7802 22800
rect 5622 22594 5678 22596
rect 5702 22594 5758 22596
rect 5782 22594 5838 22596
rect 5862 22594 5918 22596
rect 5622 22542 5648 22594
rect 5648 22542 5678 22594
rect 5702 22542 5712 22594
rect 5712 22542 5758 22594
rect 5782 22542 5828 22594
rect 5828 22542 5838 22594
rect 5862 22542 5892 22594
rect 5892 22542 5918 22594
rect 5622 22540 5678 22542
rect 5702 22540 5758 22542
rect 5782 22540 5838 22542
rect 5862 22540 5918 22542
rect 4986 22336 5042 22392
rect 5622 21506 5678 21508
rect 5702 21506 5758 21508
rect 5782 21506 5838 21508
rect 5862 21506 5918 21508
rect 5622 21454 5648 21506
rect 5648 21454 5678 21506
rect 5702 21454 5712 21506
rect 5712 21454 5758 21506
rect 5782 21454 5828 21506
rect 5828 21454 5838 21506
rect 5862 21454 5892 21506
rect 5892 21454 5918 21506
rect 5622 21452 5678 21454
rect 5702 21452 5758 21454
rect 5782 21452 5838 21454
rect 5862 21452 5918 21454
rect 10289 25314 10345 25316
rect 10369 25314 10425 25316
rect 10449 25314 10505 25316
rect 10529 25314 10585 25316
rect 10289 25262 10315 25314
rect 10315 25262 10345 25314
rect 10369 25262 10379 25314
rect 10379 25262 10425 25314
rect 10449 25262 10495 25314
rect 10495 25262 10505 25314
rect 10529 25262 10559 25314
rect 10559 25262 10585 25314
rect 10289 25260 10345 25262
rect 10369 25260 10425 25262
rect 10449 25260 10505 25262
rect 10529 25260 10585 25262
rect 10289 24226 10345 24228
rect 10369 24226 10425 24228
rect 10449 24226 10505 24228
rect 10529 24226 10585 24228
rect 10289 24174 10315 24226
rect 10315 24174 10345 24226
rect 10369 24174 10379 24226
rect 10379 24174 10425 24226
rect 10449 24174 10495 24226
rect 10495 24174 10505 24226
rect 10529 24174 10559 24226
rect 10559 24174 10585 24226
rect 10289 24172 10345 24174
rect 10369 24172 10425 24174
rect 10449 24172 10505 24174
rect 10529 24172 10585 24174
rect 10966 23188 10968 23208
rect 10968 23188 11020 23208
rect 11020 23188 11022 23208
rect 5622 20418 5678 20420
rect 5702 20418 5758 20420
rect 5782 20418 5838 20420
rect 5862 20418 5918 20420
rect 5622 20366 5648 20418
rect 5648 20366 5678 20418
rect 5702 20366 5712 20418
rect 5712 20366 5758 20418
rect 5782 20366 5828 20418
rect 5828 20366 5838 20418
rect 5862 20366 5892 20418
rect 5892 20366 5918 20418
rect 5622 20364 5678 20366
rect 5702 20364 5758 20366
rect 5782 20364 5838 20366
rect 5862 20364 5918 20366
rect 5622 19330 5678 19332
rect 5702 19330 5758 19332
rect 5782 19330 5838 19332
rect 5862 19330 5918 19332
rect 5622 19278 5648 19330
rect 5648 19278 5678 19330
rect 5702 19278 5712 19330
rect 5712 19278 5758 19330
rect 5782 19278 5828 19330
rect 5828 19278 5838 19330
rect 5862 19278 5892 19330
rect 5892 19278 5918 19330
rect 5622 19276 5678 19278
rect 5702 19276 5758 19278
rect 5782 19276 5838 19278
rect 5862 19276 5918 19278
rect 10966 23152 11022 23188
rect 10289 23138 10345 23140
rect 10369 23138 10425 23140
rect 10449 23138 10505 23140
rect 10529 23138 10585 23140
rect 10289 23086 10315 23138
rect 10315 23086 10345 23138
rect 10369 23086 10379 23138
rect 10379 23086 10425 23138
rect 10449 23086 10495 23138
rect 10495 23086 10505 23138
rect 10529 23086 10559 23138
rect 10559 23086 10585 23138
rect 10289 23084 10345 23086
rect 10369 23084 10425 23086
rect 10449 23084 10505 23086
rect 10529 23084 10585 23086
rect 10289 22050 10345 22052
rect 10369 22050 10425 22052
rect 10449 22050 10505 22052
rect 10529 22050 10585 22052
rect 10289 21998 10315 22050
rect 10315 21998 10345 22050
rect 10369 21998 10379 22050
rect 10379 21998 10425 22050
rect 10449 21998 10495 22050
rect 10495 21998 10505 22050
rect 10529 21998 10559 22050
rect 10559 21998 10585 22050
rect 10289 21996 10345 21998
rect 10369 21996 10425 21998
rect 10449 21996 10505 21998
rect 10529 21996 10585 21998
rect 10046 21792 10102 21848
rect 10598 21792 10654 21848
rect 10289 20962 10345 20964
rect 10369 20962 10425 20964
rect 10449 20962 10505 20964
rect 10529 20962 10585 20964
rect 10289 20910 10315 20962
rect 10315 20910 10345 20962
rect 10369 20910 10379 20962
rect 10379 20910 10425 20962
rect 10449 20910 10495 20962
rect 10495 20910 10505 20962
rect 10529 20910 10559 20962
rect 10559 20910 10585 20962
rect 10289 20908 10345 20910
rect 10369 20908 10425 20910
rect 10449 20908 10505 20910
rect 10529 20908 10585 20910
rect 13174 24512 13230 24568
rect 12530 23016 12586 23072
rect 12346 20976 12402 21032
rect 12070 20704 12126 20760
rect 10289 19874 10345 19876
rect 10369 19874 10425 19876
rect 10449 19874 10505 19876
rect 10529 19874 10585 19876
rect 10289 19822 10315 19874
rect 10315 19822 10345 19874
rect 10369 19822 10379 19874
rect 10379 19822 10425 19874
rect 10449 19822 10495 19874
rect 10495 19822 10505 19874
rect 10529 19822 10559 19874
rect 10559 19822 10585 19874
rect 10289 19820 10345 19822
rect 10369 19820 10425 19822
rect 10449 19820 10505 19822
rect 10529 19820 10585 19822
rect 11242 20160 11298 20216
rect 11150 19752 11206 19808
rect 9862 19072 9918 19128
rect 4342 18936 4398 18992
rect 10289 18786 10345 18788
rect 10369 18786 10425 18788
rect 10449 18786 10505 18788
rect 10529 18786 10585 18788
rect 10289 18734 10315 18786
rect 10315 18734 10345 18786
rect 10369 18734 10379 18786
rect 10379 18734 10425 18786
rect 10449 18734 10495 18786
rect 10495 18734 10505 18786
rect 10529 18734 10559 18786
rect 10559 18734 10585 18786
rect 10289 18732 10345 18734
rect 10369 18732 10425 18734
rect 10449 18732 10505 18734
rect 10529 18732 10585 18734
rect 10874 18292 10876 18312
rect 10876 18292 10928 18312
rect 10928 18292 10930 18312
rect 10874 18256 10930 18292
rect 5622 18242 5678 18244
rect 5702 18242 5758 18244
rect 5782 18242 5838 18244
rect 5862 18242 5918 18244
rect 5622 18190 5648 18242
rect 5648 18190 5678 18242
rect 5702 18190 5712 18242
rect 5712 18190 5758 18242
rect 5782 18190 5828 18242
rect 5828 18190 5838 18242
rect 5862 18190 5892 18242
rect 5892 18190 5918 18242
rect 5622 18188 5678 18190
rect 5702 18188 5758 18190
rect 5782 18188 5838 18190
rect 5862 18188 5918 18190
rect 2962 17848 3018 17904
rect 10289 17698 10345 17700
rect 10369 17698 10425 17700
rect 10449 17698 10505 17700
rect 10529 17698 10585 17700
rect 10289 17646 10315 17698
rect 10315 17646 10345 17698
rect 10369 17646 10379 17698
rect 10379 17646 10425 17698
rect 10449 17646 10495 17698
rect 10495 17646 10505 17698
rect 10529 17646 10559 17698
rect 10559 17646 10585 17698
rect 10289 17644 10345 17646
rect 10369 17644 10425 17646
rect 10449 17644 10505 17646
rect 10529 17644 10585 17646
rect 5622 17154 5678 17156
rect 5702 17154 5758 17156
rect 5782 17154 5838 17156
rect 5862 17154 5918 17156
rect 5622 17102 5648 17154
rect 5648 17102 5678 17154
rect 5702 17102 5712 17154
rect 5712 17102 5758 17154
rect 5782 17102 5828 17154
rect 5828 17102 5838 17154
rect 5862 17102 5892 17154
rect 5892 17102 5918 17154
rect 5622 17100 5678 17102
rect 5702 17100 5758 17102
rect 5782 17100 5838 17102
rect 5862 17100 5918 17102
rect 10289 16610 10345 16612
rect 10369 16610 10425 16612
rect 10449 16610 10505 16612
rect 10529 16610 10585 16612
rect 10289 16558 10315 16610
rect 10315 16558 10345 16610
rect 10369 16558 10379 16610
rect 10379 16558 10425 16610
rect 10449 16558 10495 16610
rect 10495 16558 10505 16610
rect 10529 16558 10559 16610
rect 10559 16558 10585 16610
rect 10289 16556 10345 16558
rect 10369 16556 10425 16558
rect 10449 16556 10505 16558
rect 10529 16556 10585 16558
rect 5622 16066 5678 16068
rect 5702 16066 5758 16068
rect 5782 16066 5838 16068
rect 5862 16066 5918 16068
rect 5622 16014 5648 16066
rect 5648 16014 5678 16066
rect 5702 16014 5712 16066
rect 5712 16014 5758 16066
rect 5782 16014 5828 16066
rect 5828 16014 5838 16066
rect 5862 16014 5892 16066
rect 5892 16014 5918 16066
rect 5622 16012 5678 16014
rect 5702 16012 5758 16014
rect 5782 16012 5838 16014
rect 5862 16012 5918 16014
rect 11794 18256 11850 18312
rect 12438 18256 12494 18312
rect 10289 15522 10345 15524
rect 10369 15522 10425 15524
rect 10449 15522 10505 15524
rect 10529 15522 10585 15524
rect 10289 15470 10315 15522
rect 10315 15470 10345 15522
rect 10369 15470 10379 15522
rect 10379 15470 10425 15522
rect 10449 15470 10495 15522
rect 10495 15470 10505 15522
rect 10529 15470 10559 15522
rect 10559 15470 10585 15522
rect 10289 15468 10345 15470
rect 10369 15468 10425 15470
rect 10449 15468 10505 15470
rect 10529 15468 10585 15470
rect 5622 14978 5678 14980
rect 5702 14978 5758 14980
rect 5782 14978 5838 14980
rect 5862 14978 5918 14980
rect 5622 14926 5648 14978
rect 5648 14926 5678 14978
rect 5702 14926 5712 14978
rect 5712 14926 5758 14978
rect 5782 14926 5828 14978
rect 5828 14926 5838 14978
rect 5862 14926 5892 14978
rect 5892 14926 5918 14978
rect 5622 14924 5678 14926
rect 5702 14924 5758 14926
rect 5782 14924 5838 14926
rect 5862 14924 5918 14926
rect 12622 20588 12678 20624
rect 12622 20568 12624 20588
rect 12624 20568 12676 20588
rect 12676 20568 12678 20588
rect 13634 21792 13690 21848
rect 13634 19616 13690 19672
rect 13542 18664 13598 18720
rect 13450 17868 13506 17904
rect 13450 17848 13452 17868
rect 13452 17848 13504 17868
rect 13504 17848 13506 17868
rect 14094 23016 14150 23072
rect 14278 23016 14334 23072
rect 14278 22900 14334 22936
rect 14278 22880 14280 22900
rect 14280 22880 14332 22900
rect 14332 22880 14334 22900
rect 14956 24770 15012 24772
rect 15036 24770 15092 24772
rect 15116 24770 15172 24772
rect 15196 24770 15252 24772
rect 14956 24718 14982 24770
rect 14982 24718 15012 24770
rect 15036 24718 15046 24770
rect 15046 24718 15092 24770
rect 15116 24718 15162 24770
rect 15162 24718 15172 24770
rect 15196 24718 15226 24770
rect 15226 24718 15252 24770
rect 14956 24716 15012 24718
rect 15036 24716 15092 24718
rect 15116 24716 15172 24718
rect 15196 24716 15252 24718
rect 15106 23832 15162 23888
rect 14956 23682 15012 23684
rect 15036 23682 15092 23684
rect 15116 23682 15172 23684
rect 15196 23682 15252 23684
rect 14956 23630 14982 23682
rect 14982 23630 15012 23682
rect 15036 23630 15046 23682
rect 15046 23630 15092 23682
rect 15116 23630 15162 23682
rect 15162 23630 15172 23682
rect 15196 23630 15226 23682
rect 15226 23630 15252 23682
rect 14956 23628 15012 23630
rect 15036 23628 15092 23630
rect 15116 23628 15172 23630
rect 15196 23628 15252 23630
rect 14956 22594 15012 22596
rect 15036 22594 15092 22596
rect 15116 22594 15172 22596
rect 15196 22594 15252 22596
rect 14956 22542 14982 22594
rect 14982 22542 15012 22594
rect 15036 22542 15046 22594
rect 15046 22542 15092 22594
rect 15116 22542 15162 22594
rect 15162 22542 15172 22594
rect 15196 22542 15226 22594
rect 15226 22542 15252 22594
rect 14956 22540 15012 22542
rect 15036 22540 15092 22542
rect 15116 22540 15172 22542
rect 15196 22540 15252 22542
rect 14956 21506 15012 21508
rect 15036 21506 15092 21508
rect 15116 21506 15172 21508
rect 15196 21506 15252 21508
rect 14956 21454 14982 21506
rect 14982 21454 15012 21506
rect 15036 21454 15046 21506
rect 15046 21454 15092 21506
rect 15116 21454 15162 21506
rect 15162 21454 15172 21506
rect 15196 21454 15226 21506
rect 15226 21454 15252 21506
rect 14956 21452 15012 21454
rect 15036 21452 15092 21454
rect 15116 21452 15172 21454
rect 15196 21452 15252 21454
rect 14956 20418 15012 20420
rect 15036 20418 15092 20420
rect 15116 20418 15172 20420
rect 15196 20418 15252 20420
rect 14956 20366 14982 20418
rect 14982 20366 15012 20418
rect 15036 20366 15046 20418
rect 15046 20366 15092 20418
rect 15116 20366 15162 20418
rect 15162 20366 15172 20418
rect 15196 20366 15226 20418
rect 15226 20366 15252 20418
rect 14956 20364 15012 20366
rect 15036 20364 15092 20366
rect 15116 20364 15172 20366
rect 15196 20364 15252 20366
rect 13910 17984 13966 18040
rect 14956 19330 15012 19332
rect 15036 19330 15092 19332
rect 15116 19330 15172 19332
rect 15196 19330 15252 19332
rect 14956 19278 14982 19330
rect 14982 19278 15012 19330
rect 15036 19278 15046 19330
rect 15046 19278 15092 19330
rect 15116 19278 15162 19330
rect 15162 19278 15172 19330
rect 15196 19278 15226 19330
rect 15226 19278 15252 19330
rect 14956 19276 15012 19278
rect 15036 19276 15092 19278
rect 15116 19276 15172 19278
rect 15196 19276 15252 19278
rect 16118 22780 16120 22800
rect 16120 22780 16172 22800
rect 16172 22780 16174 22800
rect 16118 22744 16174 22780
rect 16302 21384 16358 21440
rect 16026 21248 16082 21304
rect 16394 19772 16450 19808
rect 16394 19752 16396 19772
rect 16396 19752 16448 19772
rect 16448 19752 16450 19772
rect 14738 19072 14794 19128
rect 15290 19072 15346 19128
rect 12254 14584 12310 14640
rect 10289 14434 10345 14436
rect 10369 14434 10425 14436
rect 10449 14434 10505 14436
rect 10529 14434 10585 14436
rect 10289 14382 10315 14434
rect 10315 14382 10345 14434
rect 10369 14382 10379 14434
rect 10379 14382 10425 14434
rect 10449 14382 10495 14434
rect 10495 14382 10505 14434
rect 10529 14382 10559 14434
rect 10559 14382 10585 14434
rect 10289 14380 10345 14382
rect 10369 14380 10425 14382
rect 10449 14380 10505 14382
rect 10529 14380 10585 14382
rect 5622 13890 5678 13892
rect 5702 13890 5758 13892
rect 5782 13890 5838 13892
rect 5862 13890 5918 13892
rect 5622 13838 5648 13890
rect 5648 13838 5678 13890
rect 5702 13838 5712 13890
rect 5712 13838 5758 13890
rect 5782 13838 5828 13890
rect 5828 13838 5838 13890
rect 5862 13838 5892 13890
rect 5892 13838 5918 13890
rect 5622 13836 5678 13838
rect 5702 13836 5758 13838
rect 5782 13836 5838 13838
rect 5862 13836 5918 13838
rect 1490 13632 1546 13688
rect 386 13088 442 13144
rect 2778 13496 2834 13552
rect 11702 13532 11704 13552
rect 11704 13532 11756 13552
rect 11756 13532 11758 13552
rect 11702 13496 11758 13532
rect 10289 13346 10345 13348
rect 10369 13346 10425 13348
rect 10449 13346 10505 13348
rect 10529 13346 10585 13348
rect 10289 13294 10315 13346
rect 10315 13294 10345 13346
rect 10369 13294 10379 13346
rect 10379 13294 10425 13346
rect 10449 13294 10495 13346
rect 10495 13294 10505 13346
rect 10529 13294 10559 13346
rect 10559 13294 10585 13346
rect 10289 13292 10345 13294
rect 10369 13292 10425 13294
rect 10449 13292 10505 13294
rect 10529 13292 10585 13294
rect 15014 18956 15070 18992
rect 15014 18936 15016 18956
rect 15016 18936 15068 18956
rect 15068 18936 15070 18956
rect 14956 18242 15012 18244
rect 15036 18242 15092 18244
rect 15116 18242 15172 18244
rect 15196 18242 15252 18244
rect 14956 18190 14982 18242
rect 14982 18190 15012 18242
rect 15036 18190 15046 18242
rect 15046 18190 15092 18242
rect 15116 18190 15162 18242
rect 15162 18190 15172 18242
rect 15196 18190 15226 18242
rect 15226 18190 15252 18242
rect 14956 18188 15012 18190
rect 15036 18188 15092 18190
rect 15116 18188 15172 18190
rect 15196 18188 15252 18190
rect 16394 18392 16450 18448
rect 15106 17476 15108 17496
rect 15108 17476 15160 17496
rect 15160 17476 15162 17496
rect 15106 17440 15162 17476
rect 14956 17154 15012 17156
rect 15036 17154 15092 17156
rect 15116 17154 15172 17156
rect 15196 17154 15252 17156
rect 14956 17102 14982 17154
rect 14982 17102 15012 17154
rect 15036 17102 15046 17154
rect 15046 17102 15092 17154
rect 15116 17102 15162 17154
rect 15162 17102 15172 17154
rect 15196 17102 15226 17154
rect 15226 17102 15252 17154
rect 14956 17100 15012 17102
rect 15036 17100 15092 17102
rect 15116 17100 15172 17102
rect 15196 17100 15252 17102
rect 15474 16896 15530 16952
rect 15750 16796 15752 16816
rect 15752 16796 15804 16816
rect 15804 16796 15806 16816
rect 15750 16760 15806 16796
rect 14956 16066 15012 16068
rect 15036 16066 15092 16068
rect 15116 16066 15172 16068
rect 15196 16066 15252 16068
rect 14956 16014 14982 16066
rect 14982 16014 15012 16066
rect 15036 16014 15046 16066
rect 15046 16014 15092 16066
rect 15116 16014 15162 16066
rect 15162 16014 15172 16066
rect 15196 16014 15226 16066
rect 15226 16014 15252 16066
rect 14956 16012 15012 16014
rect 15036 16012 15092 16014
rect 15116 16012 15172 16014
rect 15196 16012 15252 16014
rect 14956 14978 15012 14980
rect 15036 14978 15092 14980
rect 15116 14978 15172 14980
rect 15196 14978 15252 14980
rect 14956 14926 14982 14978
rect 14982 14926 15012 14978
rect 15036 14926 15046 14978
rect 15046 14926 15092 14978
rect 15116 14926 15162 14978
rect 15162 14926 15172 14978
rect 15196 14926 15226 14978
rect 15226 14926 15252 14978
rect 14956 14924 15012 14926
rect 15036 14924 15092 14926
rect 15116 14924 15172 14926
rect 15196 14924 15252 14926
rect 14956 13890 15012 13892
rect 15036 13890 15092 13892
rect 15116 13890 15172 13892
rect 15196 13890 15252 13892
rect 14956 13838 14982 13890
rect 14982 13838 15012 13890
rect 15036 13838 15046 13890
rect 15046 13838 15092 13890
rect 15116 13838 15162 13890
rect 15162 13838 15172 13890
rect 15196 13838 15226 13890
rect 15226 13838 15252 13890
rect 14956 13836 15012 13838
rect 15036 13836 15092 13838
rect 15116 13836 15172 13838
rect 15196 13836 15252 13838
rect 14370 13632 14426 13688
rect 13358 13088 13414 13144
rect 2042 12952 2098 13008
rect 2870 12952 2926 13008
rect 12070 12952 12126 13008
rect 5622 12802 5678 12804
rect 5702 12802 5758 12804
rect 5782 12802 5838 12804
rect 5862 12802 5918 12804
rect 5622 12750 5648 12802
rect 5648 12750 5678 12802
rect 5702 12750 5712 12802
rect 5712 12750 5758 12802
rect 5782 12750 5828 12802
rect 5828 12750 5838 12802
rect 5862 12750 5892 12802
rect 5892 12750 5918 12802
rect 5622 12748 5678 12750
rect 5702 12748 5758 12750
rect 5782 12748 5838 12750
rect 5862 12748 5918 12750
rect 10289 12258 10345 12260
rect 10369 12258 10425 12260
rect 10449 12258 10505 12260
rect 10529 12258 10585 12260
rect 10289 12206 10315 12258
rect 10315 12206 10345 12258
rect 10369 12206 10379 12258
rect 10379 12206 10425 12258
rect 10449 12206 10495 12258
rect 10495 12206 10505 12258
rect 10529 12206 10559 12258
rect 10559 12206 10585 12258
rect 10289 12204 10345 12206
rect 10369 12204 10425 12206
rect 10449 12204 10505 12206
rect 10529 12204 10585 12206
rect 5622 11714 5678 11716
rect 5702 11714 5758 11716
rect 5782 11714 5838 11716
rect 5862 11714 5918 11716
rect 5622 11662 5648 11714
rect 5648 11662 5678 11714
rect 5702 11662 5712 11714
rect 5712 11662 5758 11714
rect 5782 11662 5828 11714
rect 5828 11662 5838 11714
rect 5862 11662 5892 11714
rect 5892 11662 5918 11714
rect 5622 11660 5678 11662
rect 5702 11660 5758 11662
rect 5782 11660 5838 11662
rect 5862 11660 5918 11662
rect 10289 11170 10345 11172
rect 10369 11170 10425 11172
rect 10449 11170 10505 11172
rect 10529 11170 10585 11172
rect 10289 11118 10315 11170
rect 10315 11118 10345 11170
rect 10369 11118 10379 11170
rect 10379 11118 10425 11170
rect 10449 11118 10495 11170
rect 10495 11118 10505 11170
rect 10529 11118 10559 11170
rect 10559 11118 10585 11170
rect 10289 11116 10345 11118
rect 10369 11116 10425 11118
rect 10449 11116 10505 11118
rect 10529 11116 10585 11118
rect 5622 10626 5678 10628
rect 5702 10626 5758 10628
rect 5782 10626 5838 10628
rect 5862 10626 5918 10628
rect 5622 10574 5648 10626
rect 5648 10574 5678 10626
rect 5702 10574 5712 10626
rect 5712 10574 5758 10626
rect 5782 10574 5828 10626
rect 5828 10574 5838 10626
rect 5862 10574 5892 10626
rect 5892 10574 5918 10626
rect 5622 10572 5678 10574
rect 5702 10572 5758 10574
rect 5782 10572 5838 10574
rect 5862 10572 5918 10574
rect 10289 10082 10345 10084
rect 10369 10082 10425 10084
rect 10449 10082 10505 10084
rect 10529 10082 10585 10084
rect 10289 10030 10315 10082
rect 10315 10030 10345 10082
rect 10369 10030 10379 10082
rect 10379 10030 10425 10082
rect 10449 10030 10495 10082
rect 10495 10030 10505 10082
rect 10529 10030 10559 10082
rect 10559 10030 10585 10082
rect 10289 10028 10345 10030
rect 10369 10028 10425 10030
rect 10449 10028 10505 10030
rect 10529 10028 10585 10030
rect 5622 9538 5678 9540
rect 5702 9538 5758 9540
rect 5782 9538 5838 9540
rect 5862 9538 5918 9540
rect 5622 9486 5648 9538
rect 5648 9486 5678 9538
rect 5702 9486 5712 9538
rect 5712 9486 5758 9538
rect 5782 9486 5828 9538
rect 5828 9486 5838 9538
rect 5862 9486 5892 9538
rect 5892 9486 5918 9538
rect 5622 9484 5678 9486
rect 5702 9484 5758 9486
rect 5782 9484 5838 9486
rect 5862 9484 5918 9486
rect 10289 8994 10345 8996
rect 10369 8994 10425 8996
rect 10449 8994 10505 8996
rect 10529 8994 10585 8996
rect 10289 8942 10315 8994
rect 10315 8942 10345 8994
rect 10369 8942 10379 8994
rect 10379 8942 10425 8994
rect 10449 8942 10495 8994
rect 10495 8942 10505 8994
rect 10529 8942 10559 8994
rect 10559 8942 10585 8994
rect 10289 8940 10345 8942
rect 10369 8940 10425 8942
rect 10449 8940 10505 8942
rect 10529 8940 10585 8942
rect 5622 8450 5678 8452
rect 5702 8450 5758 8452
rect 5782 8450 5838 8452
rect 5862 8450 5918 8452
rect 5622 8398 5648 8450
rect 5648 8398 5678 8450
rect 5702 8398 5712 8450
rect 5712 8398 5758 8450
rect 5782 8398 5828 8450
rect 5828 8398 5838 8450
rect 5862 8398 5892 8450
rect 5892 8398 5918 8450
rect 5622 8396 5678 8398
rect 5702 8396 5758 8398
rect 5782 8396 5838 8398
rect 5862 8396 5918 8398
rect 10289 7906 10345 7908
rect 10369 7906 10425 7908
rect 10449 7906 10505 7908
rect 10529 7906 10585 7908
rect 10289 7854 10315 7906
rect 10315 7854 10345 7906
rect 10369 7854 10379 7906
rect 10379 7854 10425 7906
rect 10449 7854 10495 7906
rect 10495 7854 10505 7906
rect 10529 7854 10559 7906
rect 10559 7854 10585 7906
rect 10289 7852 10345 7854
rect 10369 7852 10425 7854
rect 10449 7852 10505 7854
rect 10529 7852 10585 7854
rect 5622 7362 5678 7364
rect 5702 7362 5758 7364
rect 5782 7362 5838 7364
rect 5862 7362 5918 7364
rect 5622 7310 5648 7362
rect 5648 7310 5678 7362
rect 5702 7310 5712 7362
rect 5712 7310 5758 7362
rect 5782 7310 5828 7362
rect 5828 7310 5838 7362
rect 5862 7310 5892 7362
rect 5892 7310 5918 7362
rect 5622 7308 5678 7310
rect 5702 7308 5758 7310
rect 5782 7308 5838 7310
rect 5862 7308 5918 7310
rect 10289 6818 10345 6820
rect 10369 6818 10425 6820
rect 10449 6818 10505 6820
rect 10529 6818 10585 6820
rect 10289 6766 10315 6818
rect 10315 6766 10345 6818
rect 10369 6766 10379 6818
rect 10379 6766 10425 6818
rect 10449 6766 10495 6818
rect 10495 6766 10505 6818
rect 10529 6766 10559 6818
rect 10559 6766 10585 6818
rect 10289 6764 10345 6766
rect 10369 6764 10425 6766
rect 10449 6764 10505 6766
rect 10529 6764 10585 6766
rect 5622 6274 5678 6276
rect 5702 6274 5758 6276
rect 5782 6274 5838 6276
rect 5862 6274 5918 6276
rect 5622 6222 5648 6274
rect 5648 6222 5678 6274
rect 5702 6222 5712 6274
rect 5712 6222 5758 6274
rect 5782 6222 5828 6274
rect 5828 6222 5838 6274
rect 5862 6222 5892 6274
rect 5892 6222 5918 6274
rect 5622 6220 5678 6222
rect 5702 6220 5758 6222
rect 5782 6220 5838 6222
rect 5862 6220 5918 6222
rect 10289 5730 10345 5732
rect 10369 5730 10425 5732
rect 10449 5730 10505 5732
rect 10529 5730 10585 5732
rect 10289 5678 10315 5730
rect 10315 5678 10345 5730
rect 10369 5678 10379 5730
rect 10379 5678 10425 5730
rect 10449 5678 10495 5730
rect 10495 5678 10505 5730
rect 10529 5678 10559 5730
rect 10559 5678 10585 5730
rect 10289 5676 10345 5678
rect 10369 5676 10425 5678
rect 10449 5676 10505 5678
rect 10529 5676 10585 5678
rect 5622 5186 5678 5188
rect 5702 5186 5758 5188
rect 5782 5186 5838 5188
rect 5862 5186 5918 5188
rect 5622 5134 5648 5186
rect 5648 5134 5678 5186
rect 5702 5134 5712 5186
rect 5712 5134 5758 5186
rect 5782 5134 5828 5186
rect 5828 5134 5838 5186
rect 5862 5134 5892 5186
rect 5892 5134 5918 5186
rect 5622 5132 5678 5134
rect 5702 5132 5758 5134
rect 5782 5132 5838 5134
rect 5862 5132 5918 5134
rect 10289 4642 10345 4644
rect 10369 4642 10425 4644
rect 10449 4642 10505 4644
rect 10529 4642 10585 4644
rect 10289 4590 10315 4642
rect 10315 4590 10345 4642
rect 10369 4590 10379 4642
rect 10379 4590 10425 4642
rect 10449 4590 10495 4642
rect 10495 4590 10505 4642
rect 10529 4590 10559 4642
rect 10559 4590 10585 4642
rect 10289 4588 10345 4590
rect 10369 4588 10425 4590
rect 10449 4588 10505 4590
rect 10529 4588 10585 4590
rect 2870 4384 2926 4440
rect 5622 4098 5678 4100
rect 5702 4098 5758 4100
rect 5782 4098 5838 4100
rect 5862 4098 5918 4100
rect 5622 4046 5648 4098
rect 5648 4046 5678 4098
rect 5702 4046 5712 4098
rect 5712 4046 5758 4098
rect 5782 4046 5828 4098
rect 5828 4046 5838 4098
rect 5862 4046 5892 4098
rect 5892 4046 5918 4098
rect 5622 4044 5678 4046
rect 5702 4044 5758 4046
rect 5782 4044 5838 4046
rect 5862 4044 5918 4046
rect 10289 3554 10345 3556
rect 10369 3554 10425 3556
rect 10449 3554 10505 3556
rect 10529 3554 10585 3556
rect 10289 3502 10315 3554
rect 10315 3502 10345 3554
rect 10369 3502 10379 3554
rect 10379 3502 10425 3554
rect 10449 3502 10495 3554
rect 10495 3502 10505 3554
rect 10529 3502 10559 3554
rect 10559 3502 10585 3554
rect 10289 3500 10345 3502
rect 10369 3500 10425 3502
rect 10449 3500 10505 3502
rect 10529 3500 10585 3502
rect 5622 3010 5678 3012
rect 5702 3010 5758 3012
rect 5782 3010 5838 3012
rect 5862 3010 5918 3012
rect 5622 2958 5648 3010
rect 5648 2958 5678 3010
rect 5702 2958 5712 3010
rect 5712 2958 5758 3010
rect 5782 2958 5828 3010
rect 5828 2958 5838 3010
rect 5862 2958 5892 3010
rect 5892 2958 5918 3010
rect 5622 2956 5678 2958
rect 5702 2956 5758 2958
rect 5782 2956 5838 2958
rect 5862 2956 5918 2958
rect 10289 2466 10345 2468
rect 10369 2466 10425 2468
rect 10449 2466 10505 2468
rect 10529 2466 10585 2468
rect 10289 2414 10315 2466
rect 10315 2414 10345 2466
rect 10369 2414 10379 2466
rect 10379 2414 10425 2466
rect 10449 2414 10495 2466
rect 10495 2414 10505 2466
rect 10529 2414 10559 2466
rect 10559 2414 10585 2466
rect 10289 2412 10345 2414
rect 10369 2412 10425 2414
rect 10449 2412 10505 2414
rect 10529 2412 10585 2414
rect 5622 1922 5678 1924
rect 5702 1922 5758 1924
rect 5782 1922 5838 1924
rect 5862 1922 5918 1924
rect 5622 1870 5648 1922
rect 5648 1870 5678 1922
rect 5702 1870 5712 1922
rect 5712 1870 5758 1922
rect 5782 1870 5828 1922
rect 5828 1870 5838 1922
rect 5862 1870 5892 1922
rect 5892 1870 5918 1922
rect 5622 1868 5678 1870
rect 5702 1868 5758 1870
rect 5782 1868 5838 1870
rect 5862 1868 5918 1870
rect 14956 12802 15012 12804
rect 15036 12802 15092 12804
rect 15116 12802 15172 12804
rect 15196 12802 15252 12804
rect 14956 12750 14982 12802
rect 14982 12750 15012 12802
rect 15036 12750 15046 12802
rect 15046 12750 15092 12802
rect 15116 12750 15162 12802
rect 15162 12750 15172 12802
rect 15196 12750 15226 12802
rect 15226 12750 15252 12802
rect 14956 12748 15012 12750
rect 15036 12748 15092 12750
rect 15116 12748 15172 12750
rect 15196 12748 15252 12750
rect 13358 12444 13360 12464
rect 13360 12444 13412 12464
rect 13412 12444 13414 12464
rect 13358 12408 13414 12444
rect 14956 11714 15012 11716
rect 15036 11714 15092 11716
rect 15116 11714 15172 11716
rect 15196 11714 15252 11716
rect 14956 11662 14982 11714
rect 14982 11662 15012 11714
rect 15036 11662 15046 11714
rect 15046 11662 15092 11714
rect 15116 11662 15162 11714
rect 15162 11662 15172 11714
rect 15196 11662 15226 11714
rect 15226 11662 15252 11714
rect 14956 11660 15012 11662
rect 15036 11660 15092 11662
rect 15116 11660 15172 11662
rect 15196 11660 15252 11662
rect 14956 10626 15012 10628
rect 15036 10626 15092 10628
rect 15116 10626 15172 10628
rect 15196 10626 15252 10628
rect 14956 10574 14982 10626
rect 14982 10574 15012 10626
rect 15036 10574 15046 10626
rect 15046 10574 15092 10626
rect 15116 10574 15162 10626
rect 15162 10574 15172 10626
rect 15196 10574 15226 10626
rect 15226 10574 15252 10626
rect 14956 10572 15012 10574
rect 15036 10572 15092 10574
rect 15116 10572 15172 10574
rect 15196 10572 15252 10574
rect 14956 9538 15012 9540
rect 15036 9538 15092 9540
rect 15116 9538 15172 9540
rect 15196 9538 15252 9540
rect 14956 9486 14982 9538
rect 14982 9486 15012 9538
rect 15036 9486 15046 9538
rect 15046 9486 15092 9538
rect 15116 9486 15162 9538
rect 15162 9486 15172 9538
rect 15196 9486 15226 9538
rect 15226 9486 15252 9538
rect 14956 9484 15012 9486
rect 15036 9484 15092 9486
rect 15116 9484 15172 9486
rect 15196 9484 15252 9486
rect 14956 8450 15012 8452
rect 15036 8450 15092 8452
rect 15116 8450 15172 8452
rect 15196 8450 15252 8452
rect 14956 8398 14982 8450
rect 14982 8398 15012 8450
rect 15036 8398 15046 8450
rect 15046 8398 15092 8450
rect 15116 8398 15162 8450
rect 15162 8398 15172 8450
rect 15196 8398 15226 8450
rect 15226 8398 15252 8450
rect 14956 8396 15012 8398
rect 15036 8396 15092 8398
rect 15116 8396 15172 8398
rect 15196 8396 15252 8398
rect 14956 7362 15012 7364
rect 15036 7362 15092 7364
rect 15116 7362 15172 7364
rect 15196 7362 15252 7364
rect 14956 7310 14982 7362
rect 14982 7310 15012 7362
rect 15036 7310 15046 7362
rect 15046 7310 15092 7362
rect 15116 7310 15162 7362
rect 15162 7310 15172 7362
rect 15196 7310 15226 7362
rect 15226 7310 15252 7362
rect 14956 7308 15012 7310
rect 15036 7308 15092 7310
rect 15116 7308 15172 7310
rect 15196 7308 15252 7310
rect 14956 6274 15012 6276
rect 15036 6274 15092 6276
rect 15116 6274 15172 6276
rect 15196 6274 15252 6276
rect 14956 6222 14982 6274
rect 14982 6222 15012 6274
rect 15036 6222 15046 6274
rect 15046 6222 15092 6274
rect 15116 6222 15162 6274
rect 15162 6222 15172 6274
rect 15196 6222 15226 6274
rect 15226 6222 15252 6274
rect 14956 6220 15012 6222
rect 15036 6220 15092 6222
rect 15116 6220 15172 6222
rect 15196 6220 15252 6222
rect 14956 5186 15012 5188
rect 15036 5186 15092 5188
rect 15116 5186 15172 5188
rect 15196 5186 15252 5188
rect 14956 5134 14982 5186
rect 14982 5134 15012 5186
rect 15036 5134 15046 5186
rect 15046 5134 15092 5186
rect 15116 5134 15162 5186
rect 15162 5134 15172 5186
rect 15196 5134 15226 5186
rect 15226 5134 15252 5186
rect 14956 5132 15012 5134
rect 15036 5132 15092 5134
rect 15116 5132 15172 5134
rect 15196 5132 15252 5134
rect 14956 4098 15012 4100
rect 15036 4098 15092 4100
rect 15116 4098 15172 4100
rect 15196 4098 15252 4100
rect 14956 4046 14982 4098
rect 14982 4046 15012 4098
rect 15036 4046 15046 4098
rect 15046 4046 15092 4098
rect 15116 4046 15162 4098
rect 15162 4046 15172 4098
rect 15196 4046 15226 4098
rect 15226 4046 15252 4098
rect 14956 4044 15012 4046
rect 15036 4044 15092 4046
rect 15116 4044 15172 4046
rect 15196 4044 15252 4046
rect 14956 3010 15012 3012
rect 15036 3010 15092 3012
rect 15116 3010 15172 3012
rect 15196 3010 15252 3012
rect 14956 2958 14982 3010
rect 14982 2958 15012 3010
rect 15036 2958 15046 3010
rect 15046 2958 15092 3010
rect 15116 2958 15162 3010
rect 15162 2958 15172 3010
rect 15196 2958 15226 3010
rect 15226 2958 15252 3010
rect 14956 2956 15012 2958
rect 15036 2956 15092 2958
rect 15116 2956 15172 2958
rect 15196 2956 15252 2958
rect 14956 1922 15012 1924
rect 15036 1922 15092 1924
rect 15116 1922 15172 1924
rect 15196 1922 15252 1924
rect 14956 1870 14982 1922
rect 14982 1870 15012 1922
rect 15036 1870 15046 1922
rect 15046 1870 15092 1922
rect 15116 1870 15162 1922
rect 15162 1870 15172 1922
rect 15196 1870 15226 1922
rect 15226 1870 15252 1922
rect 14956 1868 15012 1870
rect 15036 1868 15092 1870
rect 15116 1868 15172 1870
rect 15196 1868 15252 1870
rect 15934 12444 15936 12464
rect 15936 12444 15988 12464
rect 15988 12444 15990 12464
rect 15934 12408 15990 12444
rect 17866 23832 17922 23888
rect 16854 22236 16856 22256
rect 16856 22236 16908 22256
rect 16908 22236 16910 22256
rect 16854 22200 16910 22236
rect 16762 19752 16818 19808
rect 16762 19344 16818 19400
rect 18510 22336 18566 22392
rect 18234 21792 18290 21848
rect 18142 21404 18198 21440
rect 18142 21384 18144 21404
rect 18144 21384 18196 21404
rect 18196 21384 18198 21404
rect 18326 18936 18382 18992
rect 18786 18970 18842 19026
rect 18142 18256 18198 18312
rect 18234 17476 18236 17496
rect 18236 17476 18288 17496
rect 18288 17476 18290 17496
rect 18234 17440 18290 17476
rect 18234 12952 18290 13008
rect 18510 12408 18566 12464
rect 19622 25314 19678 25316
rect 19702 25314 19758 25316
rect 19782 25314 19838 25316
rect 19862 25314 19918 25316
rect 19622 25262 19648 25314
rect 19648 25262 19678 25314
rect 19702 25262 19712 25314
rect 19712 25262 19758 25314
rect 19782 25262 19828 25314
rect 19828 25262 19838 25314
rect 19862 25262 19892 25314
rect 19892 25262 19918 25314
rect 19622 25260 19678 25262
rect 19702 25260 19758 25262
rect 19782 25260 19838 25262
rect 19862 25260 19918 25262
rect 19622 24226 19678 24228
rect 19702 24226 19758 24228
rect 19782 24226 19838 24228
rect 19862 24226 19918 24228
rect 19622 24174 19648 24226
rect 19648 24174 19678 24226
rect 19702 24174 19712 24226
rect 19712 24174 19758 24226
rect 19782 24174 19828 24226
rect 19828 24174 19838 24226
rect 19862 24174 19892 24226
rect 19892 24174 19918 24226
rect 19622 24172 19678 24174
rect 19702 24172 19758 24174
rect 19782 24172 19838 24174
rect 19862 24172 19918 24174
rect 19890 23832 19946 23888
rect 19062 23308 19118 23344
rect 19062 23288 19064 23308
rect 19064 23288 19116 23308
rect 19116 23288 19118 23308
rect 19622 23138 19678 23140
rect 19702 23138 19758 23140
rect 19782 23138 19838 23140
rect 19862 23138 19918 23140
rect 19622 23086 19648 23138
rect 19648 23086 19678 23138
rect 19702 23086 19712 23138
rect 19712 23086 19758 23138
rect 19782 23086 19828 23138
rect 19828 23086 19838 23138
rect 19862 23086 19892 23138
rect 19892 23086 19918 23138
rect 19622 23084 19678 23086
rect 19702 23084 19758 23086
rect 19782 23084 19838 23086
rect 19862 23084 19918 23086
rect 19622 22050 19678 22052
rect 19702 22050 19758 22052
rect 19782 22050 19838 22052
rect 19862 22050 19918 22052
rect 19622 21998 19648 22050
rect 19648 21998 19678 22050
rect 19702 21998 19712 22050
rect 19712 21998 19758 22050
rect 19782 21998 19828 22050
rect 19828 21998 19838 22050
rect 19862 21998 19892 22050
rect 19892 21998 19918 22050
rect 19622 21996 19678 21998
rect 19702 21996 19758 21998
rect 19782 21996 19838 21998
rect 19862 21996 19918 21998
rect 19430 21384 19486 21440
rect 19062 20160 19118 20216
rect 19622 20962 19678 20964
rect 19702 20962 19758 20964
rect 19782 20962 19838 20964
rect 19862 20962 19918 20964
rect 19622 20910 19648 20962
rect 19648 20910 19678 20962
rect 19702 20910 19712 20962
rect 19712 20910 19758 20962
rect 19782 20910 19828 20962
rect 19828 20910 19838 20962
rect 19862 20910 19892 20962
rect 19892 20910 19918 20962
rect 19622 20908 19678 20910
rect 19702 20908 19758 20910
rect 19782 20908 19838 20910
rect 19862 20908 19918 20910
rect 19798 20316 19854 20352
rect 19798 20296 19800 20316
rect 19800 20296 19852 20316
rect 19852 20296 19854 20316
rect 19622 19874 19678 19876
rect 19702 19874 19758 19876
rect 19782 19874 19838 19876
rect 19862 19874 19918 19876
rect 19622 19822 19648 19874
rect 19648 19822 19678 19874
rect 19702 19822 19712 19874
rect 19712 19822 19758 19874
rect 19782 19822 19828 19874
rect 19828 19822 19838 19874
rect 19862 19822 19892 19874
rect 19892 19822 19918 19874
rect 19622 19820 19678 19822
rect 19702 19820 19758 19822
rect 19782 19820 19838 19822
rect 19862 19820 19918 19822
rect 18970 18528 19026 18584
rect 19338 18684 19394 18720
rect 19338 18664 19340 18684
rect 19340 18664 19392 18684
rect 19392 18664 19394 18684
rect 19622 18786 19678 18788
rect 19702 18786 19758 18788
rect 19782 18786 19838 18788
rect 19862 18786 19918 18788
rect 19622 18734 19648 18786
rect 19648 18734 19678 18786
rect 19702 18734 19712 18786
rect 19712 18734 19758 18786
rect 19782 18734 19828 18786
rect 19828 18734 19838 18786
rect 19862 18734 19892 18786
rect 19892 18734 19918 18786
rect 19622 18732 19678 18734
rect 19702 18732 19758 18734
rect 19782 18732 19838 18734
rect 19862 18732 19918 18734
rect 20166 18836 20168 18856
rect 20168 18836 20220 18856
rect 20220 18836 20222 18856
rect 20166 18800 20222 18836
rect 19246 17848 19302 17904
rect 19622 17698 19678 17700
rect 19702 17698 19758 17700
rect 19782 17698 19838 17700
rect 19862 17698 19918 17700
rect 19622 17646 19648 17698
rect 19648 17646 19678 17698
rect 19702 17646 19712 17698
rect 19712 17646 19758 17698
rect 19782 17646 19828 17698
rect 19828 17646 19838 17698
rect 19862 17646 19892 17698
rect 19892 17646 19918 17698
rect 19622 17644 19678 17646
rect 19702 17644 19758 17646
rect 19782 17644 19838 17646
rect 19862 17644 19918 17646
rect 19622 16610 19678 16612
rect 19702 16610 19758 16612
rect 19782 16610 19838 16612
rect 19862 16610 19918 16612
rect 19622 16558 19648 16610
rect 19648 16558 19678 16610
rect 19702 16558 19712 16610
rect 19712 16558 19758 16610
rect 19782 16558 19828 16610
rect 19828 16558 19838 16610
rect 19862 16558 19892 16610
rect 19892 16558 19918 16610
rect 19622 16556 19678 16558
rect 19702 16556 19758 16558
rect 19782 16556 19838 16558
rect 19862 16556 19918 16558
rect 19622 15522 19678 15524
rect 19702 15522 19758 15524
rect 19782 15522 19838 15524
rect 19862 15522 19918 15524
rect 19622 15470 19648 15522
rect 19648 15470 19678 15522
rect 19702 15470 19712 15522
rect 19712 15470 19758 15522
rect 19782 15470 19828 15522
rect 19828 15470 19838 15522
rect 19862 15470 19892 15522
rect 19892 15470 19918 15522
rect 19622 15468 19678 15470
rect 19702 15468 19758 15470
rect 19782 15468 19838 15470
rect 19862 15468 19918 15470
rect 19622 14434 19678 14436
rect 19702 14434 19758 14436
rect 19782 14434 19838 14436
rect 19862 14434 19918 14436
rect 19622 14382 19648 14434
rect 19648 14382 19678 14434
rect 19702 14382 19712 14434
rect 19712 14382 19758 14434
rect 19782 14382 19828 14434
rect 19828 14382 19838 14434
rect 19862 14382 19892 14434
rect 19892 14382 19918 14434
rect 19622 14380 19678 14382
rect 19702 14380 19758 14382
rect 19782 14380 19838 14382
rect 19862 14380 19918 14382
rect 19622 13346 19678 13348
rect 19702 13346 19758 13348
rect 19782 13346 19838 13348
rect 19862 13346 19918 13348
rect 19622 13294 19648 13346
rect 19648 13294 19678 13346
rect 19702 13294 19712 13346
rect 19712 13294 19758 13346
rect 19782 13294 19828 13346
rect 19828 13294 19838 13346
rect 19862 13294 19892 13346
rect 19892 13294 19918 13346
rect 19622 13292 19678 13294
rect 19702 13292 19758 13294
rect 19782 13292 19838 13294
rect 19862 13292 19918 13294
rect 18878 12272 18934 12328
rect 18878 12000 18934 12056
rect 18326 5336 18382 5392
rect 19622 12258 19678 12260
rect 19702 12258 19758 12260
rect 19782 12258 19838 12260
rect 19862 12258 19918 12260
rect 19622 12206 19648 12258
rect 19648 12206 19678 12258
rect 19702 12206 19712 12258
rect 19712 12206 19758 12258
rect 19782 12206 19828 12258
rect 19828 12206 19838 12258
rect 19862 12206 19892 12258
rect 19892 12206 19918 12258
rect 19622 12204 19678 12206
rect 19702 12204 19758 12206
rect 19782 12204 19838 12206
rect 19862 12204 19918 12206
rect 19622 11170 19678 11172
rect 19702 11170 19758 11172
rect 19782 11170 19838 11172
rect 19862 11170 19918 11172
rect 19622 11118 19648 11170
rect 19648 11118 19678 11170
rect 19702 11118 19712 11170
rect 19712 11118 19758 11170
rect 19782 11118 19828 11170
rect 19828 11118 19838 11170
rect 19862 11118 19892 11170
rect 19892 11118 19918 11170
rect 19622 11116 19678 11118
rect 19702 11116 19758 11118
rect 19782 11116 19838 11118
rect 19862 11116 19918 11118
rect 19622 10082 19678 10084
rect 19702 10082 19758 10084
rect 19782 10082 19838 10084
rect 19862 10082 19918 10084
rect 19622 10030 19648 10082
rect 19648 10030 19678 10082
rect 19702 10030 19712 10082
rect 19712 10030 19758 10082
rect 19782 10030 19828 10082
rect 19828 10030 19838 10082
rect 19862 10030 19892 10082
rect 19892 10030 19918 10082
rect 19622 10028 19678 10030
rect 19702 10028 19758 10030
rect 19782 10028 19838 10030
rect 19862 10028 19918 10030
rect 19622 8994 19678 8996
rect 19702 8994 19758 8996
rect 19782 8994 19838 8996
rect 19862 8994 19918 8996
rect 19622 8942 19648 8994
rect 19648 8942 19678 8994
rect 19702 8942 19712 8994
rect 19712 8942 19758 8994
rect 19782 8942 19828 8994
rect 19828 8942 19838 8994
rect 19862 8942 19892 8994
rect 19892 8942 19918 8994
rect 19622 8940 19678 8942
rect 19702 8940 19758 8942
rect 19782 8940 19838 8942
rect 19862 8940 19918 8942
rect 19622 7906 19678 7908
rect 19702 7906 19758 7908
rect 19782 7906 19838 7908
rect 19862 7906 19918 7908
rect 19622 7854 19648 7906
rect 19648 7854 19678 7906
rect 19702 7854 19712 7906
rect 19712 7854 19758 7906
rect 19782 7854 19828 7906
rect 19828 7854 19838 7906
rect 19862 7854 19892 7906
rect 19892 7854 19918 7906
rect 19622 7852 19678 7854
rect 19702 7852 19758 7854
rect 19782 7852 19838 7854
rect 19862 7852 19918 7854
rect 19622 6818 19678 6820
rect 19702 6818 19758 6820
rect 19782 6818 19838 6820
rect 19862 6818 19918 6820
rect 19622 6766 19648 6818
rect 19648 6766 19678 6818
rect 19702 6766 19712 6818
rect 19712 6766 19758 6818
rect 19782 6766 19828 6818
rect 19828 6766 19838 6818
rect 19862 6766 19892 6818
rect 19892 6766 19918 6818
rect 19622 6764 19678 6766
rect 19702 6764 19758 6766
rect 19782 6764 19838 6766
rect 19862 6764 19918 6766
rect 20350 6424 20406 6480
rect 20074 5780 20076 5800
rect 20076 5780 20128 5800
rect 20128 5780 20130 5800
rect 20074 5744 20130 5780
rect 19622 5730 19678 5732
rect 19702 5730 19758 5732
rect 19782 5730 19838 5732
rect 19862 5730 19918 5732
rect 19622 5678 19648 5730
rect 19648 5678 19678 5730
rect 19702 5678 19712 5730
rect 19712 5678 19758 5730
rect 19782 5678 19828 5730
rect 19828 5678 19838 5730
rect 19862 5678 19892 5730
rect 19892 5678 19918 5730
rect 19622 5676 19678 5678
rect 19702 5676 19758 5678
rect 19782 5676 19838 5678
rect 19862 5676 19918 5678
rect 20534 22200 20590 22256
rect 20718 21404 20774 21440
rect 20718 21384 20720 21404
rect 20720 21384 20772 21404
rect 20772 21384 20774 21404
rect 20534 18428 20536 18448
rect 20536 18428 20588 18448
rect 20588 18428 20590 18448
rect 20534 18392 20590 18428
rect 20534 17748 20536 17768
rect 20536 17748 20588 17768
rect 20588 17748 20590 17768
rect 20534 17712 20590 17748
rect 20718 16796 20720 16816
rect 20720 16796 20772 16816
rect 20772 16796 20774 16816
rect 20718 16760 20774 16796
rect 21086 16352 21142 16408
rect 21362 20860 21418 20896
rect 21362 20840 21364 20860
rect 21364 20840 21416 20860
rect 21416 20840 21418 20860
rect 23202 24396 23258 24432
rect 23202 24376 23204 24396
rect 23204 24376 23256 24396
rect 23256 24376 23258 24396
rect 23202 23424 23258 23480
rect 22742 22336 22798 22392
rect 22650 19344 22706 19400
rect 23754 26280 23810 26336
rect 23478 20044 23534 20080
rect 23478 20024 23480 20044
rect 23480 20024 23532 20044
rect 23532 20024 23534 20044
rect 23202 18800 23258 18856
rect 21730 18120 21786 18176
rect 21822 17848 21878 17904
rect 21638 16488 21694 16544
rect 22190 17868 22246 17904
rect 22190 17848 22192 17868
rect 22192 17848 22244 17868
rect 22244 17848 22246 17868
rect 22926 14604 22982 14640
rect 22926 14584 22928 14604
rect 22928 14584 22980 14604
rect 22980 14584 22982 14604
rect 22282 12408 22338 12464
rect 22006 11728 22062 11784
rect 23662 18392 23718 18448
rect 23662 16760 23718 16816
rect 23570 14992 23626 15048
rect 23846 20160 23902 20216
rect 24030 20316 24086 20352
rect 24030 20296 24032 20316
rect 24032 20296 24084 20316
rect 24084 20296 24086 20316
rect 23938 18120 23994 18176
rect 23846 17712 23902 17768
rect 21638 6868 21640 6888
rect 21640 6868 21692 6888
rect 21692 6868 21694 6888
rect 21638 6832 21694 6868
rect 20442 5064 20498 5120
rect 23478 5084 23534 5120
rect 23478 5064 23480 5084
rect 23480 5064 23532 5084
rect 23532 5064 23534 5084
rect 19062 4792 19118 4848
rect 19622 4642 19678 4644
rect 19702 4642 19758 4644
rect 19782 4642 19838 4644
rect 19862 4642 19918 4644
rect 19622 4590 19648 4642
rect 19648 4590 19678 4642
rect 19702 4590 19712 4642
rect 19712 4590 19758 4642
rect 19782 4590 19828 4642
rect 19828 4590 19838 4642
rect 19862 4590 19892 4642
rect 19892 4590 19918 4642
rect 19622 4588 19678 4590
rect 19702 4588 19758 4590
rect 19782 4588 19838 4590
rect 19862 4588 19918 4590
rect 18878 3704 18934 3760
rect 19622 3554 19678 3556
rect 19702 3554 19758 3556
rect 19782 3554 19838 3556
rect 19862 3554 19918 3556
rect 19622 3502 19648 3554
rect 19648 3502 19678 3554
rect 19702 3502 19712 3554
rect 19712 3502 19758 3554
rect 19782 3502 19828 3554
rect 19828 3502 19838 3554
rect 19862 3502 19892 3554
rect 19892 3502 19918 3554
rect 19622 3500 19678 3502
rect 19702 3500 19758 3502
rect 19782 3500 19838 3502
rect 19862 3500 19918 3502
rect 16762 2772 16818 2808
rect 16762 2752 16764 2772
rect 16764 2752 16816 2772
rect 16816 2752 16818 2772
rect 19622 2466 19678 2468
rect 19702 2466 19758 2468
rect 19782 2466 19838 2468
rect 19862 2466 19918 2468
rect 19622 2414 19648 2466
rect 19648 2414 19678 2466
rect 19702 2414 19712 2466
rect 19712 2414 19758 2466
rect 19782 2414 19828 2466
rect 19828 2414 19838 2466
rect 19862 2414 19892 2466
rect 19892 2414 19918 2466
rect 19622 2412 19678 2414
rect 19702 2412 19758 2414
rect 19782 2412 19838 2414
rect 19862 2412 19918 2414
rect 16670 2072 16726 2128
rect 15842 1256 15898 1312
rect 13266 1120 13322 1176
rect 23662 13088 23718 13144
rect 23662 11728 23718 11784
rect 24766 26824 24822 26880
rect 24766 25736 24822 25792
rect 24674 25056 24730 25112
rect 24289 24770 24345 24772
rect 24369 24770 24425 24772
rect 24449 24770 24505 24772
rect 24529 24770 24585 24772
rect 24289 24718 24315 24770
rect 24315 24718 24345 24770
rect 24369 24718 24379 24770
rect 24379 24718 24425 24770
rect 24449 24718 24495 24770
rect 24495 24718 24505 24770
rect 24529 24718 24559 24770
rect 24559 24718 24585 24770
rect 24289 24716 24345 24718
rect 24369 24716 24425 24718
rect 24449 24716 24505 24718
rect 24529 24716 24585 24718
rect 24950 24512 25006 24568
rect 24674 23868 24676 23888
rect 24676 23868 24728 23888
rect 24728 23868 24730 23888
rect 24674 23832 24730 23868
rect 24289 23682 24345 23684
rect 24369 23682 24425 23684
rect 24449 23682 24505 23684
rect 24529 23682 24585 23684
rect 24289 23630 24315 23682
rect 24315 23630 24345 23682
rect 24369 23630 24379 23682
rect 24379 23630 24425 23682
rect 24449 23630 24495 23682
rect 24495 23630 24505 23682
rect 24529 23630 24559 23682
rect 24559 23630 24585 23682
rect 24289 23628 24345 23630
rect 24369 23628 24425 23630
rect 24449 23628 24505 23630
rect 24529 23628 24585 23630
rect 24289 22594 24345 22596
rect 24369 22594 24425 22596
rect 24449 22594 24505 22596
rect 24529 22594 24585 22596
rect 24289 22542 24315 22594
rect 24315 22542 24345 22594
rect 24369 22542 24379 22594
rect 24379 22542 24425 22594
rect 24449 22542 24495 22594
rect 24495 22542 24505 22594
rect 24529 22542 24559 22594
rect 24559 22542 24585 22594
rect 24289 22540 24345 22542
rect 24369 22540 24425 22542
rect 24449 22540 24505 22542
rect 24529 22540 24585 22542
rect 25686 24512 25742 24568
rect 25502 23968 25558 24024
rect 25134 22880 25190 22936
rect 25042 22336 25098 22392
rect 24582 21792 24638 21848
rect 24289 21506 24345 21508
rect 24369 21506 24425 21508
rect 24449 21506 24505 21508
rect 24529 21506 24585 21508
rect 24289 21454 24315 21506
rect 24315 21454 24345 21506
rect 24369 21454 24379 21506
rect 24379 21454 24425 21506
rect 24449 21454 24495 21506
rect 24495 21454 24505 21506
rect 24529 21454 24559 21506
rect 24559 21454 24585 21506
rect 24289 21452 24345 21454
rect 24369 21452 24425 21454
rect 24449 21452 24505 21454
rect 24529 21452 24585 21454
rect 24766 21656 24822 21712
rect 24766 21112 24822 21168
rect 24289 20418 24345 20420
rect 24369 20418 24425 20420
rect 24449 20418 24505 20420
rect 24529 20418 24585 20420
rect 24289 20366 24315 20418
rect 24315 20366 24345 20418
rect 24369 20366 24379 20418
rect 24379 20366 24425 20418
rect 24449 20366 24495 20418
rect 24495 20366 24505 20418
rect 24529 20366 24559 20418
rect 24559 20366 24585 20418
rect 24289 20364 24345 20366
rect 24369 20364 24425 20366
rect 24449 20364 24505 20366
rect 24529 20364 24585 20366
rect 24289 19330 24345 19332
rect 24369 19330 24425 19332
rect 24449 19330 24505 19332
rect 24529 19330 24585 19332
rect 24289 19278 24315 19330
rect 24315 19278 24345 19330
rect 24369 19278 24379 19330
rect 24379 19278 24425 19330
rect 24449 19278 24495 19330
rect 24495 19278 24505 19330
rect 24529 19278 24559 19330
rect 24559 19278 24585 19330
rect 24289 19276 24345 19278
rect 24369 19276 24425 19278
rect 24449 19276 24505 19278
rect 24529 19276 24585 19278
rect 24214 18392 24270 18448
rect 24289 18242 24345 18244
rect 24369 18242 24425 18244
rect 24449 18242 24505 18244
rect 24529 18242 24585 18244
rect 24289 18190 24315 18242
rect 24315 18190 24345 18242
rect 24369 18190 24379 18242
rect 24379 18190 24425 18242
rect 24449 18190 24495 18242
rect 24495 18190 24505 18242
rect 24529 18190 24559 18242
rect 24559 18190 24585 18242
rect 24289 18188 24345 18190
rect 24369 18188 24425 18190
rect 24449 18188 24505 18190
rect 24529 18188 24585 18190
rect 23938 16488 23994 16544
rect 24289 17154 24345 17156
rect 24369 17154 24425 17156
rect 24449 17154 24505 17156
rect 24529 17154 24585 17156
rect 24289 17102 24315 17154
rect 24315 17102 24345 17154
rect 24369 17102 24379 17154
rect 24379 17102 24425 17154
rect 24449 17102 24495 17154
rect 24495 17102 24505 17154
rect 24529 17102 24559 17154
rect 24559 17102 24585 17154
rect 24289 17100 24345 17102
rect 24369 17100 24425 17102
rect 24449 17100 24505 17102
rect 24529 17100 24585 17102
rect 24214 16488 24270 16544
rect 24122 14992 24178 15048
rect 24289 16066 24345 16068
rect 24369 16066 24425 16068
rect 24449 16066 24505 16068
rect 24529 16066 24585 16068
rect 24289 16014 24315 16066
rect 24315 16014 24345 16066
rect 24369 16014 24379 16066
rect 24379 16014 24425 16066
rect 24449 16014 24495 16066
rect 24495 16014 24505 16066
rect 24529 16014 24559 16066
rect 24559 16014 24585 16066
rect 24289 16012 24345 16014
rect 24369 16012 24425 16014
rect 24449 16012 24505 16014
rect 24529 16012 24585 16014
rect 25318 20724 25374 20760
rect 25318 20704 25320 20724
rect 25320 20704 25372 20724
rect 25372 20704 25374 20724
rect 25134 19616 25190 19672
rect 25410 19344 25466 19400
rect 25318 18836 25320 18856
rect 25320 18836 25372 18856
rect 25372 18836 25374 18856
rect 25318 18800 25374 18836
rect 24766 17712 24822 17768
rect 25410 17168 25466 17224
rect 25134 16896 25190 16952
rect 25042 16760 25098 16816
rect 24289 14978 24345 14980
rect 24369 14978 24425 14980
rect 24449 14978 24505 14980
rect 24529 14978 24585 14980
rect 24289 14926 24315 14978
rect 24315 14926 24345 14978
rect 24369 14926 24379 14978
rect 24379 14926 24425 14978
rect 24449 14926 24495 14978
rect 24495 14926 24505 14978
rect 24529 14926 24559 14978
rect 24559 14926 24585 14978
rect 24289 14924 24345 14926
rect 24369 14924 24425 14926
rect 24449 14924 24505 14926
rect 24529 14924 24585 14926
rect 24674 14876 24730 14912
rect 24674 14856 24676 14876
rect 24676 14856 24728 14876
rect 24728 14856 24730 14876
rect 25226 16372 25282 16408
rect 25226 16352 25228 16372
rect 25228 16352 25280 16372
rect 25280 16352 25282 16372
rect 25410 15944 25466 16000
rect 25410 15420 25466 15456
rect 25410 15400 25412 15420
rect 25412 15400 25464 15420
rect 25464 15400 25466 15420
rect 24858 14312 24914 14368
rect 24289 13890 24345 13892
rect 24369 13890 24425 13892
rect 24449 13890 24505 13892
rect 24529 13890 24585 13892
rect 24289 13838 24315 13890
rect 24315 13838 24345 13890
rect 24369 13838 24379 13890
rect 24379 13838 24425 13890
rect 24449 13838 24495 13890
rect 24495 13838 24505 13890
rect 24529 13838 24559 13890
rect 24559 13838 24585 13890
rect 24289 13836 24345 13838
rect 24369 13836 24425 13838
rect 24449 13836 24505 13838
rect 24529 13836 24585 13838
rect 24582 13632 24638 13688
rect 24766 13632 24822 13688
rect 24582 12952 24638 13008
rect 24289 12802 24345 12804
rect 24369 12802 24425 12804
rect 24449 12802 24505 12804
rect 24529 12802 24585 12804
rect 24289 12750 24315 12802
rect 24315 12750 24345 12802
rect 24369 12750 24379 12802
rect 24379 12750 24425 12802
rect 24449 12750 24495 12802
rect 24495 12750 24505 12802
rect 24529 12750 24559 12802
rect 24559 12750 24585 12802
rect 24289 12748 24345 12750
rect 24369 12748 24425 12750
rect 24449 12748 24505 12750
rect 24529 12748 24585 12750
rect 24766 12580 24768 12600
rect 24768 12580 24820 12600
rect 24820 12580 24822 12600
rect 24766 12544 24822 12580
rect 24766 12000 24822 12056
rect 24289 11714 24345 11716
rect 24369 11714 24425 11716
rect 24449 11714 24505 11716
rect 24529 11714 24585 11716
rect 24289 11662 24315 11714
rect 24315 11662 24345 11714
rect 24369 11662 24379 11714
rect 24379 11662 24425 11714
rect 24449 11662 24495 11714
rect 24495 11662 24505 11714
rect 24529 11662 24559 11714
rect 24559 11662 24585 11714
rect 24289 11660 24345 11662
rect 24369 11660 24425 11662
rect 24449 11660 24505 11662
rect 24529 11660 24585 11662
rect 24766 11612 24822 11648
rect 24766 11592 24768 11612
rect 24768 11592 24820 11612
rect 24820 11592 24822 11612
rect 25226 11476 25282 11512
rect 25226 11456 25228 11476
rect 25228 11456 25280 11476
rect 25280 11456 25282 11476
rect 24582 10776 24638 10832
rect 24289 10626 24345 10628
rect 24369 10626 24425 10628
rect 24449 10626 24505 10628
rect 24529 10626 24585 10628
rect 24289 10574 24315 10626
rect 24315 10574 24345 10626
rect 24369 10574 24379 10626
rect 24379 10574 24425 10626
rect 24449 10574 24495 10626
rect 24495 10574 24505 10626
rect 24529 10574 24559 10626
rect 24559 10574 24585 10626
rect 24289 10572 24345 10574
rect 24369 10572 24425 10574
rect 24449 10572 24505 10574
rect 24529 10572 24585 10574
rect 24766 10524 24822 10560
rect 24766 10504 24768 10524
rect 24768 10504 24820 10524
rect 24820 10504 24822 10524
rect 25594 10504 25650 10560
rect 25226 10252 25282 10288
rect 25226 10232 25228 10252
rect 25228 10232 25280 10252
rect 25280 10232 25282 10252
rect 24582 9688 24638 9744
rect 24289 9538 24345 9540
rect 24369 9538 24425 9540
rect 24449 9538 24505 9540
rect 24529 9538 24585 9540
rect 24289 9486 24315 9538
rect 24315 9486 24345 9538
rect 24369 9486 24379 9538
rect 24379 9486 24425 9538
rect 24449 9486 24495 9538
rect 24495 9486 24505 9538
rect 24529 9486 24559 9538
rect 24559 9486 24585 9538
rect 24289 9484 24345 9486
rect 24369 9484 24425 9486
rect 24449 9484 24505 9486
rect 24529 9484 24585 9486
rect 24398 9164 24454 9200
rect 24398 9144 24400 9164
rect 24400 9144 24452 9164
rect 24452 9144 24454 9164
rect 24398 8600 24454 8656
rect 24674 8600 24730 8656
rect 24289 8450 24345 8452
rect 24369 8450 24425 8452
rect 24449 8450 24505 8452
rect 24529 8450 24585 8452
rect 24289 8398 24315 8450
rect 24315 8398 24345 8450
rect 24369 8398 24379 8450
rect 24379 8398 24425 8450
rect 24449 8398 24495 8450
rect 24495 8398 24505 8450
rect 24529 8398 24559 8450
rect 24559 8398 24585 8450
rect 24289 8396 24345 8398
rect 24369 8396 24425 8398
rect 24449 8396 24505 8398
rect 24529 8396 24585 8398
rect 23662 7920 23718 7976
rect 24674 7376 24730 7432
rect 24289 7362 24345 7364
rect 24369 7362 24425 7364
rect 24449 7362 24505 7364
rect 24529 7362 24585 7364
rect 24289 7310 24315 7362
rect 24315 7310 24345 7362
rect 24369 7310 24379 7362
rect 24379 7310 24425 7362
rect 24449 7310 24495 7362
rect 24495 7310 24505 7362
rect 24529 7310 24559 7362
rect 24559 7310 24585 7362
rect 24289 7308 24345 7310
rect 24369 7308 24425 7310
rect 24449 7308 24505 7310
rect 24529 7308 24585 7310
rect 24289 6274 24345 6276
rect 24369 6274 24425 6276
rect 24449 6274 24505 6276
rect 24529 6274 24585 6276
rect 24289 6222 24315 6274
rect 24315 6222 24345 6274
rect 24369 6222 24379 6274
rect 24379 6222 24425 6274
rect 24449 6222 24495 6274
rect 24495 6222 24505 6274
rect 24529 6222 24559 6274
rect 24559 6222 24585 6274
rect 24289 6220 24345 6222
rect 24369 6220 24425 6222
rect 24449 6220 24505 6222
rect 24529 6220 24585 6222
rect 23938 5336 23994 5392
rect 24289 5186 24345 5188
rect 24369 5186 24425 5188
rect 24449 5186 24505 5188
rect 24529 5186 24585 5188
rect 24289 5134 24315 5186
rect 24315 5134 24345 5186
rect 24369 5134 24379 5186
rect 24379 5134 24425 5186
rect 24449 5134 24495 5186
rect 24495 5134 24505 5186
rect 24529 5134 24559 5186
rect 24559 5134 24585 5186
rect 24289 5132 24345 5134
rect 24369 5132 24425 5134
rect 24449 5132 24505 5134
rect 24529 5132 24585 5134
rect 25226 5084 25282 5120
rect 25226 5064 25228 5084
rect 25228 5064 25280 5084
rect 25280 5064 25282 5084
rect 24766 4792 24822 4848
rect 24582 4520 24638 4576
rect 24289 4098 24345 4100
rect 24369 4098 24425 4100
rect 24449 4098 24505 4100
rect 24529 4098 24585 4100
rect 24289 4046 24315 4098
rect 24315 4046 24345 4098
rect 24369 4046 24379 4098
rect 24379 4046 24425 4098
rect 24449 4046 24495 4098
rect 24495 4046 24505 4098
rect 24529 4046 24559 4098
rect 24559 4046 24585 4098
rect 24289 4044 24345 4046
rect 24369 4044 24425 4046
rect 24449 4044 24505 4046
rect 24529 4044 24585 4046
rect 25226 3976 25282 4032
rect 24766 3704 24822 3760
rect 23938 3432 23994 3488
rect 26882 11592 26938 11648
rect 24766 3024 24822 3080
rect 26238 3024 26294 3080
rect 24289 3010 24345 3012
rect 24369 3010 24425 3012
rect 24449 3010 24505 3012
rect 24529 3010 24585 3012
rect 24289 2958 24315 3010
rect 24315 2958 24345 3010
rect 24369 2958 24379 3010
rect 24379 2958 24425 3010
rect 24449 2958 24495 3010
rect 24495 2958 24505 3010
rect 24529 2958 24559 3010
rect 24559 2958 24585 3010
rect 24289 2956 24345 2958
rect 24369 2956 24425 2958
rect 24449 2956 24505 2958
rect 24529 2956 24585 2958
rect 24289 1922 24345 1924
rect 24369 1922 24425 1924
rect 24449 1922 24505 1924
rect 24529 1922 24585 1924
rect 24289 1870 24315 1922
rect 24315 1870 24345 1922
rect 24369 1870 24379 1922
rect 24379 1870 24425 1922
rect 24449 1870 24495 1922
rect 24495 1870 24505 1922
rect 24529 1870 24559 1922
rect 24559 1870 24585 1922
rect 24289 1868 24345 1870
rect 24369 1868 24425 1870
rect 24449 1868 24505 1870
rect 24529 1868 24585 1870
rect 24766 2092 24822 2128
rect 24766 2072 24768 2092
rect 24768 2072 24820 2092
rect 24820 2072 24822 2092
rect 25226 1664 25282 1720
rect 24674 576 24730 632
rect 23570 32 23626 88
<< metal3 >>
rect 25865 27426 25931 27429
rect 27520 27426 28000 27456
rect 25865 27424 28000 27426
rect 25865 27368 25870 27424
rect 25926 27368 28000 27424
rect 25865 27366 28000 27368
rect 25865 27363 25931 27366
rect 27520 27336 28000 27366
rect 24761 26882 24827 26885
rect 27520 26882 28000 26912
rect 24761 26880 28000 26882
rect 24761 26824 24766 26880
rect 24822 26824 28000 26880
rect 24761 26822 28000 26824
rect 24761 26819 24827 26822
rect 27520 26792 28000 26822
rect 23749 26338 23815 26341
rect 27520 26338 28000 26368
rect 23749 26336 28000 26338
rect 23749 26280 23754 26336
rect 23810 26280 28000 26336
rect 23749 26278 28000 26280
rect 23749 26275 23815 26278
rect 27520 26248 28000 26278
rect 24761 25794 24827 25797
rect 27520 25794 28000 25824
rect 24761 25792 28000 25794
rect 24761 25736 24766 25792
rect 24822 25736 28000 25792
rect 24761 25734 28000 25736
rect 24761 25731 24827 25734
rect 27520 25704 28000 25734
rect 10277 25320 10597 25321
rect 10277 25256 10285 25320
rect 10349 25256 10365 25320
rect 10429 25256 10445 25320
rect 10509 25256 10525 25320
rect 10589 25256 10597 25320
rect 10277 25255 10597 25256
rect 19610 25320 19930 25321
rect 19610 25256 19618 25320
rect 19682 25256 19698 25320
rect 19762 25256 19778 25320
rect 19842 25256 19858 25320
rect 19922 25256 19930 25320
rect 19610 25255 19930 25256
rect 24669 25114 24735 25117
rect 27520 25114 28000 25144
rect 24669 25112 28000 25114
rect 24669 25056 24674 25112
rect 24730 25056 28000 25112
rect 24669 25054 28000 25056
rect 24669 25051 24735 25054
rect 27520 25024 28000 25054
rect 5610 24776 5930 24777
rect 5610 24712 5618 24776
rect 5682 24712 5698 24776
rect 5762 24712 5778 24776
rect 5842 24712 5858 24776
rect 5922 24712 5930 24776
rect 5610 24711 5930 24712
rect 14944 24776 15264 24777
rect 14944 24712 14952 24776
rect 15016 24712 15032 24776
rect 15096 24712 15112 24776
rect 15176 24712 15192 24776
rect 15256 24712 15264 24776
rect 14944 24711 15264 24712
rect 24277 24776 24597 24777
rect 24277 24712 24285 24776
rect 24349 24712 24365 24776
rect 24429 24712 24445 24776
rect 24509 24712 24525 24776
rect 24589 24712 24597 24776
rect 24277 24711 24597 24712
rect 13169 24570 13235 24573
rect 24945 24570 25011 24573
rect 13169 24568 25011 24570
rect 13169 24512 13174 24568
rect 13230 24512 24950 24568
rect 25006 24512 25011 24568
rect 13169 24510 25011 24512
rect 13169 24507 13235 24510
rect 24945 24507 25011 24510
rect 25681 24570 25747 24573
rect 27520 24570 28000 24600
rect 25681 24568 28000 24570
rect 25681 24512 25686 24568
rect 25742 24512 28000 24568
rect 25681 24510 28000 24512
rect 25681 24507 25747 24510
rect 27520 24480 28000 24510
rect 6361 24434 6427 24437
rect 23197 24434 23263 24437
rect 6361 24432 23263 24434
rect 6361 24376 6366 24432
rect 6422 24376 23202 24432
rect 23258 24376 23263 24432
rect 6361 24374 23263 24376
rect 6361 24371 6427 24374
rect 23197 24371 23263 24374
rect 10277 24232 10597 24233
rect 10277 24168 10285 24232
rect 10349 24168 10365 24232
rect 10429 24168 10445 24232
rect 10509 24168 10525 24232
rect 10589 24168 10597 24232
rect 10277 24167 10597 24168
rect 19610 24232 19930 24233
rect 19610 24168 19618 24232
rect 19682 24168 19698 24232
rect 19762 24168 19778 24232
rect 19842 24168 19858 24232
rect 19922 24168 19930 24232
rect 19610 24167 19930 24168
rect 25497 24026 25563 24029
rect 27520 24026 28000 24056
rect 25497 24024 28000 24026
rect 25497 23968 25502 24024
rect 25558 23968 28000 24024
rect 25497 23966 28000 23968
rect 25497 23963 25563 23966
rect 27520 23936 28000 23966
rect 5993 23890 6059 23893
rect 6126 23890 6132 23892
rect 5993 23888 6132 23890
rect 5993 23832 5998 23888
rect 6054 23832 6132 23888
rect 5993 23830 6132 23832
rect 5993 23827 6059 23830
rect 6126 23828 6132 23830
rect 6196 23828 6202 23892
rect 15101 23890 15167 23893
rect 17861 23890 17927 23893
rect 15101 23888 17927 23890
rect 15101 23832 15106 23888
rect 15162 23832 17866 23888
rect 17922 23832 17927 23888
rect 15101 23830 17927 23832
rect 15101 23827 15167 23830
rect 17861 23827 17927 23830
rect 19885 23890 19951 23893
rect 24669 23890 24735 23893
rect 19885 23888 24735 23890
rect 19885 23832 19890 23888
rect 19946 23832 24674 23888
rect 24730 23832 24735 23888
rect 19885 23830 24735 23832
rect 19885 23827 19951 23830
rect 24669 23827 24735 23830
rect 5610 23688 5930 23689
rect 5610 23624 5618 23688
rect 5682 23624 5698 23688
rect 5762 23624 5778 23688
rect 5842 23624 5858 23688
rect 5922 23624 5930 23688
rect 5610 23623 5930 23624
rect 14944 23688 15264 23689
rect 14944 23624 14952 23688
rect 15016 23624 15032 23688
rect 15096 23624 15112 23688
rect 15176 23624 15192 23688
rect 15256 23624 15264 23688
rect 14944 23623 15264 23624
rect 24277 23688 24597 23689
rect 24277 23624 24285 23688
rect 24349 23624 24365 23688
rect 24429 23624 24445 23688
rect 24509 23624 24525 23688
rect 24589 23624 24597 23688
rect 24277 23623 24597 23624
rect 23197 23482 23263 23485
rect 27520 23482 28000 23512
rect 23197 23480 28000 23482
rect 23197 23424 23202 23480
rect 23258 23424 28000 23480
rect 23197 23422 28000 23424
rect 23197 23419 23263 23422
rect 27520 23392 28000 23422
rect 7097 23346 7163 23349
rect 19057 23346 19123 23349
rect 7097 23344 19123 23346
rect 7097 23288 7102 23344
rect 7158 23288 19062 23344
rect 19118 23288 19123 23344
rect 7097 23286 19123 23288
rect 7097 23283 7163 23286
rect 19057 23283 19123 23286
rect 10961 23212 11027 23213
rect 10910 23210 10916 23212
rect 10870 23150 10916 23210
rect 10980 23208 11027 23212
rect 11022 23152 11027 23208
rect 10910 23148 10916 23150
rect 10980 23148 11027 23152
rect 10961 23147 11027 23148
rect 10277 23144 10597 23145
rect 0 23074 480 23104
rect 10277 23080 10285 23144
rect 10349 23080 10365 23144
rect 10429 23080 10445 23144
rect 10509 23080 10525 23144
rect 10589 23080 10597 23144
rect 10277 23079 10597 23080
rect 19610 23144 19930 23145
rect 19610 23080 19618 23144
rect 19682 23080 19698 23144
rect 19762 23080 19778 23144
rect 19842 23080 19858 23144
rect 19922 23080 19930 23144
rect 19610 23079 19930 23080
rect 12525 23074 12591 23077
rect 14089 23074 14155 23077
rect 0 23014 3250 23074
rect 0 22984 480 23014
rect 3190 21850 3250 23014
rect 12525 23072 14155 23074
rect 12525 23016 12530 23072
rect 12586 23016 14094 23072
rect 14150 23016 14155 23072
rect 12525 23014 14155 23016
rect 12525 23011 12591 23014
rect 14089 23011 14155 23014
rect 14273 23074 14339 23077
rect 14273 23072 19442 23074
rect 14273 23016 14278 23072
rect 14334 23016 19442 23072
rect 14273 23014 19442 23016
rect 14273 23011 14339 23014
rect 8385 22938 8451 22941
rect 14273 22938 14339 22941
rect 8385 22936 14339 22938
rect 8385 22880 8390 22936
rect 8446 22880 14278 22936
rect 14334 22880 14339 22936
rect 8385 22878 14339 22880
rect 8385 22875 8451 22878
rect 14273 22875 14339 22878
rect 7741 22802 7807 22805
rect 16113 22802 16179 22805
rect 7741 22800 16179 22802
rect 7741 22744 7746 22800
rect 7802 22744 16118 22800
rect 16174 22744 16179 22800
rect 7741 22742 16179 22744
rect 7741 22739 7807 22742
rect 16113 22739 16179 22742
rect 5610 22600 5930 22601
rect 5610 22536 5618 22600
rect 5682 22536 5698 22600
rect 5762 22536 5778 22600
rect 5842 22536 5858 22600
rect 5922 22536 5930 22600
rect 5610 22535 5930 22536
rect 14944 22600 15264 22601
rect 14944 22536 14952 22600
rect 15016 22536 15032 22600
rect 15096 22536 15112 22600
rect 15176 22536 15192 22600
rect 15256 22536 15264 22600
rect 14944 22535 15264 22536
rect 4981 22394 5047 22397
rect 18505 22394 18571 22397
rect 4981 22392 18571 22394
rect 4981 22336 4986 22392
rect 5042 22336 18510 22392
rect 18566 22336 18571 22392
rect 4981 22334 18571 22336
rect 19382 22394 19442 23014
rect 25129 22938 25195 22941
rect 27520 22938 28000 22968
rect 25129 22936 28000 22938
rect 25129 22880 25134 22936
rect 25190 22880 28000 22936
rect 25129 22878 28000 22880
rect 25129 22875 25195 22878
rect 27520 22848 28000 22878
rect 24277 22600 24597 22601
rect 24277 22536 24285 22600
rect 24349 22536 24365 22600
rect 24429 22536 24445 22600
rect 24509 22536 24525 22600
rect 24589 22536 24597 22600
rect 24277 22535 24597 22536
rect 22737 22394 22803 22397
rect 25037 22394 25103 22397
rect 19382 22334 20730 22394
rect 4981 22331 5047 22334
rect 18505 22331 18571 22334
rect 16849 22258 16915 22261
rect 20529 22258 20595 22261
rect 16849 22256 20595 22258
rect 16849 22200 16854 22256
rect 16910 22200 20534 22256
rect 20590 22200 20595 22256
rect 16849 22198 20595 22200
rect 20670 22258 20730 22334
rect 22737 22392 25103 22394
rect 22737 22336 22742 22392
rect 22798 22336 25042 22392
rect 25098 22336 25103 22392
rect 22737 22334 25103 22336
rect 22737 22331 22803 22334
rect 25037 22331 25103 22334
rect 27520 22258 28000 22288
rect 20670 22198 28000 22258
rect 16849 22195 16915 22198
rect 20529 22195 20595 22198
rect 27520 22168 28000 22198
rect 10277 22056 10597 22057
rect 10277 21992 10285 22056
rect 10349 21992 10365 22056
rect 10429 21992 10445 22056
rect 10509 21992 10525 22056
rect 10589 21992 10597 22056
rect 10277 21991 10597 21992
rect 19610 22056 19930 22057
rect 19610 21992 19618 22056
rect 19682 21992 19698 22056
rect 19762 21992 19778 22056
rect 19842 21992 19858 22056
rect 19922 21992 19930 22056
rect 19610 21991 19930 21992
rect 10041 21850 10107 21853
rect 3190 21848 10107 21850
rect 3190 21792 10046 21848
rect 10102 21792 10107 21848
rect 3190 21790 10107 21792
rect 10041 21787 10107 21790
rect 10593 21850 10659 21853
rect 13629 21850 13695 21853
rect 10593 21848 13695 21850
rect 10593 21792 10598 21848
rect 10654 21792 13634 21848
rect 13690 21792 13695 21848
rect 10593 21790 13695 21792
rect 10593 21787 10659 21790
rect 13629 21787 13695 21790
rect 18229 21850 18295 21853
rect 24577 21850 24643 21853
rect 18229 21848 24643 21850
rect 18229 21792 18234 21848
rect 18290 21792 24582 21848
rect 24638 21792 24643 21848
rect 18229 21790 24643 21792
rect 18229 21787 18295 21790
rect 24577 21787 24643 21790
rect 24761 21714 24827 21717
rect 27520 21714 28000 21744
rect 24761 21712 28000 21714
rect 24761 21656 24766 21712
rect 24822 21656 28000 21712
rect 24761 21654 28000 21656
rect 24761 21651 24827 21654
rect 27520 21624 28000 21654
rect 5610 21512 5930 21513
rect 5610 21448 5618 21512
rect 5682 21448 5698 21512
rect 5762 21448 5778 21512
rect 5842 21448 5858 21512
rect 5922 21448 5930 21512
rect 5610 21447 5930 21448
rect 14944 21512 15264 21513
rect 14944 21448 14952 21512
rect 15016 21448 15032 21512
rect 15096 21448 15112 21512
rect 15176 21448 15192 21512
rect 15256 21448 15264 21512
rect 14944 21447 15264 21448
rect 24277 21512 24597 21513
rect 24277 21448 24285 21512
rect 24349 21448 24365 21512
rect 24429 21448 24445 21512
rect 24509 21448 24525 21512
rect 24589 21448 24597 21512
rect 24277 21447 24597 21448
rect 16297 21442 16363 21445
rect 18137 21442 18203 21445
rect 19425 21442 19491 21445
rect 20713 21442 20779 21445
rect 16297 21440 20779 21442
rect 16297 21384 16302 21440
rect 16358 21384 18142 21440
rect 18198 21384 19430 21440
rect 19486 21384 20718 21440
rect 20774 21384 20779 21440
rect 16297 21382 20779 21384
rect 16297 21379 16363 21382
rect 18137 21379 18203 21382
rect 19425 21379 19491 21382
rect 20713 21379 20779 21382
rect 2313 21306 2379 21309
rect 16021 21306 16087 21309
rect 2313 21304 16087 21306
rect 2313 21248 2318 21304
rect 2374 21248 16026 21304
rect 16082 21248 16087 21304
rect 2313 21246 16087 21248
rect 2313 21243 2379 21246
rect 16021 21243 16087 21246
rect 16990 21246 24962 21306
rect 12341 21034 12407 21037
rect 16990 21034 17050 21246
rect 24761 21170 24827 21173
rect 12341 21032 17050 21034
rect 12341 20976 12346 21032
rect 12402 20976 17050 21032
rect 12341 20974 17050 20976
rect 17174 21168 24827 21170
rect 17174 21112 24766 21168
rect 24822 21112 24827 21168
rect 17174 21110 24827 21112
rect 24902 21170 24962 21246
rect 27520 21170 28000 21200
rect 24902 21110 28000 21170
rect 12341 20971 12407 20974
rect 10277 20968 10597 20969
rect 10277 20904 10285 20968
rect 10349 20904 10365 20968
rect 10429 20904 10445 20968
rect 10509 20904 10525 20968
rect 10589 20904 10597 20968
rect 10277 20903 10597 20904
rect 12065 20762 12131 20765
rect 17174 20762 17234 21110
rect 24761 21107 24827 21110
rect 27520 21080 28000 21110
rect 19610 20968 19930 20969
rect 19610 20904 19618 20968
rect 19682 20904 19698 20968
rect 19762 20904 19778 20968
rect 19842 20904 19858 20968
rect 19922 20904 19930 20968
rect 19610 20903 19930 20904
rect 21214 20836 21220 20900
rect 21284 20898 21290 20900
rect 21357 20898 21423 20901
rect 21284 20896 21423 20898
rect 21284 20840 21362 20896
rect 21418 20840 21423 20896
rect 21284 20838 21423 20840
rect 21284 20836 21290 20838
rect 21357 20835 21423 20838
rect 25313 20762 25379 20765
rect 12065 20760 17234 20762
rect 12065 20704 12070 20760
rect 12126 20704 17234 20760
rect 12065 20702 17234 20704
rect 17358 20760 25379 20762
rect 17358 20704 25318 20760
rect 25374 20704 25379 20760
rect 17358 20702 25379 20704
rect 12065 20699 12131 20702
rect 12617 20626 12683 20629
rect 17358 20626 17418 20702
rect 25313 20699 25379 20702
rect 12617 20624 17418 20626
rect 12617 20568 12622 20624
rect 12678 20568 17418 20624
rect 12617 20566 17418 20568
rect 12617 20563 12683 20566
rect 23974 20564 23980 20628
rect 24044 20626 24050 20628
rect 27520 20626 28000 20656
rect 24044 20566 28000 20626
rect 24044 20564 24050 20566
rect 27520 20536 28000 20566
rect 5610 20424 5930 20425
rect 5610 20360 5618 20424
rect 5682 20360 5698 20424
rect 5762 20360 5778 20424
rect 5842 20360 5858 20424
rect 5922 20360 5930 20424
rect 5610 20359 5930 20360
rect 14944 20424 15264 20425
rect 14944 20360 14952 20424
rect 15016 20360 15032 20424
rect 15096 20360 15112 20424
rect 15176 20360 15192 20424
rect 15256 20360 15264 20424
rect 14944 20359 15264 20360
rect 24277 20424 24597 20425
rect 24277 20360 24285 20424
rect 24349 20360 24365 20424
rect 24429 20360 24445 20424
rect 24509 20360 24525 20424
rect 24589 20360 24597 20424
rect 24277 20359 24597 20360
rect 19793 20354 19859 20357
rect 24025 20354 24091 20357
rect 19793 20352 24091 20354
rect 19793 20296 19798 20352
rect 19854 20296 24030 20352
rect 24086 20296 24091 20352
rect 19793 20294 24091 20296
rect 19793 20291 19859 20294
rect 24025 20291 24091 20294
rect 3693 20218 3759 20221
rect 11237 20218 11303 20221
rect 3693 20216 11303 20218
rect 3693 20160 3698 20216
rect 3754 20160 11242 20216
rect 11298 20160 11303 20216
rect 3693 20158 11303 20160
rect 3693 20155 3759 20158
rect 11237 20155 11303 20158
rect 19057 20218 19123 20221
rect 23841 20218 23907 20221
rect 19057 20216 23907 20218
rect 19057 20160 19062 20216
rect 19118 20160 23846 20216
rect 23902 20160 23907 20216
rect 19057 20158 23907 20160
rect 19057 20155 19123 20158
rect 23841 20155 23907 20158
rect 933 20082 999 20085
rect 23473 20082 23539 20085
rect 27520 20082 28000 20112
rect 933 20080 23539 20082
rect 933 20024 938 20080
rect 994 20024 23478 20080
rect 23534 20024 23539 20080
rect 933 20022 23539 20024
rect 933 20019 999 20022
rect 23473 20019 23539 20022
rect 25270 20022 28000 20082
rect 10277 19880 10597 19881
rect 10277 19816 10285 19880
rect 10349 19816 10365 19880
rect 10429 19816 10445 19880
rect 10509 19816 10525 19880
rect 10589 19816 10597 19880
rect 10277 19815 10597 19816
rect 19610 19880 19930 19881
rect 19610 19816 19618 19880
rect 19682 19816 19698 19880
rect 19762 19816 19778 19880
rect 19842 19816 19858 19880
rect 19922 19816 19930 19880
rect 19610 19815 19930 19816
rect 11145 19810 11211 19813
rect 16389 19810 16455 19813
rect 16757 19810 16823 19813
rect 11145 19808 16823 19810
rect 11145 19752 11150 19808
rect 11206 19752 16394 19808
rect 16450 19752 16762 19808
rect 16818 19752 16823 19808
rect 11145 19750 16823 19752
rect 11145 19747 11211 19750
rect 16389 19747 16455 19750
rect 16757 19747 16823 19750
rect 13629 19674 13695 19677
rect 25129 19674 25195 19677
rect 13629 19672 25195 19674
rect 13629 19616 13634 19672
rect 13690 19616 25134 19672
rect 25190 19616 25195 19672
rect 13629 19614 25195 19616
rect 13629 19611 13695 19614
rect 25129 19611 25195 19614
rect 25270 19538 25330 20022
rect 27520 19992 28000 20022
rect 14598 19478 25330 19538
rect 5610 19336 5930 19337
rect 5610 19272 5618 19336
rect 5682 19272 5698 19336
rect 5762 19272 5778 19336
rect 5842 19272 5858 19336
rect 5922 19272 5930 19336
rect 5610 19271 5930 19272
rect 9857 19130 9923 19133
rect 14598 19130 14658 19478
rect 16757 19402 16823 19405
rect 22645 19402 22711 19405
rect 16757 19400 22711 19402
rect 16757 19344 16762 19400
rect 16818 19344 22650 19400
rect 22706 19344 22711 19400
rect 16757 19342 22711 19344
rect 16757 19339 16823 19342
rect 22645 19339 22711 19342
rect 25405 19402 25471 19405
rect 27520 19402 28000 19432
rect 25405 19400 28000 19402
rect 25405 19344 25410 19400
rect 25466 19344 28000 19400
rect 25405 19342 28000 19344
rect 25405 19339 25471 19342
rect 14944 19336 15264 19337
rect 14944 19272 14952 19336
rect 15016 19272 15032 19336
rect 15096 19272 15112 19336
rect 15176 19272 15192 19336
rect 15256 19272 15264 19336
rect 14944 19271 15264 19272
rect 24277 19336 24597 19337
rect 24277 19272 24285 19336
rect 24349 19272 24365 19336
rect 24429 19272 24445 19336
rect 24509 19272 24525 19336
rect 24589 19272 24597 19336
rect 27520 19312 28000 19342
rect 24277 19271 24597 19272
rect 9857 19128 14658 19130
rect 9857 19072 9862 19128
rect 9918 19072 14658 19128
rect 9857 19070 14658 19072
rect 14733 19130 14799 19133
rect 15285 19130 15351 19133
rect 14733 19128 15351 19130
rect 14733 19072 14738 19128
rect 14794 19072 15290 19128
rect 15346 19072 15351 19128
rect 14733 19070 15351 19072
rect 9857 19067 9923 19070
rect 14733 19067 14799 19070
rect 15285 19067 15351 19070
rect 18781 19028 18847 19031
rect 18646 19026 18847 19028
rect 4337 18994 4403 18997
rect 15009 18994 15075 18997
rect 4337 18992 15075 18994
rect 4337 18936 4342 18992
rect 4398 18936 15014 18992
rect 15070 18936 15075 18992
rect 4337 18934 15075 18936
rect 4337 18931 4403 18934
rect 15009 18931 15075 18934
rect 18321 18994 18387 18997
rect 18646 18994 18786 19026
rect 18321 18992 18786 18994
rect 18321 18936 18326 18992
rect 18382 18970 18786 18992
rect 18842 18970 18847 19026
rect 18382 18968 18847 18970
rect 18382 18936 18706 18968
rect 18781 18965 18847 18968
rect 18321 18934 18706 18936
rect 18321 18931 18387 18934
rect 20161 18858 20227 18861
rect 23197 18858 23263 18861
rect 20161 18856 23263 18858
rect 20161 18800 20166 18856
rect 20222 18800 23202 18856
rect 23258 18800 23263 18856
rect 20161 18798 23263 18800
rect 20161 18795 20227 18798
rect 23197 18795 23263 18798
rect 25313 18858 25379 18861
rect 27520 18858 28000 18888
rect 25313 18856 28000 18858
rect 25313 18800 25318 18856
rect 25374 18800 28000 18856
rect 25313 18798 28000 18800
rect 25313 18795 25379 18798
rect 10277 18792 10597 18793
rect 10277 18728 10285 18792
rect 10349 18728 10365 18792
rect 10429 18728 10445 18792
rect 10509 18728 10525 18792
rect 10589 18728 10597 18792
rect 10277 18727 10597 18728
rect 19610 18792 19930 18793
rect 19610 18728 19618 18792
rect 19682 18728 19698 18792
rect 19762 18728 19778 18792
rect 19842 18728 19858 18792
rect 19922 18728 19930 18792
rect 27520 18768 28000 18798
rect 19610 18727 19930 18728
rect 13537 18722 13603 18725
rect 19333 18722 19399 18725
rect 13537 18720 19399 18722
rect 13537 18664 13542 18720
rect 13598 18664 19338 18720
rect 19394 18664 19399 18720
rect 13537 18662 19399 18664
rect 13537 18659 13603 18662
rect 19333 18659 19399 18662
rect 1577 18586 1643 18589
rect 18965 18586 19031 18589
rect 1577 18584 19031 18586
rect 1577 18528 1582 18584
rect 1638 18528 18970 18584
rect 19026 18528 19031 18584
rect 1577 18526 19031 18528
rect 1577 18523 1643 18526
rect 18965 18523 19031 18526
rect 16389 18450 16455 18453
rect 20529 18450 20595 18453
rect 23657 18450 23723 18453
rect 16389 18448 20595 18450
rect 16389 18392 16394 18448
rect 16450 18392 20534 18448
rect 20590 18392 20595 18448
rect 16389 18390 20595 18392
rect 16389 18387 16455 18390
rect 20529 18387 20595 18390
rect 20670 18448 23723 18450
rect 20670 18392 23662 18448
rect 23718 18392 23723 18448
rect 20670 18390 23723 18392
rect 10869 18314 10935 18317
rect 11789 18314 11855 18317
rect 12433 18314 12499 18317
rect 10869 18312 12499 18314
rect 10869 18256 10874 18312
rect 10930 18256 11794 18312
rect 11850 18256 12438 18312
rect 12494 18256 12499 18312
rect 10869 18254 12499 18256
rect 10869 18251 10935 18254
rect 11789 18251 11855 18254
rect 12433 18251 12499 18254
rect 18137 18314 18203 18317
rect 20670 18314 20730 18390
rect 23657 18387 23723 18390
rect 24209 18450 24275 18453
rect 24209 18448 24778 18450
rect 24209 18392 24214 18448
rect 24270 18392 24778 18448
rect 24209 18390 24778 18392
rect 24209 18387 24275 18390
rect 18137 18312 20730 18314
rect 18137 18256 18142 18312
rect 18198 18256 20730 18312
rect 18137 18254 20730 18256
rect 24718 18314 24778 18390
rect 27520 18314 28000 18344
rect 24718 18254 28000 18314
rect 18137 18251 18203 18254
rect 5610 18248 5930 18249
rect 5610 18184 5618 18248
rect 5682 18184 5698 18248
rect 5762 18184 5778 18248
rect 5842 18184 5858 18248
rect 5922 18184 5930 18248
rect 5610 18183 5930 18184
rect 14944 18248 15264 18249
rect 14944 18184 14952 18248
rect 15016 18184 15032 18248
rect 15096 18184 15112 18248
rect 15176 18184 15192 18248
rect 15256 18184 15264 18248
rect 14944 18183 15264 18184
rect 24277 18248 24597 18249
rect 24277 18184 24285 18248
rect 24349 18184 24365 18248
rect 24429 18184 24445 18248
rect 24509 18184 24525 18248
rect 24589 18184 24597 18248
rect 27520 18224 28000 18254
rect 24277 18183 24597 18184
rect 21725 18178 21791 18181
rect 23933 18178 23999 18181
rect 21725 18176 23999 18178
rect 21725 18120 21730 18176
rect 21786 18120 23938 18176
rect 23994 18120 23999 18176
rect 21725 18118 23999 18120
rect 21725 18115 21791 18118
rect 23933 18115 23999 18118
rect 13905 18042 13971 18045
rect 13905 18040 22018 18042
rect 13905 17984 13910 18040
rect 13966 17984 22018 18040
rect 13905 17982 22018 17984
rect 13905 17979 13971 17982
rect 2957 17906 3023 17909
rect 13445 17906 13511 17909
rect 2957 17904 13511 17906
rect 2957 17848 2962 17904
rect 3018 17848 13450 17904
rect 13506 17848 13511 17904
rect 2957 17846 13511 17848
rect 2957 17843 3023 17846
rect 13445 17843 13511 17846
rect 19241 17906 19307 17909
rect 21817 17906 21883 17909
rect 19241 17904 21883 17906
rect 19241 17848 19246 17904
rect 19302 17848 21822 17904
rect 21878 17848 21883 17904
rect 19241 17846 21883 17848
rect 21958 17906 22018 17982
rect 22185 17906 22251 17909
rect 21958 17904 22251 17906
rect 21958 17848 22190 17904
rect 22246 17848 22251 17904
rect 21958 17846 22251 17848
rect 19241 17843 19307 17846
rect 21817 17843 21883 17846
rect 22185 17843 22251 17846
rect 20529 17770 20595 17773
rect 23841 17770 23907 17773
rect 20529 17768 23907 17770
rect 20529 17712 20534 17768
rect 20590 17712 23846 17768
rect 23902 17712 23907 17768
rect 20529 17710 23907 17712
rect 20529 17707 20595 17710
rect 23841 17707 23907 17710
rect 24761 17770 24827 17773
rect 27520 17770 28000 17800
rect 24761 17768 28000 17770
rect 24761 17712 24766 17768
rect 24822 17712 28000 17768
rect 24761 17710 28000 17712
rect 24761 17707 24827 17710
rect 10277 17704 10597 17705
rect 10277 17640 10285 17704
rect 10349 17640 10365 17704
rect 10429 17640 10445 17704
rect 10509 17640 10525 17704
rect 10589 17640 10597 17704
rect 10277 17639 10597 17640
rect 19610 17704 19930 17705
rect 19610 17640 19618 17704
rect 19682 17640 19698 17704
rect 19762 17640 19778 17704
rect 19842 17640 19858 17704
rect 19922 17640 19930 17704
rect 27520 17680 28000 17710
rect 19610 17639 19930 17640
rect 15101 17498 15167 17501
rect 18229 17498 18295 17501
rect 15101 17496 18295 17498
rect 15101 17440 15106 17496
rect 15162 17440 18234 17496
rect 18290 17440 18295 17496
rect 15101 17438 18295 17440
rect 15101 17435 15167 17438
rect 18229 17435 18295 17438
rect 25405 17226 25471 17229
rect 27520 17226 28000 17256
rect 25405 17224 28000 17226
rect 25405 17168 25410 17224
rect 25466 17168 28000 17224
rect 25405 17166 28000 17168
rect 25405 17163 25471 17166
rect 5610 17160 5930 17161
rect 5610 17096 5618 17160
rect 5682 17096 5698 17160
rect 5762 17096 5778 17160
rect 5842 17096 5858 17160
rect 5922 17096 5930 17160
rect 5610 17095 5930 17096
rect 14944 17160 15264 17161
rect 14944 17096 14952 17160
rect 15016 17096 15032 17160
rect 15096 17096 15112 17160
rect 15176 17096 15192 17160
rect 15256 17096 15264 17160
rect 14944 17095 15264 17096
rect 24277 17160 24597 17161
rect 24277 17096 24285 17160
rect 24349 17096 24365 17160
rect 24429 17096 24445 17160
rect 24509 17096 24525 17160
rect 24589 17096 24597 17160
rect 27520 17136 28000 17166
rect 24277 17095 24597 17096
rect 15469 16954 15535 16957
rect 25129 16954 25195 16957
rect 15469 16952 25195 16954
rect 15469 16896 15474 16952
rect 15530 16896 25134 16952
rect 25190 16896 25195 16952
rect 15469 16894 25195 16896
rect 15469 16891 15535 16894
rect 25129 16891 25195 16894
rect 15745 16818 15811 16821
rect 20713 16818 20779 16821
rect 23657 16818 23723 16821
rect 25037 16818 25103 16821
rect 15745 16816 25103 16818
rect 15745 16760 15750 16816
rect 15806 16760 20718 16816
rect 20774 16760 23662 16816
rect 23718 16760 25042 16816
rect 25098 16760 25103 16816
rect 15745 16758 25103 16760
rect 15745 16755 15811 16758
rect 20713 16755 20779 16758
rect 23657 16755 23723 16758
rect 25037 16755 25103 16758
rect 10277 16616 10597 16617
rect 10277 16552 10285 16616
rect 10349 16552 10365 16616
rect 10429 16552 10445 16616
rect 10509 16552 10525 16616
rect 10589 16552 10597 16616
rect 10277 16551 10597 16552
rect 19610 16616 19930 16617
rect 19610 16552 19618 16616
rect 19682 16552 19698 16616
rect 19762 16552 19778 16616
rect 19842 16552 19858 16616
rect 19922 16552 19930 16616
rect 19610 16551 19930 16552
rect 21633 16546 21699 16549
rect 23933 16546 23999 16549
rect 21633 16544 23999 16546
rect 21633 16488 21638 16544
rect 21694 16488 23938 16544
rect 23994 16488 23999 16544
rect 21633 16486 23999 16488
rect 21633 16483 21699 16486
rect 23933 16483 23999 16486
rect 24209 16546 24275 16549
rect 27520 16546 28000 16576
rect 24209 16544 28000 16546
rect 24209 16488 24214 16544
rect 24270 16488 28000 16544
rect 24209 16486 28000 16488
rect 24209 16483 24275 16486
rect 27520 16456 28000 16486
rect 21081 16410 21147 16413
rect 25221 16410 25287 16413
rect 21081 16408 25287 16410
rect 21081 16352 21086 16408
rect 21142 16352 25226 16408
rect 25282 16352 25287 16408
rect 21081 16350 25287 16352
rect 21081 16347 21147 16350
rect 25221 16347 25287 16350
rect 5610 16072 5930 16073
rect 5610 16008 5618 16072
rect 5682 16008 5698 16072
rect 5762 16008 5778 16072
rect 5842 16008 5858 16072
rect 5922 16008 5930 16072
rect 5610 16007 5930 16008
rect 14944 16072 15264 16073
rect 14944 16008 14952 16072
rect 15016 16008 15032 16072
rect 15096 16008 15112 16072
rect 15176 16008 15192 16072
rect 15256 16008 15264 16072
rect 14944 16007 15264 16008
rect 24277 16072 24597 16073
rect 24277 16008 24285 16072
rect 24349 16008 24365 16072
rect 24429 16008 24445 16072
rect 24509 16008 24525 16072
rect 24589 16008 24597 16072
rect 24277 16007 24597 16008
rect 25405 16002 25471 16005
rect 27520 16002 28000 16032
rect 25405 16000 28000 16002
rect 25405 15944 25410 16000
rect 25466 15944 28000 16000
rect 25405 15942 28000 15944
rect 25405 15939 25471 15942
rect 27520 15912 28000 15942
rect 10277 15528 10597 15529
rect 10277 15464 10285 15528
rect 10349 15464 10365 15528
rect 10429 15464 10445 15528
rect 10509 15464 10525 15528
rect 10589 15464 10597 15528
rect 10277 15463 10597 15464
rect 19610 15528 19930 15529
rect 19610 15464 19618 15528
rect 19682 15464 19698 15528
rect 19762 15464 19778 15528
rect 19842 15464 19858 15528
rect 19922 15464 19930 15528
rect 19610 15463 19930 15464
rect 25405 15458 25471 15461
rect 27520 15458 28000 15488
rect 25405 15456 28000 15458
rect 25405 15400 25410 15456
rect 25466 15400 28000 15456
rect 25405 15398 28000 15400
rect 25405 15395 25471 15398
rect 27520 15368 28000 15398
rect 23565 15050 23631 15053
rect 24117 15050 24183 15053
rect 23565 15048 24183 15050
rect 23565 14992 23570 15048
rect 23626 14992 24122 15048
rect 24178 14992 24183 15048
rect 23565 14990 24183 14992
rect 23565 14987 23631 14990
rect 24117 14987 24183 14990
rect 5610 14984 5930 14985
rect 5610 14920 5618 14984
rect 5682 14920 5698 14984
rect 5762 14920 5778 14984
rect 5842 14920 5858 14984
rect 5922 14920 5930 14984
rect 5610 14919 5930 14920
rect 14944 14984 15264 14985
rect 14944 14920 14952 14984
rect 15016 14920 15032 14984
rect 15096 14920 15112 14984
rect 15176 14920 15192 14984
rect 15256 14920 15264 14984
rect 14944 14919 15264 14920
rect 24277 14984 24597 14985
rect 24277 14920 24285 14984
rect 24349 14920 24365 14984
rect 24429 14920 24445 14984
rect 24509 14920 24525 14984
rect 24589 14920 24597 14984
rect 24277 14919 24597 14920
rect 24669 14914 24735 14917
rect 27520 14914 28000 14944
rect 24669 14912 28000 14914
rect 24669 14856 24674 14912
rect 24730 14856 28000 14912
rect 24669 14854 28000 14856
rect 24669 14851 24735 14854
rect 27520 14824 28000 14854
rect 12249 14642 12315 14645
rect 22921 14642 22987 14645
rect 12249 14640 22987 14642
rect 12249 14584 12254 14640
rect 12310 14584 22926 14640
rect 22982 14584 22987 14640
rect 12249 14582 22987 14584
rect 12249 14579 12315 14582
rect 22921 14579 22987 14582
rect 10277 14440 10597 14441
rect 10277 14376 10285 14440
rect 10349 14376 10365 14440
rect 10429 14376 10445 14440
rect 10509 14376 10525 14440
rect 10589 14376 10597 14440
rect 10277 14375 10597 14376
rect 19610 14440 19930 14441
rect 19610 14376 19618 14440
rect 19682 14376 19698 14440
rect 19762 14376 19778 14440
rect 19842 14376 19858 14440
rect 19922 14376 19930 14440
rect 19610 14375 19930 14376
rect 24853 14370 24919 14373
rect 27520 14370 28000 14400
rect 24853 14368 28000 14370
rect 24853 14312 24858 14368
rect 24914 14312 28000 14368
rect 24853 14310 28000 14312
rect 24853 14307 24919 14310
rect 27520 14280 28000 14310
rect 5610 13896 5930 13897
rect 5610 13832 5618 13896
rect 5682 13832 5698 13896
rect 5762 13832 5778 13896
rect 5842 13832 5858 13896
rect 5922 13832 5930 13896
rect 5610 13831 5930 13832
rect 14944 13896 15264 13897
rect 14944 13832 14952 13896
rect 15016 13832 15032 13896
rect 15096 13832 15112 13896
rect 15176 13832 15192 13896
rect 15256 13832 15264 13896
rect 14944 13831 15264 13832
rect 24277 13896 24597 13897
rect 24277 13832 24285 13896
rect 24349 13832 24365 13896
rect 24429 13832 24445 13896
rect 24509 13832 24525 13896
rect 24589 13832 24597 13896
rect 24277 13831 24597 13832
rect 0 13690 480 13720
rect 1485 13690 1551 13693
rect 0 13688 1551 13690
rect 0 13632 1490 13688
rect 1546 13632 1551 13688
rect 0 13630 1551 13632
rect 0 13600 480 13630
rect 1485 13627 1551 13630
rect 14365 13690 14431 13693
rect 24577 13690 24643 13693
rect 14365 13688 24643 13690
rect 14365 13632 14370 13688
rect 14426 13632 24582 13688
rect 24638 13632 24643 13688
rect 14365 13630 24643 13632
rect 14365 13627 14431 13630
rect 24577 13627 24643 13630
rect 24761 13690 24827 13693
rect 27520 13690 28000 13720
rect 24761 13688 28000 13690
rect 24761 13632 24766 13688
rect 24822 13632 28000 13688
rect 24761 13630 28000 13632
rect 24761 13627 24827 13630
rect 27520 13600 28000 13630
rect 2773 13554 2839 13557
rect 11697 13554 11763 13557
rect 2773 13552 11763 13554
rect 2773 13496 2778 13552
rect 2834 13496 11702 13552
rect 11758 13496 11763 13552
rect 2773 13494 11763 13496
rect 2773 13491 2839 13494
rect 11697 13491 11763 13494
rect 10277 13352 10597 13353
rect 10277 13288 10285 13352
rect 10349 13288 10365 13352
rect 10429 13288 10445 13352
rect 10509 13288 10525 13352
rect 10589 13288 10597 13352
rect 10277 13287 10597 13288
rect 19610 13352 19930 13353
rect 19610 13288 19618 13352
rect 19682 13288 19698 13352
rect 19762 13288 19778 13352
rect 19842 13288 19858 13352
rect 19922 13288 19930 13352
rect 19610 13287 19930 13288
rect 381 13146 447 13149
rect 13353 13146 13419 13149
rect 381 13144 13419 13146
rect 381 13088 386 13144
rect 442 13088 13358 13144
rect 13414 13088 13419 13144
rect 381 13086 13419 13088
rect 381 13083 447 13086
rect 13353 13083 13419 13086
rect 23657 13146 23723 13149
rect 27520 13146 28000 13176
rect 23657 13144 28000 13146
rect 23657 13088 23662 13144
rect 23718 13088 28000 13144
rect 23657 13086 28000 13088
rect 23657 13083 23723 13086
rect 27520 13056 28000 13086
rect 2037 13010 2103 13013
rect 2865 13010 2931 13013
rect 12065 13010 12131 13013
rect 2037 13008 12131 13010
rect 2037 12952 2042 13008
rect 2098 12952 2870 13008
rect 2926 12952 12070 13008
rect 12126 12952 12131 13008
rect 2037 12950 12131 12952
rect 2037 12947 2103 12950
rect 2865 12947 2931 12950
rect 12065 12947 12131 12950
rect 18229 13010 18295 13013
rect 24577 13010 24643 13013
rect 18229 13008 24643 13010
rect 18229 12952 18234 13008
rect 18290 12952 24582 13008
rect 24638 12952 24643 13008
rect 18229 12950 24643 12952
rect 18229 12947 18295 12950
rect 24577 12947 24643 12950
rect 5610 12808 5930 12809
rect 5610 12744 5618 12808
rect 5682 12744 5698 12808
rect 5762 12744 5778 12808
rect 5842 12744 5858 12808
rect 5922 12744 5930 12808
rect 5610 12743 5930 12744
rect 14944 12808 15264 12809
rect 14944 12744 14952 12808
rect 15016 12744 15032 12808
rect 15096 12744 15112 12808
rect 15176 12744 15192 12808
rect 15256 12744 15264 12808
rect 14944 12743 15264 12744
rect 24277 12808 24597 12809
rect 24277 12744 24285 12808
rect 24349 12744 24365 12808
rect 24429 12744 24445 12808
rect 24509 12744 24525 12808
rect 24589 12744 24597 12808
rect 24277 12743 24597 12744
rect 24761 12602 24827 12605
rect 27520 12602 28000 12632
rect 24761 12600 28000 12602
rect 24761 12544 24766 12600
rect 24822 12544 28000 12600
rect 24761 12542 28000 12544
rect 24761 12539 24827 12542
rect 27520 12512 28000 12542
rect 13353 12466 13419 12469
rect 15929 12466 15995 12469
rect 18505 12466 18571 12469
rect 22277 12466 22343 12469
rect 13353 12464 22343 12466
rect 13353 12408 13358 12464
rect 13414 12408 15934 12464
rect 15990 12408 18510 12464
rect 18566 12408 22282 12464
rect 22338 12408 22343 12464
rect 13353 12406 22343 12408
rect 13353 12403 13419 12406
rect 15929 12403 15995 12406
rect 18505 12403 18571 12406
rect 22277 12403 22343 12406
rect 18873 12330 18939 12333
rect 18830 12328 18939 12330
rect 18830 12272 18878 12328
rect 18934 12272 18939 12328
rect 18830 12267 18939 12272
rect 10277 12264 10597 12265
rect 10277 12200 10285 12264
rect 10349 12200 10365 12264
rect 10429 12200 10445 12264
rect 10509 12200 10525 12264
rect 10589 12200 10597 12264
rect 10277 12199 10597 12200
rect 18830 12061 18890 12267
rect 19610 12264 19930 12265
rect 19610 12200 19618 12264
rect 19682 12200 19698 12264
rect 19762 12200 19778 12264
rect 19842 12200 19858 12264
rect 19922 12200 19930 12264
rect 19610 12199 19930 12200
rect 18830 12056 18939 12061
rect 18830 12000 18878 12056
rect 18934 12000 18939 12056
rect 18830 11998 18939 12000
rect 18873 11995 18939 11998
rect 24761 12058 24827 12061
rect 27520 12058 28000 12088
rect 24761 12056 28000 12058
rect 24761 12000 24766 12056
rect 24822 12000 28000 12056
rect 24761 11998 28000 12000
rect 24761 11995 24827 11998
rect 27520 11968 28000 11998
rect 22001 11786 22067 11789
rect 23657 11786 23723 11789
rect 22001 11784 23723 11786
rect 22001 11728 22006 11784
rect 22062 11728 23662 11784
rect 23718 11728 23723 11784
rect 22001 11726 23723 11728
rect 22001 11723 22067 11726
rect 23657 11723 23723 11726
rect 5610 11720 5930 11721
rect 5610 11656 5618 11720
rect 5682 11656 5698 11720
rect 5762 11656 5778 11720
rect 5842 11656 5858 11720
rect 5922 11656 5930 11720
rect 5610 11655 5930 11656
rect 14944 11720 15264 11721
rect 14944 11656 14952 11720
rect 15016 11656 15032 11720
rect 15096 11656 15112 11720
rect 15176 11656 15192 11720
rect 15256 11656 15264 11720
rect 14944 11655 15264 11656
rect 24277 11720 24597 11721
rect 24277 11656 24285 11720
rect 24349 11656 24365 11720
rect 24429 11656 24445 11720
rect 24509 11656 24525 11720
rect 24589 11656 24597 11720
rect 24277 11655 24597 11656
rect 24761 11650 24827 11653
rect 26877 11650 26943 11653
rect 24761 11648 26943 11650
rect 24761 11592 24766 11648
rect 24822 11592 26882 11648
rect 26938 11592 26943 11648
rect 24761 11590 26943 11592
rect 24761 11587 24827 11590
rect 26877 11587 26943 11590
rect 25221 11514 25287 11517
rect 27520 11514 28000 11544
rect 25221 11512 28000 11514
rect 25221 11456 25226 11512
rect 25282 11456 28000 11512
rect 25221 11454 28000 11456
rect 25221 11451 25287 11454
rect 27520 11424 28000 11454
rect 10277 11176 10597 11177
rect 10277 11112 10285 11176
rect 10349 11112 10365 11176
rect 10429 11112 10445 11176
rect 10509 11112 10525 11176
rect 10589 11112 10597 11176
rect 10277 11111 10597 11112
rect 19610 11176 19930 11177
rect 19610 11112 19618 11176
rect 19682 11112 19698 11176
rect 19762 11112 19778 11176
rect 19842 11112 19858 11176
rect 19922 11112 19930 11176
rect 19610 11111 19930 11112
rect 24577 10834 24643 10837
rect 27520 10834 28000 10864
rect 24577 10832 28000 10834
rect 24577 10776 24582 10832
rect 24638 10776 28000 10832
rect 24577 10774 28000 10776
rect 24577 10771 24643 10774
rect 27520 10744 28000 10774
rect 5610 10632 5930 10633
rect 5610 10568 5618 10632
rect 5682 10568 5698 10632
rect 5762 10568 5778 10632
rect 5842 10568 5858 10632
rect 5922 10568 5930 10632
rect 5610 10567 5930 10568
rect 14944 10632 15264 10633
rect 14944 10568 14952 10632
rect 15016 10568 15032 10632
rect 15096 10568 15112 10632
rect 15176 10568 15192 10632
rect 15256 10568 15264 10632
rect 14944 10567 15264 10568
rect 24277 10632 24597 10633
rect 24277 10568 24285 10632
rect 24349 10568 24365 10632
rect 24429 10568 24445 10632
rect 24509 10568 24525 10632
rect 24589 10568 24597 10632
rect 24277 10567 24597 10568
rect 24761 10562 24827 10565
rect 25589 10562 25655 10565
rect 24761 10560 25655 10562
rect 24761 10504 24766 10560
rect 24822 10504 25594 10560
rect 25650 10504 25655 10560
rect 24761 10502 25655 10504
rect 24761 10499 24827 10502
rect 25589 10499 25655 10502
rect 25221 10290 25287 10293
rect 27520 10290 28000 10320
rect 25221 10288 28000 10290
rect 25221 10232 25226 10288
rect 25282 10232 28000 10288
rect 25221 10230 28000 10232
rect 25221 10227 25287 10230
rect 27520 10200 28000 10230
rect 10277 10088 10597 10089
rect 10277 10024 10285 10088
rect 10349 10024 10365 10088
rect 10429 10024 10445 10088
rect 10509 10024 10525 10088
rect 10589 10024 10597 10088
rect 10277 10023 10597 10024
rect 19610 10088 19930 10089
rect 19610 10024 19618 10088
rect 19682 10024 19698 10088
rect 19762 10024 19778 10088
rect 19842 10024 19858 10088
rect 19922 10024 19930 10088
rect 19610 10023 19930 10024
rect 24577 9746 24643 9749
rect 27520 9746 28000 9776
rect 24577 9744 28000 9746
rect 24577 9688 24582 9744
rect 24638 9688 28000 9744
rect 24577 9686 28000 9688
rect 24577 9683 24643 9686
rect 27520 9656 28000 9686
rect 5610 9544 5930 9545
rect 5610 9480 5618 9544
rect 5682 9480 5698 9544
rect 5762 9480 5778 9544
rect 5842 9480 5858 9544
rect 5922 9480 5930 9544
rect 5610 9479 5930 9480
rect 14944 9544 15264 9545
rect 14944 9480 14952 9544
rect 15016 9480 15032 9544
rect 15096 9480 15112 9544
rect 15176 9480 15192 9544
rect 15256 9480 15264 9544
rect 14944 9479 15264 9480
rect 24277 9544 24597 9545
rect 24277 9480 24285 9544
rect 24349 9480 24365 9544
rect 24429 9480 24445 9544
rect 24509 9480 24525 9544
rect 24589 9480 24597 9544
rect 24277 9479 24597 9480
rect 24393 9202 24459 9205
rect 27520 9202 28000 9232
rect 24393 9200 28000 9202
rect 24393 9144 24398 9200
rect 24454 9144 28000 9200
rect 24393 9142 28000 9144
rect 24393 9139 24459 9142
rect 27520 9112 28000 9142
rect 10277 9000 10597 9001
rect 10277 8936 10285 9000
rect 10349 8936 10365 9000
rect 10429 8936 10445 9000
rect 10509 8936 10525 9000
rect 10589 8936 10597 9000
rect 10277 8935 10597 8936
rect 19610 9000 19930 9001
rect 19610 8936 19618 9000
rect 19682 8936 19698 9000
rect 19762 8936 19778 9000
rect 19842 8936 19858 9000
rect 19922 8936 19930 9000
rect 19610 8935 19930 8936
rect 24393 8658 24459 8661
rect 24669 8658 24735 8661
rect 27520 8658 28000 8688
rect 24393 8656 28000 8658
rect 24393 8600 24398 8656
rect 24454 8600 24674 8656
rect 24730 8600 28000 8656
rect 24393 8598 28000 8600
rect 24393 8595 24459 8598
rect 24669 8595 24735 8598
rect 27520 8568 28000 8598
rect 5610 8456 5930 8457
rect 5610 8392 5618 8456
rect 5682 8392 5698 8456
rect 5762 8392 5778 8456
rect 5842 8392 5858 8456
rect 5922 8392 5930 8456
rect 5610 8391 5930 8392
rect 14944 8456 15264 8457
rect 14944 8392 14952 8456
rect 15016 8392 15032 8456
rect 15096 8392 15112 8456
rect 15176 8392 15192 8456
rect 15256 8392 15264 8456
rect 14944 8391 15264 8392
rect 24277 8456 24597 8457
rect 24277 8392 24285 8456
rect 24349 8392 24365 8456
rect 24429 8392 24445 8456
rect 24509 8392 24525 8456
rect 24589 8392 24597 8456
rect 24277 8391 24597 8392
rect 23657 7978 23723 7981
rect 27520 7978 28000 8008
rect 23657 7976 28000 7978
rect 23657 7920 23662 7976
rect 23718 7920 28000 7976
rect 23657 7918 28000 7920
rect 23657 7915 23723 7918
rect 10277 7912 10597 7913
rect 10277 7848 10285 7912
rect 10349 7848 10365 7912
rect 10429 7848 10445 7912
rect 10509 7848 10525 7912
rect 10589 7848 10597 7912
rect 10277 7847 10597 7848
rect 19610 7912 19930 7913
rect 19610 7848 19618 7912
rect 19682 7848 19698 7912
rect 19762 7848 19778 7912
rect 19842 7848 19858 7912
rect 19922 7848 19930 7912
rect 27520 7888 28000 7918
rect 19610 7847 19930 7848
rect 24669 7434 24735 7437
rect 27520 7434 28000 7464
rect 24669 7432 28000 7434
rect 24669 7376 24674 7432
rect 24730 7376 28000 7432
rect 24669 7374 28000 7376
rect 24669 7371 24735 7374
rect 5610 7368 5930 7369
rect 5610 7304 5618 7368
rect 5682 7304 5698 7368
rect 5762 7304 5778 7368
rect 5842 7304 5858 7368
rect 5922 7304 5930 7368
rect 5610 7303 5930 7304
rect 14944 7368 15264 7369
rect 14944 7304 14952 7368
rect 15016 7304 15032 7368
rect 15096 7304 15112 7368
rect 15176 7304 15192 7368
rect 15256 7304 15264 7368
rect 14944 7303 15264 7304
rect 24277 7368 24597 7369
rect 24277 7304 24285 7368
rect 24349 7304 24365 7368
rect 24429 7304 24445 7368
rect 24509 7304 24525 7368
rect 24589 7304 24597 7368
rect 27520 7344 28000 7374
rect 24277 7303 24597 7304
rect 21633 6890 21699 6893
rect 27520 6890 28000 6920
rect 21633 6888 28000 6890
rect 21633 6832 21638 6888
rect 21694 6832 28000 6888
rect 21633 6830 28000 6832
rect 21633 6827 21699 6830
rect 10277 6824 10597 6825
rect 10277 6760 10285 6824
rect 10349 6760 10365 6824
rect 10429 6760 10445 6824
rect 10509 6760 10525 6824
rect 10589 6760 10597 6824
rect 10277 6759 10597 6760
rect 19610 6824 19930 6825
rect 19610 6760 19618 6824
rect 19682 6760 19698 6824
rect 19762 6760 19778 6824
rect 19842 6760 19858 6824
rect 19922 6760 19930 6824
rect 27520 6800 28000 6830
rect 19610 6759 19930 6760
rect 20345 6482 20411 6485
rect 20345 6480 24962 6482
rect 20345 6424 20350 6480
rect 20406 6424 24962 6480
rect 20345 6422 24962 6424
rect 20345 6419 20411 6422
rect 24902 6346 24962 6422
rect 27520 6346 28000 6376
rect 24902 6286 28000 6346
rect 5610 6280 5930 6281
rect 5610 6216 5618 6280
rect 5682 6216 5698 6280
rect 5762 6216 5778 6280
rect 5842 6216 5858 6280
rect 5922 6216 5930 6280
rect 5610 6215 5930 6216
rect 14944 6280 15264 6281
rect 14944 6216 14952 6280
rect 15016 6216 15032 6280
rect 15096 6216 15112 6280
rect 15176 6216 15192 6280
rect 15256 6216 15264 6280
rect 14944 6215 15264 6216
rect 24277 6280 24597 6281
rect 24277 6216 24285 6280
rect 24349 6216 24365 6280
rect 24429 6216 24445 6280
rect 24509 6216 24525 6280
rect 24589 6216 24597 6280
rect 27520 6256 28000 6286
rect 24277 6215 24597 6216
rect 20069 5802 20135 5805
rect 27520 5802 28000 5832
rect 20069 5800 28000 5802
rect 20069 5744 20074 5800
rect 20130 5744 28000 5800
rect 20069 5742 28000 5744
rect 20069 5739 20135 5742
rect 10277 5736 10597 5737
rect 10277 5672 10285 5736
rect 10349 5672 10365 5736
rect 10429 5672 10445 5736
rect 10509 5672 10525 5736
rect 10589 5672 10597 5736
rect 10277 5671 10597 5672
rect 19610 5736 19930 5737
rect 19610 5672 19618 5736
rect 19682 5672 19698 5736
rect 19762 5672 19778 5736
rect 19842 5672 19858 5736
rect 19922 5672 19930 5736
rect 27520 5712 28000 5742
rect 19610 5671 19930 5672
rect 18321 5394 18387 5397
rect 23933 5394 23999 5397
rect 18321 5392 23999 5394
rect 18321 5336 18326 5392
rect 18382 5336 23938 5392
rect 23994 5336 23999 5392
rect 18321 5334 23999 5336
rect 18321 5331 18387 5334
rect 23933 5331 23999 5334
rect 5610 5192 5930 5193
rect 5610 5128 5618 5192
rect 5682 5128 5698 5192
rect 5762 5128 5778 5192
rect 5842 5128 5858 5192
rect 5922 5128 5930 5192
rect 5610 5127 5930 5128
rect 14944 5192 15264 5193
rect 14944 5128 14952 5192
rect 15016 5128 15032 5192
rect 15096 5128 15112 5192
rect 15176 5128 15192 5192
rect 15256 5128 15264 5192
rect 14944 5127 15264 5128
rect 24277 5192 24597 5193
rect 24277 5128 24285 5192
rect 24349 5128 24365 5192
rect 24429 5128 24445 5192
rect 24509 5128 24525 5192
rect 24589 5128 24597 5192
rect 24277 5127 24597 5128
rect 20437 5122 20503 5125
rect 23473 5122 23539 5125
rect 20437 5120 23539 5122
rect 20437 5064 20442 5120
rect 20498 5064 23478 5120
rect 23534 5064 23539 5120
rect 20437 5062 23539 5064
rect 20437 5059 20503 5062
rect 23473 5059 23539 5062
rect 25221 5122 25287 5125
rect 27520 5122 28000 5152
rect 25221 5120 28000 5122
rect 25221 5064 25226 5120
rect 25282 5064 28000 5120
rect 25221 5062 28000 5064
rect 25221 5059 25287 5062
rect 27520 5032 28000 5062
rect 19057 4850 19123 4853
rect 24761 4850 24827 4853
rect 19057 4848 24827 4850
rect 19057 4792 19062 4848
rect 19118 4792 24766 4848
rect 24822 4792 24827 4848
rect 19057 4790 24827 4792
rect 19057 4787 19123 4790
rect 24761 4787 24827 4790
rect 10277 4648 10597 4649
rect 10277 4584 10285 4648
rect 10349 4584 10365 4648
rect 10429 4584 10445 4648
rect 10509 4584 10525 4648
rect 10589 4584 10597 4648
rect 10277 4583 10597 4584
rect 19610 4648 19930 4649
rect 19610 4584 19618 4648
rect 19682 4584 19698 4648
rect 19762 4584 19778 4648
rect 19842 4584 19858 4648
rect 19922 4584 19930 4648
rect 19610 4583 19930 4584
rect 24577 4578 24643 4581
rect 27520 4578 28000 4608
rect 24577 4576 28000 4578
rect 24577 4520 24582 4576
rect 24638 4520 28000 4576
rect 24577 4518 28000 4520
rect 24577 4515 24643 4518
rect 27520 4488 28000 4518
rect 0 4442 480 4472
rect 2865 4442 2931 4445
rect 0 4440 2931 4442
rect 0 4384 2870 4440
rect 2926 4384 2931 4440
rect 0 4382 2931 4384
rect 0 4352 480 4382
rect 2865 4379 2931 4382
rect 5610 4104 5930 4105
rect 5610 4040 5618 4104
rect 5682 4040 5698 4104
rect 5762 4040 5778 4104
rect 5842 4040 5858 4104
rect 5922 4040 5930 4104
rect 5610 4039 5930 4040
rect 14944 4104 15264 4105
rect 14944 4040 14952 4104
rect 15016 4040 15032 4104
rect 15096 4040 15112 4104
rect 15176 4040 15192 4104
rect 15256 4040 15264 4104
rect 14944 4039 15264 4040
rect 24277 4104 24597 4105
rect 24277 4040 24285 4104
rect 24349 4040 24365 4104
rect 24429 4040 24445 4104
rect 24509 4040 24525 4104
rect 24589 4040 24597 4104
rect 24277 4039 24597 4040
rect 25221 4034 25287 4037
rect 27520 4034 28000 4064
rect 25221 4032 28000 4034
rect 25221 3976 25226 4032
rect 25282 3976 28000 4032
rect 25221 3974 28000 3976
rect 25221 3971 25287 3974
rect 27520 3944 28000 3974
rect 18873 3762 18939 3765
rect 24761 3762 24827 3765
rect 18873 3760 24827 3762
rect 18873 3704 18878 3760
rect 18934 3704 24766 3760
rect 24822 3704 24827 3760
rect 18873 3702 24827 3704
rect 18873 3699 18939 3702
rect 24761 3699 24827 3702
rect 10277 3560 10597 3561
rect 10277 3496 10285 3560
rect 10349 3496 10365 3560
rect 10429 3496 10445 3560
rect 10509 3496 10525 3560
rect 10589 3496 10597 3560
rect 10277 3495 10597 3496
rect 19610 3560 19930 3561
rect 19610 3496 19618 3560
rect 19682 3496 19698 3560
rect 19762 3496 19778 3560
rect 19842 3496 19858 3560
rect 19922 3496 19930 3560
rect 19610 3495 19930 3496
rect 23933 3490 23999 3493
rect 27520 3490 28000 3520
rect 23933 3488 28000 3490
rect 23933 3432 23938 3488
rect 23994 3432 28000 3488
rect 23933 3430 28000 3432
rect 23933 3427 23999 3430
rect 27520 3400 28000 3430
rect 24761 3082 24827 3085
rect 26233 3082 26299 3085
rect 24761 3080 26299 3082
rect 24761 3024 24766 3080
rect 24822 3024 26238 3080
rect 26294 3024 26299 3080
rect 24761 3022 26299 3024
rect 24761 3019 24827 3022
rect 26233 3019 26299 3022
rect 5610 3016 5930 3017
rect 5610 2952 5618 3016
rect 5682 2952 5698 3016
rect 5762 2952 5778 3016
rect 5842 2952 5858 3016
rect 5922 2952 5930 3016
rect 5610 2951 5930 2952
rect 14944 3016 15264 3017
rect 14944 2952 14952 3016
rect 15016 2952 15032 3016
rect 15096 2952 15112 3016
rect 15176 2952 15192 3016
rect 15256 2952 15264 3016
rect 14944 2951 15264 2952
rect 24277 3016 24597 3017
rect 24277 2952 24285 3016
rect 24349 2952 24365 3016
rect 24429 2952 24445 3016
rect 24509 2952 24525 3016
rect 24589 2952 24597 3016
rect 24277 2951 24597 2952
rect 27520 2946 28000 2976
rect 24902 2886 28000 2946
rect 16757 2810 16823 2813
rect 24902 2810 24962 2886
rect 27520 2856 28000 2886
rect 16757 2808 24962 2810
rect 16757 2752 16762 2808
rect 16818 2752 24962 2808
rect 16757 2750 24962 2752
rect 16757 2747 16823 2750
rect 10277 2472 10597 2473
rect 10277 2408 10285 2472
rect 10349 2408 10365 2472
rect 10429 2408 10445 2472
rect 10509 2408 10525 2472
rect 10589 2408 10597 2472
rect 10277 2407 10597 2408
rect 19610 2472 19930 2473
rect 19610 2408 19618 2472
rect 19682 2408 19698 2472
rect 19762 2408 19778 2472
rect 19842 2408 19858 2472
rect 19922 2408 19930 2472
rect 19610 2407 19930 2408
rect 27520 2266 28000 2296
rect 24902 2206 28000 2266
rect 16665 2130 16731 2133
rect 24761 2130 24827 2133
rect 16665 2128 24827 2130
rect 16665 2072 16670 2128
rect 16726 2072 24766 2128
rect 24822 2072 24827 2128
rect 16665 2070 24827 2072
rect 16665 2067 16731 2070
rect 24761 2067 24827 2070
rect 5610 1928 5930 1929
rect 5610 1864 5618 1928
rect 5682 1864 5698 1928
rect 5762 1864 5778 1928
rect 5842 1864 5858 1928
rect 5922 1864 5930 1928
rect 5610 1863 5930 1864
rect 14944 1928 15264 1929
rect 14944 1864 14952 1928
rect 15016 1864 15032 1928
rect 15096 1864 15112 1928
rect 15176 1864 15192 1928
rect 15256 1864 15264 1928
rect 14944 1863 15264 1864
rect 24277 1928 24597 1929
rect 24277 1864 24285 1928
rect 24349 1864 24365 1928
rect 24429 1864 24445 1928
rect 24509 1864 24525 1928
rect 24589 1864 24597 1928
rect 24277 1863 24597 1864
rect 15837 1314 15903 1317
rect 24902 1314 24962 2206
rect 27520 2176 28000 2206
rect 25221 1722 25287 1725
rect 27520 1722 28000 1752
rect 25221 1720 28000 1722
rect 25221 1664 25226 1720
rect 25282 1664 28000 1720
rect 25221 1662 28000 1664
rect 25221 1659 25287 1662
rect 27520 1632 28000 1662
rect 15837 1312 24962 1314
rect 15837 1256 15842 1312
rect 15898 1256 24962 1312
rect 15837 1254 24962 1256
rect 15837 1251 15903 1254
rect 13261 1178 13327 1181
rect 27520 1178 28000 1208
rect 13261 1176 28000 1178
rect 13261 1120 13266 1176
rect 13322 1120 28000 1176
rect 13261 1118 28000 1120
rect 13261 1115 13327 1118
rect 27520 1088 28000 1118
rect 24669 634 24735 637
rect 27520 634 28000 664
rect 24669 632 28000 634
rect 24669 576 24674 632
rect 24730 576 28000 632
rect 24669 574 28000 576
rect 24669 571 24735 574
rect 27520 544 28000 574
rect 23565 90 23631 93
rect 27520 90 28000 120
rect 23565 88 28000 90
rect 23565 32 23570 88
rect 23626 32 28000 88
rect 23565 30 28000 32
rect 23565 27 23631 30
rect 27520 0 28000 30
<< via3 >>
rect 10285 25316 10349 25320
rect 10285 25260 10289 25316
rect 10289 25260 10345 25316
rect 10345 25260 10349 25316
rect 10285 25256 10349 25260
rect 10365 25316 10429 25320
rect 10365 25260 10369 25316
rect 10369 25260 10425 25316
rect 10425 25260 10429 25316
rect 10365 25256 10429 25260
rect 10445 25316 10509 25320
rect 10445 25260 10449 25316
rect 10449 25260 10505 25316
rect 10505 25260 10509 25316
rect 10445 25256 10509 25260
rect 10525 25316 10589 25320
rect 10525 25260 10529 25316
rect 10529 25260 10585 25316
rect 10585 25260 10589 25316
rect 10525 25256 10589 25260
rect 19618 25316 19682 25320
rect 19618 25260 19622 25316
rect 19622 25260 19678 25316
rect 19678 25260 19682 25316
rect 19618 25256 19682 25260
rect 19698 25316 19762 25320
rect 19698 25260 19702 25316
rect 19702 25260 19758 25316
rect 19758 25260 19762 25316
rect 19698 25256 19762 25260
rect 19778 25316 19842 25320
rect 19778 25260 19782 25316
rect 19782 25260 19838 25316
rect 19838 25260 19842 25316
rect 19778 25256 19842 25260
rect 19858 25316 19922 25320
rect 19858 25260 19862 25316
rect 19862 25260 19918 25316
rect 19918 25260 19922 25316
rect 19858 25256 19922 25260
rect 5618 24772 5682 24776
rect 5618 24716 5622 24772
rect 5622 24716 5678 24772
rect 5678 24716 5682 24772
rect 5618 24712 5682 24716
rect 5698 24772 5762 24776
rect 5698 24716 5702 24772
rect 5702 24716 5758 24772
rect 5758 24716 5762 24772
rect 5698 24712 5762 24716
rect 5778 24772 5842 24776
rect 5778 24716 5782 24772
rect 5782 24716 5838 24772
rect 5838 24716 5842 24772
rect 5778 24712 5842 24716
rect 5858 24772 5922 24776
rect 5858 24716 5862 24772
rect 5862 24716 5918 24772
rect 5918 24716 5922 24772
rect 5858 24712 5922 24716
rect 14952 24772 15016 24776
rect 14952 24716 14956 24772
rect 14956 24716 15012 24772
rect 15012 24716 15016 24772
rect 14952 24712 15016 24716
rect 15032 24772 15096 24776
rect 15032 24716 15036 24772
rect 15036 24716 15092 24772
rect 15092 24716 15096 24772
rect 15032 24712 15096 24716
rect 15112 24772 15176 24776
rect 15112 24716 15116 24772
rect 15116 24716 15172 24772
rect 15172 24716 15176 24772
rect 15112 24712 15176 24716
rect 15192 24772 15256 24776
rect 15192 24716 15196 24772
rect 15196 24716 15252 24772
rect 15252 24716 15256 24772
rect 15192 24712 15256 24716
rect 24285 24772 24349 24776
rect 24285 24716 24289 24772
rect 24289 24716 24345 24772
rect 24345 24716 24349 24772
rect 24285 24712 24349 24716
rect 24365 24772 24429 24776
rect 24365 24716 24369 24772
rect 24369 24716 24425 24772
rect 24425 24716 24429 24772
rect 24365 24712 24429 24716
rect 24445 24772 24509 24776
rect 24445 24716 24449 24772
rect 24449 24716 24505 24772
rect 24505 24716 24509 24772
rect 24445 24712 24509 24716
rect 24525 24772 24589 24776
rect 24525 24716 24529 24772
rect 24529 24716 24585 24772
rect 24585 24716 24589 24772
rect 24525 24712 24589 24716
rect 10285 24228 10349 24232
rect 10285 24172 10289 24228
rect 10289 24172 10345 24228
rect 10345 24172 10349 24228
rect 10285 24168 10349 24172
rect 10365 24228 10429 24232
rect 10365 24172 10369 24228
rect 10369 24172 10425 24228
rect 10425 24172 10429 24228
rect 10365 24168 10429 24172
rect 10445 24228 10509 24232
rect 10445 24172 10449 24228
rect 10449 24172 10505 24228
rect 10505 24172 10509 24228
rect 10445 24168 10509 24172
rect 10525 24228 10589 24232
rect 10525 24172 10529 24228
rect 10529 24172 10585 24228
rect 10585 24172 10589 24228
rect 10525 24168 10589 24172
rect 19618 24228 19682 24232
rect 19618 24172 19622 24228
rect 19622 24172 19678 24228
rect 19678 24172 19682 24228
rect 19618 24168 19682 24172
rect 19698 24228 19762 24232
rect 19698 24172 19702 24228
rect 19702 24172 19758 24228
rect 19758 24172 19762 24228
rect 19698 24168 19762 24172
rect 19778 24228 19842 24232
rect 19778 24172 19782 24228
rect 19782 24172 19838 24228
rect 19838 24172 19842 24228
rect 19778 24168 19842 24172
rect 19858 24228 19922 24232
rect 19858 24172 19862 24228
rect 19862 24172 19918 24228
rect 19918 24172 19922 24228
rect 19858 24168 19922 24172
rect 6132 23828 6196 23892
rect 5618 23684 5682 23688
rect 5618 23628 5622 23684
rect 5622 23628 5678 23684
rect 5678 23628 5682 23684
rect 5618 23624 5682 23628
rect 5698 23684 5762 23688
rect 5698 23628 5702 23684
rect 5702 23628 5758 23684
rect 5758 23628 5762 23684
rect 5698 23624 5762 23628
rect 5778 23684 5842 23688
rect 5778 23628 5782 23684
rect 5782 23628 5838 23684
rect 5838 23628 5842 23684
rect 5778 23624 5842 23628
rect 5858 23684 5922 23688
rect 5858 23628 5862 23684
rect 5862 23628 5918 23684
rect 5918 23628 5922 23684
rect 5858 23624 5922 23628
rect 14952 23684 15016 23688
rect 14952 23628 14956 23684
rect 14956 23628 15012 23684
rect 15012 23628 15016 23684
rect 14952 23624 15016 23628
rect 15032 23684 15096 23688
rect 15032 23628 15036 23684
rect 15036 23628 15092 23684
rect 15092 23628 15096 23684
rect 15032 23624 15096 23628
rect 15112 23684 15176 23688
rect 15112 23628 15116 23684
rect 15116 23628 15172 23684
rect 15172 23628 15176 23684
rect 15112 23624 15176 23628
rect 15192 23684 15256 23688
rect 15192 23628 15196 23684
rect 15196 23628 15252 23684
rect 15252 23628 15256 23684
rect 15192 23624 15256 23628
rect 24285 23684 24349 23688
rect 24285 23628 24289 23684
rect 24289 23628 24345 23684
rect 24345 23628 24349 23684
rect 24285 23624 24349 23628
rect 24365 23684 24429 23688
rect 24365 23628 24369 23684
rect 24369 23628 24425 23684
rect 24425 23628 24429 23684
rect 24365 23624 24429 23628
rect 24445 23684 24509 23688
rect 24445 23628 24449 23684
rect 24449 23628 24505 23684
rect 24505 23628 24509 23684
rect 24445 23624 24509 23628
rect 24525 23684 24589 23688
rect 24525 23628 24529 23684
rect 24529 23628 24585 23684
rect 24585 23628 24589 23684
rect 24525 23624 24589 23628
rect 10916 23208 10980 23212
rect 10916 23152 10966 23208
rect 10966 23152 10980 23208
rect 10916 23148 10980 23152
rect 10285 23140 10349 23144
rect 10285 23084 10289 23140
rect 10289 23084 10345 23140
rect 10345 23084 10349 23140
rect 10285 23080 10349 23084
rect 10365 23140 10429 23144
rect 10365 23084 10369 23140
rect 10369 23084 10425 23140
rect 10425 23084 10429 23140
rect 10365 23080 10429 23084
rect 10445 23140 10509 23144
rect 10445 23084 10449 23140
rect 10449 23084 10505 23140
rect 10505 23084 10509 23140
rect 10445 23080 10509 23084
rect 10525 23140 10589 23144
rect 10525 23084 10529 23140
rect 10529 23084 10585 23140
rect 10585 23084 10589 23140
rect 10525 23080 10589 23084
rect 19618 23140 19682 23144
rect 19618 23084 19622 23140
rect 19622 23084 19678 23140
rect 19678 23084 19682 23140
rect 19618 23080 19682 23084
rect 19698 23140 19762 23144
rect 19698 23084 19702 23140
rect 19702 23084 19758 23140
rect 19758 23084 19762 23140
rect 19698 23080 19762 23084
rect 19778 23140 19842 23144
rect 19778 23084 19782 23140
rect 19782 23084 19838 23140
rect 19838 23084 19842 23140
rect 19778 23080 19842 23084
rect 19858 23140 19922 23144
rect 19858 23084 19862 23140
rect 19862 23084 19918 23140
rect 19918 23084 19922 23140
rect 19858 23080 19922 23084
rect 5618 22596 5682 22600
rect 5618 22540 5622 22596
rect 5622 22540 5678 22596
rect 5678 22540 5682 22596
rect 5618 22536 5682 22540
rect 5698 22596 5762 22600
rect 5698 22540 5702 22596
rect 5702 22540 5758 22596
rect 5758 22540 5762 22596
rect 5698 22536 5762 22540
rect 5778 22596 5842 22600
rect 5778 22540 5782 22596
rect 5782 22540 5838 22596
rect 5838 22540 5842 22596
rect 5778 22536 5842 22540
rect 5858 22596 5922 22600
rect 5858 22540 5862 22596
rect 5862 22540 5918 22596
rect 5918 22540 5922 22596
rect 5858 22536 5922 22540
rect 14952 22596 15016 22600
rect 14952 22540 14956 22596
rect 14956 22540 15012 22596
rect 15012 22540 15016 22596
rect 14952 22536 15016 22540
rect 15032 22596 15096 22600
rect 15032 22540 15036 22596
rect 15036 22540 15092 22596
rect 15092 22540 15096 22596
rect 15032 22536 15096 22540
rect 15112 22596 15176 22600
rect 15112 22540 15116 22596
rect 15116 22540 15172 22596
rect 15172 22540 15176 22596
rect 15112 22536 15176 22540
rect 15192 22596 15256 22600
rect 15192 22540 15196 22596
rect 15196 22540 15252 22596
rect 15252 22540 15256 22596
rect 15192 22536 15256 22540
rect 24285 22596 24349 22600
rect 24285 22540 24289 22596
rect 24289 22540 24345 22596
rect 24345 22540 24349 22596
rect 24285 22536 24349 22540
rect 24365 22596 24429 22600
rect 24365 22540 24369 22596
rect 24369 22540 24425 22596
rect 24425 22540 24429 22596
rect 24365 22536 24429 22540
rect 24445 22596 24509 22600
rect 24445 22540 24449 22596
rect 24449 22540 24505 22596
rect 24505 22540 24509 22596
rect 24445 22536 24509 22540
rect 24525 22596 24589 22600
rect 24525 22540 24529 22596
rect 24529 22540 24585 22596
rect 24585 22540 24589 22596
rect 24525 22536 24589 22540
rect 10285 22052 10349 22056
rect 10285 21996 10289 22052
rect 10289 21996 10345 22052
rect 10345 21996 10349 22052
rect 10285 21992 10349 21996
rect 10365 22052 10429 22056
rect 10365 21996 10369 22052
rect 10369 21996 10425 22052
rect 10425 21996 10429 22052
rect 10365 21992 10429 21996
rect 10445 22052 10509 22056
rect 10445 21996 10449 22052
rect 10449 21996 10505 22052
rect 10505 21996 10509 22052
rect 10445 21992 10509 21996
rect 10525 22052 10589 22056
rect 10525 21996 10529 22052
rect 10529 21996 10585 22052
rect 10585 21996 10589 22052
rect 10525 21992 10589 21996
rect 19618 22052 19682 22056
rect 19618 21996 19622 22052
rect 19622 21996 19678 22052
rect 19678 21996 19682 22052
rect 19618 21992 19682 21996
rect 19698 22052 19762 22056
rect 19698 21996 19702 22052
rect 19702 21996 19758 22052
rect 19758 21996 19762 22052
rect 19698 21992 19762 21996
rect 19778 22052 19842 22056
rect 19778 21996 19782 22052
rect 19782 21996 19838 22052
rect 19838 21996 19842 22052
rect 19778 21992 19842 21996
rect 19858 22052 19922 22056
rect 19858 21996 19862 22052
rect 19862 21996 19918 22052
rect 19918 21996 19922 22052
rect 19858 21992 19922 21996
rect 5618 21508 5682 21512
rect 5618 21452 5622 21508
rect 5622 21452 5678 21508
rect 5678 21452 5682 21508
rect 5618 21448 5682 21452
rect 5698 21508 5762 21512
rect 5698 21452 5702 21508
rect 5702 21452 5758 21508
rect 5758 21452 5762 21508
rect 5698 21448 5762 21452
rect 5778 21508 5842 21512
rect 5778 21452 5782 21508
rect 5782 21452 5838 21508
rect 5838 21452 5842 21508
rect 5778 21448 5842 21452
rect 5858 21508 5922 21512
rect 5858 21452 5862 21508
rect 5862 21452 5918 21508
rect 5918 21452 5922 21508
rect 5858 21448 5922 21452
rect 14952 21508 15016 21512
rect 14952 21452 14956 21508
rect 14956 21452 15012 21508
rect 15012 21452 15016 21508
rect 14952 21448 15016 21452
rect 15032 21508 15096 21512
rect 15032 21452 15036 21508
rect 15036 21452 15092 21508
rect 15092 21452 15096 21508
rect 15032 21448 15096 21452
rect 15112 21508 15176 21512
rect 15112 21452 15116 21508
rect 15116 21452 15172 21508
rect 15172 21452 15176 21508
rect 15112 21448 15176 21452
rect 15192 21508 15256 21512
rect 15192 21452 15196 21508
rect 15196 21452 15252 21508
rect 15252 21452 15256 21508
rect 15192 21448 15256 21452
rect 24285 21508 24349 21512
rect 24285 21452 24289 21508
rect 24289 21452 24345 21508
rect 24345 21452 24349 21508
rect 24285 21448 24349 21452
rect 24365 21508 24429 21512
rect 24365 21452 24369 21508
rect 24369 21452 24425 21508
rect 24425 21452 24429 21508
rect 24365 21448 24429 21452
rect 24445 21508 24509 21512
rect 24445 21452 24449 21508
rect 24449 21452 24505 21508
rect 24505 21452 24509 21508
rect 24445 21448 24509 21452
rect 24525 21508 24589 21512
rect 24525 21452 24529 21508
rect 24529 21452 24585 21508
rect 24585 21452 24589 21508
rect 24525 21448 24589 21452
rect 10285 20964 10349 20968
rect 10285 20908 10289 20964
rect 10289 20908 10345 20964
rect 10345 20908 10349 20964
rect 10285 20904 10349 20908
rect 10365 20964 10429 20968
rect 10365 20908 10369 20964
rect 10369 20908 10425 20964
rect 10425 20908 10429 20964
rect 10365 20904 10429 20908
rect 10445 20964 10509 20968
rect 10445 20908 10449 20964
rect 10449 20908 10505 20964
rect 10505 20908 10509 20964
rect 10445 20904 10509 20908
rect 10525 20964 10589 20968
rect 10525 20908 10529 20964
rect 10529 20908 10585 20964
rect 10585 20908 10589 20964
rect 10525 20904 10589 20908
rect 19618 20964 19682 20968
rect 19618 20908 19622 20964
rect 19622 20908 19678 20964
rect 19678 20908 19682 20964
rect 19618 20904 19682 20908
rect 19698 20964 19762 20968
rect 19698 20908 19702 20964
rect 19702 20908 19758 20964
rect 19758 20908 19762 20964
rect 19698 20904 19762 20908
rect 19778 20964 19842 20968
rect 19778 20908 19782 20964
rect 19782 20908 19838 20964
rect 19838 20908 19842 20964
rect 19778 20904 19842 20908
rect 19858 20964 19922 20968
rect 19858 20908 19862 20964
rect 19862 20908 19918 20964
rect 19918 20908 19922 20964
rect 19858 20904 19922 20908
rect 21220 20836 21284 20900
rect 23980 20564 24044 20628
rect 5618 20420 5682 20424
rect 5618 20364 5622 20420
rect 5622 20364 5678 20420
rect 5678 20364 5682 20420
rect 5618 20360 5682 20364
rect 5698 20420 5762 20424
rect 5698 20364 5702 20420
rect 5702 20364 5758 20420
rect 5758 20364 5762 20420
rect 5698 20360 5762 20364
rect 5778 20420 5842 20424
rect 5778 20364 5782 20420
rect 5782 20364 5838 20420
rect 5838 20364 5842 20420
rect 5778 20360 5842 20364
rect 5858 20420 5922 20424
rect 5858 20364 5862 20420
rect 5862 20364 5918 20420
rect 5918 20364 5922 20420
rect 5858 20360 5922 20364
rect 14952 20420 15016 20424
rect 14952 20364 14956 20420
rect 14956 20364 15012 20420
rect 15012 20364 15016 20420
rect 14952 20360 15016 20364
rect 15032 20420 15096 20424
rect 15032 20364 15036 20420
rect 15036 20364 15092 20420
rect 15092 20364 15096 20420
rect 15032 20360 15096 20364
rect 15112 20420 15176 20424
rect 15112 20364 15116 20420
rect 15116 20364 15172 20420
rect 15172 20364 15176 20420
rect 15112 20360 15176 20364
rect 15192 20420 15256 20424
rect 15192 20364 15196 20420
rect 15196 20364 15252 20420
rect 15252 20364 15256 20420
rect 15192 20360 15256 20364
rect 24285 20420 24349 20424
rect 24285 20364 24289 20420
rect 24289 20364 24345 20420
rect 24345 20364 24349 20420
rect 24285 20360 24349 20364
rect 24365 20420 24429 20424
rect 24365 20364 24369 20420
rect 24369 20364 24425 20420
rect 24425 20364 24429 20420
rect 24365 20360 24429 20364
rect 24445 20420 24509 20424
rect 24445 20364 24449 20420
rect 24449 20364 24505 20420
rect 24505 20364 24509 20420
rect 24445 20360 24509 20364
rect 24525 20420 24589 20424
rect 24525 20364 24529 20420
rect 24529 20364 24585 20420
rect 24585 20364 24589 20420
rect 24525 20360 24589 20364
rect 10285 19876 10349 19880
rect 10285 19820 10289 19876
rect 10289 19820 10345 19876
rect 10345 19820 10349 19876
rect 10285 19816 10349 19820
rect 10365 19876 10429 19880
rect 10365 19820 10369 19876
rect 10369 19820 10425 19876
rect 10425 19820 10429 19876
rect 10365 19816 10429 19820
rect 10445 19876 10509 19880
rect 10445 19820 10449 19876
rect 10449 19820 10505 19876
rect 10505 19820 10509 19876
rect 10445 19816 10509 19820
rect 10525 19876 10589 19880
rect 10525 19820 10529 19876
rect 10529 19820 10585 19876
rect 10585 19820 10589 19876
rect 10525 19816 10589 19820
rect 19618 19876 19682 19880
rect 19618 19820 19622 19876
rect 19622 19820 19678 19876
rect 19678 19820 19682 19876
rect 19618 19816 19682 19820
rect 19698 19876 19762 19880
rect 19698 19820 19702 19876
rect 19702 19820 19758 19876
rect 19758 19820 19762 19876
rect 19698 19816 19762 19820
rect 19778 19876 19842 19880
rect 19778 19820 19782 19876
rect 19782 19820 19838 19876
rect 19838 19820 19842 19876
rect 19778 19816 19842 19820
rect 19858 19876 19922 19880
rect 19858 19820 19862 19876
rect 19862 19820 19918 19876
rect 19918 19820 19922 19876
rect 19858 19816 19922 19820
rect 5618 19332 5682 19336
rect 5618 19276 5622 19332
rect 5622 19276 5678 19332
rect 5678 19276 5682 19332
rect 5618 19272 5682 19276
rect 5698 19332 5762 19336
rect 5698 19276 5702 19332
rect 5702 19276 5758 19332
rect 5758 19276 5762 19332
rect 5698 19272 5762 19276
rect 5778 19332 5842 19336
rect 5778 19276 5782 19332
rect 5782 19276 5838 19332
rect 5838 19276 5842 19332
rect 5778 19272 5842 19276
rect 5858 19332 5922 19336
rect 5858 19276 5862 19332
rect 5862 19276 5918 19332
rect 5918 19276 5922 19332
rect 5858 19272 5922 19276
rect 14952 19332 15016 19336
rect 14952 19276 14956 19332
rect 14956 19276 15012 19332
rect 15012 19276 15016 19332
rect 14952 19272 15016 19276
rect 15032 19332 15096 19336
rect 15032 19276 15036 19332
rect 15036 19276 15092 19332
rect 15092 19276 15096 19332
rect 15032 19272 15096 19276
rect 15112 19332 15176 19336
rect 15112 19276 15116 19332
rect 15116 19276 15172 19332
rect 15172 19276 15176 19332
rect 15112 19272 15176 19276
rect 15192 19332 15256 19336
rect 15192 19276 15196 19332
rect 15196 19276 15252 19332
rect 15252 19276 15256 19332
rect 15192 19272 15256 19276
rect 24285 19332 24349 19336
rect 24285 19276 24289 19332
rect 24289 19276 24345 19332
rect 24345 19276 24349 19332
rect 24285 19272 24349 19276
rect 24365 19332 24429 19336
rect 24365 19276 24369 19332
rect 24369 19276 24425 19332
rect 24425 19276 24429 19332
rect 24365 19272 24429 19276
rect 24445 19332 24509 19336
rect 24445 19276 24449 19332
rect 24449 19276 24505 19332
rect 24505 19276 24509 19332
rect 24445 19272 24509 19276
rect 24525 19332 24589 19336
rect 24525 19276 24529 19332
rect 24529 19276 24585 19332
rect 24585 19276 24589 19332
rect 24525 19272 24589 19276
rect 10285 18788 10349 18792
rect 10285 18732 10289 18788
rect 10289 18732 10345 18788
rect 10345 18732 10349 18788
rect 10285 18728 10349 18732
rect 10365 18788 10429 18792
rect 10365 18732 10369 18788
rect 10369 18732 10425 18788
rect 10425 18732 10429 18788
rect 10365 18728 10429 18732
rect 10445 18788 10509 18792
rect 10445 18732 10449 18788
rect 10449 18732 10505 18788
rect 10505 18732 10509 18788
rect 10445 18728 10509 18732
rect 10525 18788 10589 18792
rect 10525 18732 10529 18788
rect 10529 18732 10585 18788
rect 10585 18732 10589 18788
rect 10525 18728 10589 18732
rect 19618 18788 19682 18792
rect 19618 18732 19622 18788
rect 19622 18732 19678 18788
rect 19678 18732 19682 18788
rect 19618 18728 19682 18732
rect 19698 18788 19762 18792
rect 19698 18732 19702 18788
rect 19702 18732 19758 18788
rect 19758 18732 19762 18788
rect 19698 18728 19762 18732
rect 19778 18788 19842 18792
rect 19778 18732 19782 18788
rect 19782 18732 19838 18788
rect 19838 18732 19842 18788
rect 19778 18728 19842 18732
rect 19858 18788 19922 18792
rect 19858 18732 19862 18788
rect 19862 18732 19918 18788
rect 19918 18732 19922 18788
rect 19858 18728 19922 18732
rect 5618 18244 5682 18248
rect 5618 18188 5622 18244
rect 5622 18188 5678 18244
rect 5678 18188 5682 18244
rect 5618 18184 5682 18188
rect 5698 18244 5762 18248
rect 5698 18188 5702 18244
rect 5702 18188 5758 18244
rect 5758 18188 5762 18244
rect 5698 18184 5762 18188
rect 5778 18244 5842 18248
rect 5778 18188 5782 18244
rect 5782 18188 5838 18244
rect 5838 18188 5842 18244
rect 5778 18184 5842 18188
rect 5858 18244 5922 18248
rect 5858 18188 5862 18244
rect 5862 18188 5918 18244
rect 5918 18188 5922 18244
rect 5858 18184 5922 18188
rect 14952 18244 15016 18248
rect 14952 18188 14956 18244
rect 14956 18188 15012 18244
rect 15012 18188 15016 18244
rect 14952 18184 15016 18188
rect 15032 18244 15096 18248
rect 15032 18188 15036 18244
rect 15036 18188 15092 18244
rect 15092 18188 15096 18244
rect 15032 18184 15096 18188
rect 15112 18244 15176 18248
rect 15112 18188 15116 18244
rect 15116 18188 15172 18244
rect 15172 18188 15176 18244
rect 15112 18184 15176 18188
rect 15192 18244 15256 18248
rect 15192 18188 15196 18244
rect 15196 18188 15252 18244
rect 15252 18188 15256 18244
rect 15192 18184 15256 18188
rect 24285 18244 24349 18248
rect 24285 18188 24289 18244
rect 24289 18188 24345 18244
rect 24345 18188 24349 18244
rect 24285 18184 24349 18188
rect 24365 18244 24429 18248
rect 24365 18188 24369 18244
rect 24369 18188 24425 18244
rect 24425 18188 24429 18244
rect 24365 18184 24429 18188
rect 24445 18244 24509 18248
rect 24445 18188 24449 18244
rect 24449 18188 24505 18244
rect 24505 18188 24509 18244
rect 24445 18184 24509 18188
rect 24525 18244 24589 18248
rect 24525 18188 24529 18244
rect 24529 18188 24585 18244
rect 24585 18188 24589 18244
rect 24525 18184 24589 18188
rect 10285 17700 10349 17704
rect 10285 17644 10289 17700
rect 10289 17644 10345 17700
rect 10345 17644 10349 17700
rect 10285 17640 10349 17644
rect 10365 17700 10429 17704
rect 10365 17644 10369 17700
rect 10369 17644 10425 17700
rect 10425 17644 10429 17700
rect 10365 17640 10429 17644
rect 10445 17700 10509 17704
rect 10445 17644 10449 17700
rect 10449 17644 10505 17700
rect 10505 17644 10509 17700
rect 10445 17640 10509 17644
rect 10525 17700 10589 17704
rect 10525 17644 10529 17700
rect 10529 17644 10585 17700
rect 10585 17644 10589 17700
rect 10525 17640 10589 17644
rect 19618 17700 19682 17704
rect 19618 17644 19622 17700
rect 19622 17644 19678 17700
rect 19678 17644 19682 17700
rect 19618 17640 19682 17644
rect 19698 17700 19762 17704
rect 19698 17644 19702 17700
rect 19702 17644 19758 17700
rect 19758 17644 19762 17700
rect 19698 17640 19762 17644
rect 19778 17700 19842 17704
rect 19778 17644 19782 17700
rect 19782 17644 19838 17700
rect 19838 17644 19842 17700
rect 19778 17640 19842 17644
rect 19858 17700 19922 17704
rect 19858 17644 19862 17700
rect 19862 17644 19918 17700
rect 19918 17644 19922 17700
rect 19858 17640 19922 17644
rect 5618 17156 5682 17160
rect 5618 17100 5622 17156
rect 5622 17100 5678 17156
rect 5678 17100 5682 17156
rect 5618 17096 5682 17100
rect 5698 17156 5762 17160
rect 5698 17100 5702 17156
rect 5702 17100 5758 17156
rect 5758 17100 5762 17156
rect 5698 17096 5762 17100
rect 5778 17156 5842 17160
rect 5778 17100 5782 17156
rect 5782 17100 5838 17156
rect 5838 17100 5842 17156
rect 5778 17096 5842 17100
rect 5858 17156 5922 17160
rect 5858 17100 5862 17156
rect 5862 17100 5918 17156
rect 5918 17100 5922 17156
rect 5858 17096 5922 17100
rect 14952 17156 15016 17160
rect 14952 17100 14956 17156
rect 14956 17100 15012 17156
rect 15012 17100 15016 17156
rect 14952 17096 15016 17100
rect 15032 17156 15096 17160
rect 15032 17100 15036 17156
rect 15036 17100 15092 17156
rect 15092 17100 15096 17156
rect 15032 17096 15096 17100
rect 15112 17156 15176 17160
rect 15112 17100 15116 17156
rect 15116 17100 15172 17156
rect 15172 17100 15176 17156
rect 15112 17096 15176 17100
rect 15192 17156 15256 17160
rect 15192 17100 15196 17156
rect 15196 17100 15252 17156
rect 15252 17100 15256 17156
rect 15192 17096 15256 17100
rect 24285 17156 24349 17160
rect 24285 17100 24289 17156
rect 24289 17100 24345 17156
rect 24345 17100 24349 17156
rect 24285 17096 24349 17100
rect 24365 17156 24429 17160
rect 24365 17100 24369 17156
rect 24369 17100 24425 17156
rect 24425 17100 24429 17156
rect 24365 17096 24429 17100
rect 24445 17156 24509 17160
rect 24445 17100 24449 17156
rect 24449 17100 24505 17156
rect 24505 17100 24509 17156
rect 24445 17096 24509 17100
rect 24525 17156 24589 17160
rect 24525 17100 24529 17156
rect 24529 17100 24585 17156
rect 24585 17100 24589 17156
rect 24525 17096 24589 17100
rect 10285 16612 10349 16616
rect 10285 16556 10289 16612
rect 10289 16556 10345 16612
rect 10345 16556 10349 16612
rect 10285 16552 10349 16556
rect 10365 16612 10429 16616
rect 10365 16556 10369 16612
rect 10369 16556 10425 16612
rect 10425 16556 10429 16612
rect 10365 16552 10429 16556
rect 10445 16612 10509 16616
rect 10445 16556 10449 16612
rect 10449 16556 10505 16612
rect 10505 16556 10509 16612
rect 10445 16552 10509 16556
rect 10525 16612 10589 16616
rect 10525 16556 10529 16612
rect 10529 16556 10585 16612
rect 10585 16556 10589 16612
rect 10525 16552 10589 16556
rect 19618 16612 19682 16616
rect 19618 16556 19622 16612
rect 19622 16556 19678 16612
rect 19678 16556 19682 16612
rect 19618 16552 19682 16556
rect 19698 16612 19762 16616
rect 19698 16556 19702 16612
rect 19702 16556 19758 16612
rect 19758 16556 19762 16612
rect 19698 16552 19762 16556
rect 19778 16612 19842 16616
rect 19778 16556 19782 16612
rect 19782 16556 19838 16612
rect 19838 16556 19842 16612
rect 19778 16552 19842 16556
rect 19858 16612 19922 16616
rect 19858 16556 19862 16612
rect 19862 16556 19918 16612
rect 19918 16556 19922 16612
rect 19858 16552 19922 16556
rect 5618 16068 5682 16072
rect 5618 16012 5622 16068
rect 5622 16012 5678 16068
rect 5678 16012 5682 16068
rect 5618 16008 5682 16012
rect 5698 16068 5762 16072
rect 5698 16012 5702 16068
rect 5702 16012 5758 16068
rect 5758 16012 5762 16068
rect 5698 16008 5762 16012
rect 5778 16068 5842 16072
rect 5778 16012 5782 16068
rect 5782 16012 5838 16068
rect 5838 16012 5842 16068
rect 5778 16008 5842 16012
rect 5858 16068 5922 16072
rect 5858 16012 5862 16068
rect 5862 16012 5918 16068
rect 5918 16012 5922 16068
rect 5858 16008 5922 16012
rect 14952 16068 15016 16072
rect 14952 16012 14956 16068
rect 14956 16012 15012 16068
rect 15012 16012 15016 16068
rect 14952 16008 15016 16012
rect 15032 16068 15096 16072
rect 15032 16012 15036 16068
rect 15036 16012 15092 16068
rect 15092 16012 15096 16068
rect 15032 16008 15096 16012
rect 15112 16068 15176 16072
rect 15112 16012 15116 16068
rect 15116 16012 15172 16068
rect 15172 16012 15176 16068
rect 15112 16008 15176 16012
rect 15192 16068 15256 16072
rect 15192 16012 15196 16068
rect 15196 16012 15252 16068
rect 15252 16012 15256 16068
rect 15192 16008 15256 16012
rect 24285 16068 24349 16072
rect 24285 16012 24289 16068
rect 24289 16012 24345 16068
rect 24345 16012 24349 16068
rect 24285 16008 24349 16012
rect 24365 16068 24429 16072
rect 24365 16012 24369 16068
rect 24369 16012 24425 16068
rect 24425 16012 24429 16068
rect 24365 16008 24429 16012
rect 24445 16068 24509 16072
rect 24445 16012 24449 16068
rect 24449 16012 24505 16068
rect 24505 16012 24509 16068
rect 24445 16008 24509 16012
rect 24525 16068 24589 16072
rect 24525 16012 24529 16068
rect 24529 16012 24585 16068
rect 24585 16012 24589 16068
rect 24525 16008 24589 16012
rect 10285 15524 10349 15528
rect 10285 15468 10289 15524
rect 10289 15468 10345 15524
rect 10345 15468 10349 15524
rect 10285 15464 10349 15468
rect 10365 15524 10429 15528
rect 10365 15468 10369 15524
rect 10369 15468 10425 15524
rect 10425 15468 10429 15524
rect 10365 15464 10429 15468
rect 10445 15524 10509 15528
rect 10445 15468 10449 15524
rect 10449 15468 10505 15524
rect 10505 15468 10509 15524
rect 10445 15464 10509 15468
rect 10525 15524 10589 15528
rect 10525 15468 10529 15524
rect 10529 15468 10585 15524
rect 10585 15468 10589 15524
rect 10525 15464 10589 15468
rect 19618 15524 19682 15528
rect 19618 15468 19622 15524
rect 19622 15468 19678 15524
rect 19678 15468 19682 15524
rect 19618 15464 19682 15468
rect 19698 15524 19762 15528
rect 19698 15468 19702 15524
rect 19702 15468 19758 15524
rect 19758 15468 19762 15524
rect 19698 15464 19762 15468
rect 19778 15524 19842 15528
rect 19778 15468 19782 15524
rect 19782 15468 19838 15524
rect 19838 15468 19842 15524
rect 19778 15464 19842 15468
rect 19858 15524 19922 15528
rect 19858 15468 19862 15524
rect 19862 15468 19918 15524
rect 19918 15468 19922 15524
rect 19858 15464 19922 15468
rect 5618 14980 5682 14984
rect 5618 14924 5622 14980
rect 5622 14924 5678 14980
rect 5678 14924 5682 14980
rect 5618 14920 5682 14924
rect 5698 14980 5762 14984
rect 5698 14924 5702 14980
rect 5702 14924 5758 14980
rect 5758 14924 5762 14980
rect 5698 14920 5762 14924
rect 5778 14980 5842 14984
rect 5778 14924 5782 14980
rect 5782 14924 5838 14980
rect 5838 14924 5842 14980
rect 5778 14920 5842 14924
rect 5858 14980 5922 14984
rect 5858 14924 5862 14980
rect 5862 14924 5918 14980
rect 5918 14924 5922 14980
rect 5858 14920 5922 14924
rect 14952 14980 15016 14984
rect 14952 14924 14956 14980
rect 14956 14924 15012 14980
rect 15012 14924 15016 14980
rect 14952 14920 15016 14924
rect 15032 14980 15096 14984
rect 15032 14924 15036 14980
rect 15036 14924 15092 14980
rect 15092 14924 15096 14980
rect 15032 14920 15096 14924
rect 15112 14980 15176 14984
rect 15112 14924 15116 14980
rect 15116 14924 15172 14980
rect 15172 14924 15176 14980
rect 15112 14920 15176 14924
rect 15192 14980 15256 14984
rect 15192 14924 15196 14980
rect 15196 14924 15252 14980
rect 15252 14924 15256 14980
rect 15192 14920 15256 14924
rect 24285 14980 24349 14984
rect 24285 14924 24289 14980
rect 24289 14924 24345 14980
rect 24345 14924 24349 14980
rect 24285 14920 24349 14924
rect 24365 14980 24429 14984
rect 24365 14924 24369 14980
rect 24369 14924 24425 14980
rect 24425 14924 24429 14980
rect 24365 14920 24429 14924
rect 24445 14980 24509 14984
rect 24445 14924 24449 14980
rect 24449 14924 24505 14980
rect 24505 14924 24509 14980
rect 24445 14920 24509 14924
rect 24525 14980 24589 14984
rect 24525 14924 24529 14980
rect 24529 14924 24585 14980
rect 24585 14924 24589 14980
rect 24525 14920 24589 14924
rect 10285 14436 10349 14440
rect 10285 14380 10289 14436
rect 10289 14380 10345 14436
rect 10345 14380 10349 14436
rect 10285 14376 10349 14380
rect 10365 14436 10429 14440
rect 10365 14380 10369 14436
rect 10369 14380 10425 14436
rect 10425 14380 10429 14436
rect 10365 14376 10429 14380
rect 10445 14436 10509 14440
rect 10445 14380 10449 14436
rect 10449 14380 10505 14436
rect 10505 14380 10509 14436
rect 10445 14376 10509 14380
rect 10525 14436 10589 14440
rect 10525 14380 10529 14436
rect 10529 14380 10585 14436
rect 10585 14380 10589 14436
rect 10525 14376 10589 14380
rect 19618 14436 19682 14440
rect 19618 14380 19622 14436
rect 19622 14380 19678 14436
rect 19678 14380 19682 14436
rect 19618 14376 19682 14380
rect 19698 14436 19762 14440
rect 19698 14380 19702 14436
rect 19702 14380 19758 14436
rect 19758 14380 19762 14436
rect 19698 14376 19762 14380
rect 19778 14436 19842 14440
rect 19778 14380 19782 14436
rect 19782 14380 19838 14436
rect 19838 14380 19842 14436
rect 19778 14376 19842 14380
rect 19858 14436 19922 14440
rect 19858 14380 19862 14436
rect 19862 14380 19918 14436
rect 19918 14380 19922 14436
rect 19858 14376 19922 14380
rect 5618 13892 5682 13896
rect 5618 13836 5622 13892
rect 5622 13836 5678 13892
rect 5678 13836 5682 13892
rect 5618 13832 5682 13836
rect 5698 13892 5762 13896
rect 5698 13836 5702 13892
rect 5702 13836 5758 13892
rect 5758 13836 5762 13892
rect 5698 13832 5762 13836
rect 5778 13892 5842 13896
rect 5778 13836 5782 13892
rect 5782 13836 5838 13892
rect 5838 13836 5842 13892
rect 5778 13832 5842 13836
rect 5858 13892 5922 13896
rect 5858 13836 5862 13892
rect 5862 13836 5918 13892
rect 5918 13836 5922 13892
rect 5858 13832 5922 13836
rect 14952 13892 15016 13896
rect 14952 13836 14956 13892
rect 14956 13836 15012 13892
rect 15012 13836 15016 13892
rect 14952 13832 15016 13836
rect 15032 13892 15096 13896
rect 15032 13836 15036 13892
rect 15036 13836 15092 13892
rect 15092 13836 15096 13892
rect 15032 13832 15096 13836
rect 15112 13892 15176 13896
rect 15112 13836 15116 13892
rect 15116 13836 15172 13892
rect 15172 13836 15176 13892
rect 15112 13832 15176 13836
rect 15192 13892 15256 13896
rect 15192 13836 15196 13892
rect 15196 13836 15252 13892
rect 15252 13836 15256 13892
rect 15192 13832 15256 13836
rect 24285 13892 24349 13896
rect 24285 13836 24289 13892
rect 24289 13836 24345 13892
rect 24345 13836 24349 13892
rect 24285 13832 24349 13836
rect 24365 13892 24429 13896
rect 24365 13836 24369 13892
rect 24369 13836 24425 13892
rect 24425 13836 24429 13892
rect 24365 13832 24429 13836
rect 24445 13892 24509 13896
rect 24445 13836 24449 13892
rect 24449 13836 24505 13892
rect 24505 13836 24509 13892
rect 24445 13832 24509 13836
rect 24525 13892 24589 13896
rect 24525 13836 24529 13892
rect 24529 13836 24585 13892
rect 24585 13836 24589 13892
rect 24525 13832 24589 13836
rect 10285 13348 10349 13352
rect 10285 13292 10289 13348
rect 10289 13292 10345 13348
rect 10345 13292 10349 13348
rect 10285 13288 10349 13292
rect 10365 13348 10429 13352
rect 10365 13292 10369 13348
rect 10369 13292 10425 13348
rect 10425 13292 10429 13348
rect 10365 13288 10429 13292
rect 10445 13348 10509 13352
rect 10445 13292 10449 13348
rect 10449 13292 10505 13348
rect 10505 13292 10509 13348
rect 10445 13288 10509 13292
rect 10525 13348 10589 13352
rect 10525 13292 10529 13348
rect 10529 13292 10585 13348
rect 10585 13292 10589 13348
rect 10525 13288 10589 13292
rect 19618 13348 19682 13352
rect 19618 13292 19622 13348
rect 19622 13292 19678 13348
rect 19678 13292 19682 13348
rect 19618 13288 19682 13292
rect 19698 13348 19762 13352
rect 19698 13292 19702 13348
rect 19702 13292 19758 13348
rect 19758 13292 19762 13348
rect 19698 13288 19762 13292
rect 19778 13348 19842 13352
rect 19778 13292 19782 13348
rect 19782 13292 19838 13348
rect 19838 13292 19842 13348
rect 19778 13288 19842 13292
rect 19858 13348 19922 13352
rect 19858 13292 19862 13348
rect 19862 13292 19918 13348
rect 19918 13292 19922 13348
rect 19858 13288 19922 13292
rect 5618 12804 5682 12808
rect 5618 12748 5622 12804
rect 5622 12748 5678 12804
rect 5678 12748 5682 12804
rect 5618 12744 5682 12748
rect 5698 12804 5762 12808
rect 5698 12748 5702 12804
rect 5702 12748 5758 12804
rect 5758 12748 5762 12804
rect 5698 12744 5762 12748
rect 5778 12804 5842 12808
rect 5778 12748 5782 12804
rect 5782 12748 5838 12804
rect 5838 12748 5842 12804
rect 5778 12744 5842 12748
rect 5858 12804 5922 12808
rect 5858 12748 5862 12804
rect 5862 12748 5918 12804
rect 5918 12748 5922 12804
rect 5858 12744 5922 12748
rect 14952 12804 15016 12808
rect 14952 12748 14956 12804
rect 14956 12748 15012 12804
rect 15012 12748 15016 12804
rect 14952 12744 15016 12748
rect 15032 12804 15096 12808
rect 15032 12748 15036 12804
rect 15036 12748 15092 12804
rect 15092 12748 15096 12804
rect 15032 12744 15096 12748
rect 15112 12804 15176 12808
rect 15112 12748 15116 12804
rect 15116 12748 15172 12804
rect 15172 12748 15176 12804
rect 15112 12744 15176 12748
rect 15192 12804 15256 12808
rect 15192 12748 15196 12804
rect 15196 12748 15252 12804
rect 15252 12748 15256 12804
rect 15192 12744 15256 12748
rect 24285 12804 24349 12808
rect 24285 12748 24289 12804
rect 24289 12748 24345 12804
rect 24345 12748 24349 12804
rect 24285 12744 24349 12748
rect 24365 12804 24429 12808
rect 24365 12748 24369 12804
rect 24369 12748 24425 12804
rect 24425 12748 24429 12804
rect 24365 12744 24429 12748
rect 24445 12804 24509 12808
rect 24445 12748 24449 12804
rect 24449 12748 24505 12804
rect 24505 12748 24509 12804
rect 24445 12744 24509 12748
rect 24525 12804 24589 12808
rect 24525 12748 24529 12804
rect 24529 12748 24585 12804
rect 24585 12748 24589 12804
rect 24525 12744 24589 12748
rect 10285 12260 10349 12264
rect 10285 12204 10289 12260
rect 10289 12204 10345 12260
rect 10345 12204 10349 12260
rect 10285 12200 10349 12204
rect 10365 12260 10429 12264
rect 10365 12204 10369 12260
rect 10369 12204 10425 12260
rect 10425 12204 10429 12260
rect 10365 12200 10429 12204
rect 10445 12260 10509 12264
rect 10445 12204 10449 12260
rect 10449 12204 10505 12260
rect 10505 12204 10509 12260
rect 10445 12200 10509 12204
rect 10525 12260 10589 12264
rect 10525 12204 10529 12260
rect 10529 12204 10585 12260
rect 10585 12204 10589 12260
rect 10525 12200 10589 12204
rect 19618 12260 19682 12264
rect 19618 12204 19622 12260
rect 19622 12204 19678 12260
rect 19678 12204 19682 12260
rect 19618 12200 19682 12204
rect 19698 12260 19762 12264
rect 19698 12204 19702 12260
rect 19702 12204 19758 12260
rect 19758 12204 19762 12260
rect 19698 12200 19762 12204
rect 19778 12260 19842 12264
rect 19778 12204 19782 12260
rect 19782 12204 19838 12260
rect 19838 12204 19842 12260
rect 19778 12200 19842 12204
rect 19858 12260 19922 12264
rect 19858 12204 19862 12260
rect 19862 12204 19918 12260
rect 19918 12204 19922 12260
rect 19858 12200 19922 12204
rect 5618 11716 5682 11720
rect 5618 11660 5622 11716
rect 5622 11660 5678 11716
rect 5678 11660 5682 11716
rect 5618 11656 5682 11660
rect 5698 11716 5762 11720
rect 5698 11660 5702 11716
rect 5702 11660 5758 11716
rect 5758 11660 5762 11716
rect 5698 11656 5762 11660
rect 5778 11716 5842 11720
rect 5778 11660 5782 11716
rect 5782 11660 5838 11716
rect 5838 11660 5842 11716
rect 5778 11656 5842 11660
rect 5858 11716 5922 11720
rect 5858 11660 5862 11716
rect 5862 11660 5918 11716
rect 5918 11660 5922 11716
rect 5858 11656 5922 11660
rect 14952 11716 15016 11720
rect 14952 11660 14956 11716
rect 14956 11660 15012 11716
rect 15012 11660 15016 11716
rect 14952 11656 15016 11660
rect 15032 11716 15096 11720
rect 15032 11660 15036 11716
rect 15036 11660 15092 11716
rect 15092 11660 15096 11716
rect 15032 11656 15096 11660
rect 15112 11716 15176 11720
rect 15112 11660 15116 11716
rect 15116 11660 15172 11716
rect 15172 11660 15176 11716
rect 15112 11656 15176 11660
rect 15192 11716 15256 11720
rect 15192 11660 15196 11716
rect 15196 11660 15252 11716
rect 15252 11660 15256 11716
rect 15192 11656 15256 11660
rect 24285 11716 24349 11720
rect 24285 11660 24289 11716
rect 24289 11660 24345 11716
rect 24345 11660 24349 11716
rect 24285 11656 24349 11660
rect 24365 11716 24429 11720
rect 24365 11660 24369 11716
rect 24369 11660 24425 11716
rect 24425 11660 24429 11716
rect 24365 11656 24429 11660
rect 24445 11716 24509 11720
rect 24445 11660 24449 11716
rect 24449 11660 24505 11716
rect 24505 11660 24509 11716
rect 24445 11656 24509 11660
rect 24525 11716 24589 11720
rect 24525 11660 24529 11716
rect 24529 11660 24585 11716
rect 24585 11660 24589 11716
rect 24525 11656 24589 11660
rect 10285 11172 10349 11176
rect 10285 11116 10289 11172
rect 10289 11116 10345 11172
rect 10345 11116 10349 11172
rect 10285 11112 10349 11116
rect 10365 11172 10429 11176
rect 10365 11116 10369 11172
rect 10369 11116 10425 11172
rect 10425 11116 10429 11172
rect 10365 11112 10429 11116
rect 10445 11172 10509 11176
rect 10445 11116 10449 11172
rect 10449 11116 10505 11172
rect 10505 11116 10509 11172
rect 10445 11112 10509 11116
rect 10525 11172 10589 11176
rect 10525 11116 10529 11172
rect 10529 11116 10585 11172
rect 10585 11116 10589 11172
rect 10525 11112 10589 11116
rect 19618 11172 19682 11176
rect 19618 11116 19622 11172
rect 19622 11116 19678 11172
rect 19678 11116 19682 11172
rect 19618 11112 19682 11116
rect 19698 11172 19762 11176
rect 19698 11116 19702 11172
rect 19702 11116 19758 11172
rect 19758 11116 19762 11172
rect 19698 11112 19762 11116
rect 19778 11172 19842 11176
rect 19778 11116 19782 11172
rect 19782 11116 19838 11172
rect 19838 11116 19842 11172
rect 19778 11112 19842 11116
rect 19858 11172 19922 11176
rect 19858 11116 19862 11172
rect 19862 11116 19918 11172
rect 19918 11116 19922 11172
rect 19858 11112 19922 11116
rect 5618 10628 5682 10632
rect 5618 10572 5622 10628
rect 5622 10572 5678 10628
rect 5678 10572 5682 10628
rect 5618 10568 5682 10572
rect 5698 10628 5762 10632
rect 5698 10572 5702 10628
rect 5702 10572 5758 10628
rect 5758 10572 5762 10628
rect 5698 10568 5762 10572
rect 5778 10628 5842 10632
rect 5778 10572 5782 10628
rect 5782 10572 5838 10628
rect 5838 10572 5842 10628
rect 5778 10568 5842 10572
rect 5858 10628 5922 10632
rect 5858 10572 5862 10628
rect 5862 10572 5918 10628
rect 5918 10572 5922 10628
rect 5858 10568 5922 10572
rect 14952 10628 15016 10632
rect 14952 10572 14956 10628
rect 14956 10572 15012 10628
rect 15012 10572 15016 10628
rect 14952 10568 15016 10572
rect 15032 10628 15096 10632
rect 15032 10572 15036 10628
rect 15036 10572 15092 10628
rect 15092 10572 15096 10628
rect 15032 10568 15096 10572
rect 15112 10628 15176 10632
rect 15112 10572 15116 10628
rect 15116 10572 15172 10628
rect 15172 10572 15176 10628
rect 15112 10568 15176 10572
rect 15192 10628 15256 10632
rect 15192 10572 15196 10628
rect 15196 10572 15252 10628
rect 15252 10572 15256 10628
rect 15192 10568 15256 10572
rect 24285 10628 24349 10632
rect 24285 10572 24289 10628
rect 24289 10572 24345 10628
rect 24345 10572 24349 10628
rect 24285 10568 24349 10572
rect 24365 10628 24429 10632
rect 24365 10572 24369 10628
rect 24369 10572 24425 10628
rect 24425 10572 24429 10628
rect 24365 10568 24429 10572
rect 24445 10628 24509 10632
rect 24445 10572 24449 10628
rect 24449 10572 24505 10628
rect 24505 10572 24509 10628
rect 24445 10568 24509 10572
rect 24525 10628 24589 10632
rect 24525 10572 24529 10628
rect 24529 10572 24585 10628
rect 24585 10572 24589 10628
rect 24525 10568 24589 10572
rect 10285 10084 10349 10088
rect 10285 10028 10289 10084
rect 10289 10028 10345 10084
rect 10345 10028 10349 10084
rect 10285 10024 10349 10028
rect 10365 10084 10429 10088
rect 10365 10028 10369 10084
rect 10369 10028 10425 10084
rect 10425 10028 10429 10084
rect 10365 10024 10429 10028
rect 10445 10084 10509 10088
rect 10445 10028 10449 10084
rect 10449 10028 10505 10084
rect 10505 10028 10509 10084
rect 10445 10024 10509 10028
rect 10525 10084 10589 10088
rect 10525 10028 10529 10084
rect 10529 10028 10585 10084
rect 10585 10028 10589 10084
rect 10525 10024 10589 10028
rect 19618 10084 19682 10088
rect 19618 10028 19622 10084
rect 19622 10028 19678 10084
rect 19678 10028 19682 10084
rect 19618 10024 19682 10028
rect 19698 10084 19762 10088
rect 19698 10028 19702 10084
rect 19702 10028 19758 10084
rect 19758 10028 19762 10084
rect 19698 10024 19762 10028
rect 19778 10084 19842 10088
rect 19778 10028 19782 10084
rect 19782 10028 19838 10084
rect 19838 10028 19842 10084
rect 19778 10024 19842 10028
rect 19858 10084 19922 10088
rect 19858 10028 19862 10084
rect 19862 10028 19918 10084
rect 19918 10028 19922 10084
rect 19858 10024 19922 10028
rect 5618 9540 5682 9544
rect 5618 9484 5622 9540
rect 5622 9484 5678 9540
rect 5678 9484 5682 9540
rect 5618 9480 5682 9484
rect 5698 9540 5762 9544
rect 5698 9484 5702 9540
rect 5702 9484 5758 9540
rect 5758 9484 5762 9540
rect 5698 9480 5762 9484
rect 5778 9540 5842 9544
rect 5778 9484 5782 9540
rect 5782 9484 5838 9540
rect 5838 9484 5842 9540
rect 5778 9480 5842 9484
rect 5858 9540 5922 9544
rect 5858 9484 5862 9540
rect 5862 9484 5918 9540
rect 5918 9484 5922 9540
rect 5858 9480 5922 9484
rect 14952 9540 15016 9544
rect 14952 9484 14956 9540
rect 14956 9484 15012 9540
rect 15012 9484 15016 9540
rect 14952 9480 15016 9484
rect 15032 9540 15096 9544
rect 15032 9484 15036 9540
rect 15036 9484 15092 9540
rect 15092 9484 15096 9540
rect 15032 9480 15096 9484
rect 15112 9540 15176 9544
rect 15112 9484 15116 9540
rect 15116 9484 15172 9540
rect 15172 9484 15176 9540
rect 15112 9480 15176 9484
rect 15192 9540 15256 9544
rect 15192 9484 15196 9540
rect 15196 9484 15252 9540
rect 15252 9484 15256 9540
rect 15192 9480 15256 9484
rect 24285 9540 24349 9544
rect 24285 9484 24289 9540
rect 24289 9484 24345 9540
rect 24345 9484 24349 9540
rect 24285 9480 24349 9484
rect 24365 9540 24429 9544
rect 24365 9484 24369 9540
rect 24369 9484 24425 9540
rect 24425 9484 24429 9540
rect 24365 9480 24429 9484
rect 24445 9540 24509 9544
rect 24445 9484 24449 9540
rect 24449 9484 24505 9540
rect 24505 9484 24509 9540
rect 24445 9480 24509 9484
rect 24525 9540 24589 9544
rect 24525 9484 24529 9540
rect 24529 9484 24585 9540
rect 24585 9484 24589 9540
rect 24525 9480 24589 9484
rect 10285 8996 10349 9000
rect 10285 8940 10289 8996
rect 10289 8940 10345 8996
rect 10345 8940 10349 8996
rect 10285 8936 10349 8940
rect 10365 8996 10429 9000
rect 10365 8940 10369 8996
rect 10369 8940 10425 8996
rect 10425 8940 10429 8996
rect 10365 8936 10429 8940
rect 10445 8996 10509 9000
rect 10445 8940 10449 8996
rect 10449 8940 10505 8996
rect 10505 8940 10509 8996
rect 10445 8936 10509 8940
rect 10525 8996 10589 9000
rect 10525 8940 10529 8996
rect 10529 8940 10585 8996
rect 10585 8940 10589 8996
rect 10525 8936 10589 8940
rect 19618 8996 19682 9000
rect 19618 8940 19622 8996
rect 19622 8940 19678 8996
rect 19678 8940 19682 8996
rect 19618 8936 19682 8940
rect 19698 8996 19762 9000
rect 19698 8940 19702 8996
rect 19702 8940 19758 8996
rect 19758 8940 19762 8996
rect 19698 8936 19762 8940
rect 19778 8996 19842 9000
rect 19778 8940 19782 8996
rect 19782 8940 19838 8996
rect 19838 8940 19842 8996
rect 19778 8936 19842 8940
rect 19858 8996 19922 9000
rect 19858 8940 19862 8996
rect 19862 8940 19918 8996
rect 19918 8940 19922 8996
rect 19858 8936 19922 8940
rect 5618 8452 5682 8456
rect 5618 8396 5622 8452
rect 5622 8396 5678 8452
rect 5678 8396 5682 8452
rect 5618 8392 5682 8396
rect 5698 8452 5762 8456
rect 5698 8396 5702 8452
rect 5702 8396 5758 8452
rect 5758 8396 5762 8452
rect 5698 8392 5762 8396
rect 5778 8452 5842 8456
rect 5778 8396 5782 8452
rect 5782 8396 5838 8452
rect 5838 8396 5842 8452
rect 5778 8392 5842 8396
rect 5858 8452 5922 8456
rect 5858 8396 5862 8452
rect 5862 8396 5918 8452
rect 5918 8396 5922 8452
rect 5858 8392 5922 8396
rect 14952 8452 15016 8456
rect 14952 8396 14956 8452
rect 14956 8396 15012 8452
rect 15012 8396 15016 8452
rect 14952 8392 15016 8396
rect 15032 8452 15096 8456
rect 15032 8396 15036 8452
rect 15036 8396 15092 8452
rect 15092 8396 15096 8452
rect 15032 8392 15096 8396
rect 15112 8452 15176 8456
rect 15112 8396 15116 8452
rect 15116 8396 15172 8452
rect 15172 8396 15176 8452
rect 15112 8392 15176 8396
rect 15192 8452 15256 8456
rect 15192 8396 15196 8452
rect 15196 8396 15252 8452
rect 15252 8396 15256 8452
rect 15192 8392 15256 8396
rect 24285 8452 24349 8456
rect 24285 8396 24289 8452
rect 24289 8396 24345 8452
rect 24345 8396 24349 8452
rect 24285 8392 24349 8396
rect 24365 8452 24429 8456
rect 24365 8396 24369 8452
rect 24369 8396 24425 8452
rect 24425 8396 24429 8452
rect 24365 8392 24429 8396
rect 24445 8452 24509 8456
rect 24445 8396 24449 8452
rect 24449 8396 24505 8452
rect 24505 8396 24509 8452
rect 24445 8392 24509 8396
rect 24525 8452 24589 8456
rect 24525 8396 24529 8452
rect 24529 8396 24585 8452
rect 24585 8396 24589 8452
rect 24525 8392 24589 8396
rect 10285 7908 10349 7912
rect 10285 7852 10289 7908
rect 10289 7852 10345 7908
rect 10345 7852 10349 7908
rect 10285 7848 10349 7852
rect 10365 7908 10429 7912
rect 10365 7852 10369 7908
rect 10369 7852 10425 7908
rect 10425 7852 10429 7908
rect 10365 7848 10429 7852
rect 10445 7908 10509 7912
rect 10445 7852 10449 7908
rect 10449 7852 10505 7908
rect 10505 7852 10509 7908
rect 10445 7848 10509 7852
rect 10525 7908 10589 7912
rect 10525 7852 10529 7908
rect 10529 7852 10585 7908
rect 10585 7852 10589 7908
rect 10525 7848 10589 7852
rect 19618 7908 19682 7912
rect 19618 7852 19622 7908
rect 19622 7852 19678 7908
rect 19678 7852 19682 7908
rect 19618 7848 19682 7852
rect 19698 7908 19762 7912
rect 19698 7852 19702 7908
rect 19702 7852 19758 7908
rect 19758 7852 19762 7908
rect 19698 7848 19762 7852
rect 19778 7908 19842 7912
rect 19778 7852 19782 7908
rect 19782 7852 19838 7908
rect 19838 7852 19842 7908
rect 19778 7848 19842 7852
rect 19858 7908 19922 7912
rect 19858 7852 19862 7908
rect 19862 7852 19918 7908
rect 19918 7852 19922 7908
rect 19858 7848 19922 7852
rect 5618 7364 5682 7368
rect 5618 7308 5622 7364
rect 5622 7308 5678 7364
rect 5678 7308 5682 7364
rect 5618 7304 5682 7308
rect 5698 7364 5762 7368
rect 5698 7308 5702 7364
rect 5702 7308 5758 7364
rect 5758 7308 5762 7364
rect 5698 7304 5762 7308
rect 5778 7364 5842 7368
rect 5778 7308 5782 7364
rect 5782 7308 5838 7364
rect 5838 7308 5842 7364
rect 5778 7304 5842 7308
rect 5858 7364 5922 7368
rect 5858 7308 5862 7364
rect 5862 7308 5918 7364
rect 5918 7308 5922 7364
rect 5858 7304 5922 7308
rect 14952 7364 15016 7368
rect 14952 7308 14956 7364
rect 14956 7308 15012 7364
rect 15012 7308 15016 7364
rect 14952 7304 15016 7308
rect 15032 7364 15096 7368
rect 15032 7308 15036 7364
rect 15036 7308 15092 7364
rect 15092 7308 15096 7364
rect 15032 7304 15096 7308
rect 15112 7364 15176 7368
rect 15112 7308 15116 7364
rect 15116 7308 15172 7364
rect 15172 7308 15176 7364
rect 15112 7304 15176 7308
rect 15192 7364 15256 7368
rect 15192 7308 15196 7364
rect 15196 7308 15252 7364
rect 15252 7308 15256 7364
rect 15192 7304 15256 7308
rect 24285 7364 24349 7368
rect 24285 7308 24289 7364
rect 24289 7308 24345 7364
rect 24345 7308 24349 7364
rect 24285 7304 24349 7308
rect 24365 7364 24429 7368
rect 24365 7308 24369 7364
rect 24369 7308 24425 7364
rect 24425 7308 24429 7364
rect 24365 7304 24429 7308
rect 24445 7364 24509 7368
rect 24445 7308 24449 7364
rect 24449 7308 24505 7364
rect 24505 7308 24509 7364
rect 24445 7304 24509 7308
rect 24525 7364 24589 7368
rect 24525 7308 24529 7364
rect 24529 7308 24585 7364
rect 24585 7308 24589 7364
rect 24525 7304 24589 7308
rect 10285 6820 10349 6824
rect 10285 6764 10289 6820
rect 10289 6764 10345 6820
rect 10345 6764 10349 6820
rect 10285 6760 10349 6764
rect 10365 6820 10429 6824
rect 10365 6764 10369 6820
rect 10369 6764 10425 6820
rect 10425 6764 10429 6820
rect 10365 6760 10429 6764
rect 10445 6820 10509 6824
rect 10445 6764 10449 6820
rect 10449 6764 10505 6820
rect 10505 6764 10509 6820
rect 10445 6760 10509 6764
rect 10525 6820 10589 6824
rect 10525 6764 10529 6820
rect 10529 6764 10585 6820
rect 10585 6764 10589 6820
rect 10525 6760 10589 6764
rect 19618 6820 19682 6824
rect 19618 6764 19622 6820
rect 19622 6764 19678 6820
rect 19678 6764 19682 6820
rect 19618 6760 19682 6764
rect 19698 6820 19762 6824
rect 19698 6764 19702 6820
rect 19702 6764 19758 6820
rect 19758 6764 19762 6820
rect 19698 6760 19762 6764
rect 19778 6820 19842 6824
rect 19778 6764 19782 6820
rect 19782 6764 19838 6820
rect 19838 6764 19842 6820
rect 19778 6760 19842 6764
rect 19858 6820 19922 6824
rect 19858 6764 19862 6820
rect 19862 6764 19918 6820
rect 19918 6764 19922 6820
rect 19858 6760 19922 6764
rect 5618 6276 5682 6280
rect 5618 6220 5622 6276
rect 5622 6220 5678 6276
rect 5678 6220 5682 6276
rect 5618 6216 5682 6220
rect 5698 6276 5762 6280
rect 5698 6220 5702 6276
rect 5702 6220 5758 6276
rect 5758 6220 5762 6276
rect 5698 6216 5762 6220
rect 5778 6276 5842 6280
rect 5778 6220 5782 6276
rect 5782 6220 5838 6276
rect 5838 6220 5842 6276
rect 5778 6216 5842 6220
rect 5858 6276 5922 6280
rect 5858 6220 5862 6276
rect 5862 6220 5918 6276
rect 5918 6220 5922 6276
rect 5858 6216 5922 6220
rect 14952 6276 15016 6280
rect 14952 6220 14956 6276
rect 14956 6220 15012 6276
rect 15012 6220 15016 6276
rect 14952 6216 15016 6220
rect 15032 6276 15096 6280
rect 15032 6220 15036 6276
rect 15036 6220 15092 6276
rect 15092 6220 15096 6276
rect 15032 6216 15096 6220
rect 15112 6276 15176 6280
rect 15112 6220 15116 6276
rect 15116 6220 15172 6276
rect 15172 6220 15176 6276
rect 15112 6216 15176 6220
rect 15192 6276 15256 6280
rect 15192 6220 15196 6276
rect 15196 6220 15252 6276
rect 15252 6220 15256 6276
rect 15192 6216 15256 6220
rect 24285 6276 24349 6280
rect 24285 6220 24289 6276
rect 24289 6220 24345 6276
rect 24345 6220 24349 6276
rect 24285 6216 24349 6220
rect 24365 6276 24429 6280
rect 24365 6220 24369 6276
rect 24369 6220 24425 6276
rect 24425 6220 24429 6276
rect 24365 6216 24429 6220
rect 24445 6276 24509 6280
rect 24445 6220 24449 6276
rect 24449 6220 24505 6276
rect 24505 6220 24509 6276
rect 24445 6216 24509 6220
rect 24525 6276 24589 6280
rect 24525 6220 24529 6276
rect 24529 6220 24585 6276
rect 24585 6220 24589 6276
rect 24525 6216 24589 6220
rect 10285 5732 10349 5736
rect 10285 5676 10289 5732
rect 10289 5676 10345 5732
rect 10345 5676 10349 5732
rect 10285 5672 10349 5676
rect 10365 5732 10429 5736
rect 10365 5676 10369 5732
rect 10369 5676 10425 5732
rect 10425 5676 10429 5732
rect 10365 5672 10429 5676
rect 10445 5732 10509 5736
rect 10445 5676 10449 5732
rect 10449 5676 10505 5732
rect 10505 5676 10509 5732
rect 10445 5672 10509 5676
rect 10525 5732 10589 5736
rect 10525 5676 10529 5732
rect 10529 5676 10585 5732
rect 10585 5676 10589 5732
rect 10525 5672 10589 5676
rect 19618 5732 19682 5736
rect 19618 5676 19622 5732
rect 19622 5676 19678 5732
rect 19678 5676 19682 5732
rect 19618 5672 19682 5676
rect 19698 5732 19762 5736
rect 19698 5676 19702 5732
rect 19702 5676 19758 5732
rect 19758 5676 19762 5732
rect 19698 5672 19762 5676
rect 19778 5732 19842 5736
rect 19778 5676 19782 5732
rect 19782 5676 19838 5732
rect 19838 5676 19842 5732
rect 19778 5672 19842 5676
rect 19858 5732 19922 5736
rect 19858 5676 19862 5732
rect 19862 5676 19918 5732
rect 19918 5676 19922 5732
rect 19858 5672 19922 5676
rect 5618 5188 5682 5192
rect 5618 5132 5622 5188
rect 5622 5132 5678 5188
rect 5678 5132 5682 5188
rect 5618 5128 5682 5132
rect 5698 5188 5762 5192
rect 5698 5132 5702 5188
rect 5702 5132 5758 5188
rect 5758 5132 5762 5188
rect 5698 5128 5762 5132
rect 5778 5188 5842 5192
rect 5778 5132 5782 5188
rect 5782 5132 5838 5188
rect 5838 5132 5842 5188
rect 5778 5128 5842 5132
rect 5858 5188 5922 5192
rect 5858 5132 5862 5188
rect 5862 5132 5918 5188
rect 5918 5132 5922 5188
rect 5858 5128 5922 5132
rect 14952 5188 15016 5192
rect 14952 5132 14956 5188
rect 14956 5132 15012 5188
rect 15012 5132 15016 5188
rect 14952 5128 15016 5132
rect 15032 5188 15096 5192
rect 15032 5132 15036 5188
rect 15036 5132 15092 5188
rect 15092 5132 15096 5188
rect 15032 5128 15096 5132
rect 15112 5188 15176 5192
rect 15112 5132 15116 5188
rect 15116 5132 15172 5188
rect 15172 5132 15176 5188
rect 15112 5128 15176 5132
rect 15192 5188 15256 5192
rect 15192 5132 15196 5188
rect 15196 5132 15252 5188
rect 15252 5132 15256 5188
rect 15192 5128 15256 5132
rect 24285 5188 24349 5192
rect 24285 5132 24289 5188
rect 24289 5132 24345 5188
rect 24345 5132 24349 5188
rect 24285 5128 24349 5132
rect 24365 5188 24429 5192
rect 24365 5132 24369 5188
rect 24369 5132 24425 5188
rect 24425 5132 24429 5188
rect 24365 5128 24429 5132
rect 24445 5188 24509 5192
rect 24445 5132 24449 5188
rect 24449 5132 24505 5188
rect 24505 5132 24509 5188
rect 24445 5128 24509 5132
rect 24525 5188 24589 5192
rect 24525 5132 24529 5188
rect 24529 5132 24585 5188
rect 24585 5132 24589 5188
rect 24525 5128 24589 5132
rect 10285 4644 10349 4648
rect 10285 4588 10289 4644
rect 10289 4588 10345 4644
rect 10345 4588 10349 4644
rect 10285 4584 10349 4588
rect 10365 4644 10429 4648
rect 10365 4588 10369 4644
rect 10369 4588 10425 4644
rect 10425 4588 10429 4644
rect 10365 4584 10429 4588
rect 10445 4644 10509 4648
rect 10445 4588 10449 4644
rect 10449 4588 10505 4644
rect 10505 4588 10509 4644
rect 10445 4584 10509 4588
rect 10525 4644 10589 4648
rect 10525 4588 10529 4644
rect 10529 4588 10585 4644
rect 10585 4588 10589 4644
rect 10525 4584 10589 4588
rect 19618 4644 19682 4648
rect 19618 4588 19622 4644
rect 19622 4588 19678 4644
rect 19678 4588 19682 4644
rect 19618 4584 19682 4588
rect 19698 4644 19762 4648
rect 19698 4588 19702 4644
rect 19702 4588 19758 4644
rect 19758 4588 19762 4644
rect 19698 4584 19762 4588
rect 19778 4644 19842 4648
rect 19778 4588 19782 4644
rect 19782 4588 19838 4644
rect 19838 4588 19842 4644
rect 19778 4584 19842 4588
rect 19858 4644 19922 4648
rect 19858 4588 19862 4644
rect 19862 4588 19918 4644
rect 19918 4588 19922 4644
rect 19858 4584 19922 4588
rect 5618 4100 5682 4104
rect 5618 4044 5622 4100
rect 5622 4044 5678 4100
rect 5678 4044 5682 4100
rect 5618 4040 5682 4044
rect 5698 4100 5762 4104
rect 5698 4044 5702 4100
rect 5702 4044 5758 4100
rect 5758 4044 5762 4100
rect 5698 4040 5762 4044
rect 5778 4100 5842 4104
rect 5778 4044 5782 4100
rect 5782 4044 5838 4100
rect 5838 4044 5842 4100
rect 5778 4040 5842 4044
rect 5858 4100 5922 4104
rect 5858 4044 5862 4100
rect 5862 4044 5918 4100
rect 5918 4044 5922 4100
rect 5858 4040 5922 4044
rect 14952 4100 15016 4104
rect 14952 4044 14956 4100
rect 14956 4044 15012 4100
rect 15012 4044 15016 4100
rect 14952 4040 15016 4044
rect 15032 4100 15096 4104
rect 15032 4044 15036 4100
rect 15036 4044 15092 4100
rect 15092 4044 15096 4100
rect 15032 4040 15096 4044
rect 15112 4100 15176 4104
rect 15112 4044 15116 4100
rect 15116 4044 15172 4100
rect 15172 4044 15176 4100
rect 15112 4040 15176 4044
rect 15192 4100 15256 4104
rect 15192 4044 15196 4100
rect 15196 4044 15252 4100
rect 15252 4044 15256 4100
rect 15192 4040 15256 4044
rect 24285 4100 24349 4104
rect 24285 4044 24289 4100
rect 24289 4044 24345 4100
rect 24345 4044 24349 4100
rect 24285 4040 24349 4044
rect 24365 4100 24429 4104
rect 24365 4044 24369 4100
rect 24369 4044 24425 4100
rect 24425 4044 24429 4100
rect 24365 4040 24429 4044
rect 24445 4100 24509 4104
rect 24445 4044 24449 4100
rect 24449 4044 24505 4100
rect 24505 4044 24509 4100
rect 24445 4040 24509 4044
rect 24525 4100 24589 4104
rect 24525 4044 24529 4100
rect 24529 4044 24585 4100
rect 24585 4044 24589 4100
rect 24525 4040 24589 4044
rect 10285 3556 10349 3560
rect 10285 3500 10289 3556
rect 10289 3500 10345 3556
rect 10345 3500 10349 3556
rect 10285 3496 10349 3500
rect 10365 3556 10429 3560
rect 10365 3500 10369 3556
rect 10369 3500 10425 3556
rect 10425 3500 10429 3556
rect 10365 3496 10429 3500
rect 10445 3556 10509 3560
rect 10445 3500 10449 3556
rect 10449 3500 10505 3556
rect 10505 3500 10509 3556
rect 10445 3496 10509 3500
rect 10525 3556 10589 3560
rect 10525 3500 10529 3556
rect 10529 3500 10585 3556
rect 10585 3500 10589 3556
rect 10525 3496 10589 3500
rect 19618 3556 19682 3560
rect 19618 3500 19622 3556
rect 19622 3500 19678 3556
rect 19678 3500 19682 3556
rect 19618 3496 19682 3500
rect 19698 3556 19762 3560
rect 19698 3500 19702 3556
rect 19702 3500 19758 3556
rect 19758 3500 19762 3556
rect 19698 3496 19762 3500
rect 19778 3556 19842 3560
rect 19778 3500 19782 3556
rect 19782 3500 19838 3556
rect 19838 3500 19842 3556
rect 19778 3496 19842 3500
rect 19858 3556 19922 3560
rect 19858 3500 19862 3556
rect 19862 3500 19918 3556
rect 19918 3500 19922 3556
rect 19858 3496 19922 3500
rect 5618 3012 5682 3016
rect 5618 2956 5622 3012
rect 5622 2956 5678 3012
rect 5678 2956 5682 3012
rect 5618 2952 5682 2956
rect 5698 3012 5762 3016
rect 5698 2956 5702 3012
rect 5702 2956 5758 3012
rect 5758 2956 5762 3012
rect 5698 2952 5762 2956
rect 5778 3012 5842 3016
rect 5778 2956 5782 3012
rect 5782 2956 5838 3012
rect 5838 2956 5842 3012
rect 5778 2952 5842 2956
rect 5858 3012 5922 3016
rect 5858 2956 5862 3012
rect 5862 2956 5918 3012
rect 5918 2956 5922 3012
rect 5858 2952 5922 2956
rect 14952 3012 15016 3016
rect 14952 2956 14956 3012
rect 14956 2956 15012 3012
rect 15012 2956 15016 3012
rect 14952 2952 15016 2956
rect 15032 3012 15096 3016
rect 15032 2956 15036 3012
rect 15036 2956 15092 3012
rect 15092 2956 15096 3012
rect 15032 2952 15096 2956
rect 15112 3012 15176 3016
rect 15112 2956 15116 3012
rect 15116 2956 15172 3012
rect 15172 2956 15176 3012
rect 15112 2952 15176 2956
rect 15192 3012 15256 3016
rect 15192 2956 15196 3012
rect 15196 2956 15252 3012
rect 15252 2956 15256 3012
rect 15192 2952 15256 2956
rect 24285 3012 24349 3016
rect 24285 2956 24289 3012
rect 24289 2956 24345 3012
rect 24345 2956 24349 3012
rect 24285 2952 24349 2956
rect 24365 3012 24429 3016
rect 24365 2956 24369 3012
rect 24369 2956 24425 3012
rect 24425 2956 24429 3012
rect 24365 2952 24429 2956
rect 24445 3012 24509 3016
rect 24445 2956 24449 3012
rect 24449 2956 24505 3012
rect 24505 2956 24509 3012
rect 24445 2952 24509 2956
rect 24525 3012 24589 3016
rect 24525 2956 24529 3012
rect 24529 2956 24585 3012
rect 24585 2956 24589 3012
rect 24525 2952 24589 2956
rect 10285 2468 10349 2472
rect 10285 2412 10289 2468
rect 10289 2412 10345 2468
rect 10345 2412 10349 2468
rect 10285 2408 10349 2412
rect 10365 2468 10429 2472
rect 10365 2412 10369 2468
rect 10369 2412 10425 2468
rect 10425 2412 10429 2468
rect 10365 2408 10429 2412
rect 10445 2468 10509 2472
rect 10445 2412 10449 2468
rect 10449 2412 10505 2468
rect 10505 2412 10509 2468
rect 10445 2408 10509 2412
rect 10525 2468 10589 2472
rect 10525 2412 10529 2468
rect 10529 2412 10585 2468
rect 10585 2412 10589 2468
rect 10525 2408 10589 2412
rect 19618 2468 19682 2472
rect 19618 2412 19622 2468
rect 19622 2412 19678 2468
rect 19678 2412 19682 2468
rect 19618 2408 19682 2412
rect 19698 2468 19762 2472
rect 19698 2412 19702 2468
rect 19702 2412 19758 2468
rect 19758 2412 19762 2468
rect 19698 2408 19762 2412
rect 19778 2468 19842 2472
rect 19778 2412 19782 2468
rect 19782 2412 19838 2468
rect 19838 2412 19842 2468
rect 19778 2408 19842 2412
rect 19858 2468 19922 2472
rect 19858 2412 19862 2468
rect 19862 2412 19918 2468
rect 19918 2412 19922 2468
rect 19858 2408 19922 2412
rect 5618 1924 5682 1928
rect 5618 1868 5622 1924
rect 5622 1868 5678 1924
rect 5678 1868 5682 1924
rect 5618 1864 5682 1868
rect 5698 1924 5762 1928
rect 5698 1868 5702 1924
rect 5702 1868 5758 1924
rect 5758 1868 5762 1924
rect 5698 1864 5762 1868
rect 5778 1924 5842 1928
rect 5778 1868 5782 1924
rect 5782 1868 5838 1924
rect 5838 1868 5842 1924
rect 5778 1864 5842 1868
rect 5858 1924 5922 1928
rect 5858 1868 5862 1924
rect 5862 1868 5918 1924
rect 5918 1868 5922 1924
rect 5858 1864 5922 1868
rect 14952 1924 15016 1928
rect 14952 1868 14956 1924
rect 14956 1868 15012 1924
rect 15012 1868 15016 1924
rect 14952 1864 15016 1868
rect 15032 1924 15096 1928
rect 15032 1868 15036 1924
rect 15036 1868 15092 1924
rect 15092 1868 15096 1924
rect 15032 1864 15096 1868
rect 15112 1924 15176 1928
rect 15112 1868 15116 1924
rect 15116 1868 15172 1924
rect 15172 1868 15176 1924
rect 15112 1864 15176 1868
rect 15192 1924 15256 1928
rect 15192 1868 15196 1924
rect 15196 1868 15252 1924
rect 15252 1868 15256 1924
rect 15192 1864 15256 1868
rect 24285 1924 24349 1928
rect 24285 1868 24289 1924
rect 24289 1868 24345 1924
rect 24345 1868 24349 1924
rect 24285 1864 24349 1868
rect 24365 1924 24429 1928
rect 24365 1868 24369 1924
rect 24369 1868 24425 1924
rect 24425 1868 24429 1924
rect 24365 1864 24429 1868
rect 24445 1924 24509 1928
rect 24445 1868 24449 1924
rect 24449 1868 24505 1924
rect 24505 1868 24509 1924
rect 24445 1864 24509 1868
rect 24525 1924 24589 1928
rect 24525 1868 24529 1924
rect 24529 1868 24585 1924
rect 24585 1868 24589 1924
rect 24525 1864 24589 1868
<< metal4 >>
rect 5610 24776 5931 25336
rect 5610 24712 5618 24776
rect 5682 24712 5698 24776
rect 5762 24712 5778 24776
rect 5842 24712 5858 24776
rect 5922 24712 5931 24776
rect 5610 23688 5931 24712
rect 10277 25320 10597 25336
rect 10277 25256 10285 25320
rect 10349 25256 10365 25320
rect 10429 25256 10445 25320
rect 10509 25256 10525 25320
rect 10589 25256 10597 25320
rect 10277 24232 10597 25256
rect 10277 24168 10285 24232
rect 10349 24168 10365 24232
rect 10429 24168 10445 24232
rect 10509 24168 10525 24232
rect 10589 24168 10597 24232
rect 6131 23892 6197 23893
rect 6131 23828 6132 23892
rect 6196 23828 6197 23892
rect 6131 23827 6197 23828
rect 5610 23624 5618 23688
rect 5682 23624 5698 23688
rect 5762 23624 5778 23688
rect 5842 23624 5858 23688
rect 5922 23624 5931 23688
rect 5610 22600 5931 23624
rect 5610 22536 5618 22600
rect 5682 22536 5698 22600
rect 5762 22536 5778 22600
rect 5842 22536 5858 22600
rect 5922 22536 5931 22600
rect 5610 21512 5931 22536
rect 5610 21448 5618 21512
rect 5682 21448 5698 21512
rect 5762 21448 5778 21512
rect 5842 21448 5858 21512
rect 5922 21448 5931 21512
rect 5610 20424 5931 21448
rect 6134 21258 6194 23827
rect 10277 23144 10597 24168
rect 14944 24776 15264 25336
rect 14944 24712 14952 24776
rect 15016 24712 15032 24776
rect 15096 24712 15112 24776
rect 15176 24712 15192 24776
rect 15256 24712 15264 24776
rect 14944 23688 15264 24712
rect 14944 23624 14952 23688
rect 15016 23624 15032 23688
rect 15096 23624 15112 23688
rect 15176 23624 15192 23688
rect 15256 23624 15264 23688
rect 10915 23212 10981 23213
rect 10915 23148 10916 23212
rect 10980 23148 10981 23212
rect 10915 23147 10981 23148
rect 10277 23080 10285 23144
rect 10349 23080 10365 23144
rect 10429 23080 10445 23144
rect 10509 23080 10525 23144
rect 10589 23080 10597 23144
rect 10277 22056 10597 23080
rect 10277 21992 10285 22056
rect 10349 21992 10365 22056
rect 10429 21992 10445 22056
rect 10509 21992 10525 22056
rect 10589 21992 10597 22056
rect 5610 20360 5618 20424
rect 5682 20360 5698 20424
rect 5762 20360 5778 20424
rect 5842 20360 5858 20424
rect 5922 20360 5931 20424
rect 5610 19336 5931 20360
rect 5610 19272 5618 19336
rect 5682 19272 5698 19336
rect 5762 19272 5778 19336
rect 5842 19272 5858 19336
rect 5922 19272 5931 19336
rect 5610 18248 5931 19272
rect 5610 18184 5618 18248
rect 5682 18184 5698 18248
rect 5762 18184 5778 18248
rect 5842 18184 5858 18248
rect 5922 18184 5931 18248
rect 5610 17160 5931 18184
rect 5610 17096 5618 17160
rect 5682 17096 5698 17160
rect 5762 17096 5778 17160
rect 5842 17096 5858 17160
rect 5922 17096 5931 17160
rect 5610 16072 5931 17096
rect 5610 16008 5618 16072
rect 5682 16008 5698 16072
rect 5762 16008 5778 16072
rect 5842 16008 5858 16072
rect 5922 16008 5931 16072
rect 5610 14984 5931 16008
rect 5610 14920 5618 14984
rect 5682 14920 5698 14984
rect 5762 14920 5778 14984
rect 5842 14920 5858 14984
rect 5922 14920 5931 14984
rect 5610 13896 5931 14920
rect 5610 13832 5618 13896
rect 5682 13832 5698 13896
rect 5762 13832 5778 13896
rect 5842 13832 5858 13896
rect 5922 13832 5931 13896
rect 5610 12808 5931 13832
rect 5610 12744 5618 12808
rect 5682 12744 5698 12808
rect 5762 12744 5778 12808
rect 5842 12744 5858 12808
rect 5922 12744 5931 12808
rect 5610 11720 5931 12744
rect 5610 11656 5618 11720
rect 5682 11656 5698 11720
rect 5762 11656 5778 11720
rect 5842 11656 5858 11720
rect 5922 11656 5931 11720
rect 5610 10632 5931 11656
rect 5610 10568 5618 10632
rect 5682 10568 5698 10632
rect 5762 10568 5778 10632
rect 5842 10568 5858 10632
rect 5922 10568 5931 10632
rect 5610 9544 5931 10568
rect 5610 9480 5618 9544
rect 5682 9480 5698 9544
rect 5762 9480 5778 9544
rect 5842 9480 5858 9544
rect 5922 9480 5931 9544
rect 5610 8456 5931 9480
rect 5610 8392 5618 8456
rect 5682 8392 5698 8456
rect 5762 8392 5778 8456
rect 5842 8392 5858 8456
rect 5922 8392 5931 8456
rect 5610 7368 5931 8392
rect 5610 7304 5618 7368
rect 5682 7304 5698 7368
rect 5762 7304 5778 7368
rect 5842 7304 5858 7368
rect 5922 7304 5931 7368
rect 5610 6280 5931 7304
rect 5610 6216 5618 6280
rect 5682 6216 5698 6280
rect 5762 6216 5778 6280
rect 5842 6216 5858 6280
rect 5922 6216 5931 6280
rect 5610 5192 5931 6216
rect 5610 5128 5618 5192
rect 5682 5128 5698 5192
rect 5762 5128 5778 5192
rect 5842 5128 5858 5192
rect 5922 5128 5931 5192
rect 5610 4104 5931 5128
rect 5610 4040 5618 4104
rect 5682 4040 5698 4104
rect 5762 4040 5778 4104
rect 5842 4040 5858 4104
rect 5922 4040 5931 4104
rect 5610 3016 5931 4040
rect 5610 2952 5618 3016
rect 5682 2952 5698 3016
rect 5762 2952 5778 3016
rect 5842 2952 5858 3016
rect 5922 2952 5931 3016
rect 5610 1928 5931 2952
rect 5610 1864 5618 1928
rect 5682 1864 5698 1928
rect 5762 1864 5778 1928
rect 5842 1864 5858 1928
rect 5922 1864 5931 1928
rect 5610 1848 5931 1864
rect 10277 20968 10597 21992
rect 10277 20904 10285 20968
rect 10349 20904 10365 20968
rect 10429 20904 10445 20968
rect 10509 20904 10525 20968
rect 10589 20904 10597 20968
rect 10277 19880 10597 20904
rect 10918 20578 10978 23147
rect 14944 22600 15264 23624
rect 14944 22536 14952 22600
rect 15016 22536 15032 22600
rect 15096 22536 15112 22600
rect 15176 22536 15192 22600
rect 15256 22536 15264 22600
rect 14944 21512 15264 22536
rect 14944 21448 14952 21512
rect 15016 21448 15032 21512
rect 15096 21448 15112 21512
rect 15176 21448 15192 21512
rect 15256 21448 15264 21512
rect 14944 20424 15264 21448
rect 14944 20360 14952 20424
rect 15016 20360 15032 20424
rect 15096 20360 15112 20424
rect 15176 20360 15192 20424
rect 15256 20360 15264 20424
rect 10277 19816 10285 19880
rect 10349 19816 10365 19880
rect 10429 19816 10445 19880
rect 10509 19816 10525 19880
rect 10589 19816 10597 19880
rect 10277 18792 10597 19816
rect 10277 18728 10285 18792
rect 10349 18728 10365 18792
rect 10429 18728 10445 18792
rect 10509 18728 10525 18792
rect 10589 18728 10597 18792
rect 10277 17704 10597 18728
rect 10277 17640 10285 17704
rect 10349 17640 10365 17704
rect 10429 17640 10445 17704
rect 10509 17640 10525 17704
rect 10589 17640 10597 17704
rect 10277 16616 10597 17640
rect 10277 16552 10285 16616
rect 10349 16552 10365 16616
rect 10429 16552 10445 16616
rect 10509 16552 10525 16616
rect 10589 16552 10597 16616
rect 10277 15528 10597 16552
rect 10277 15464 10285 15528
rect 10349 15464 10365 15528
rect 10429 15464 10445 15528
rect 10509 15464 10525 15528
rect 10589 15464 10597 15528
rect 10277 14440 10597 15464
rect 10277 14376 10285 14440
rect 10349 14376 10365 14440
rect 10429 14376 10445 14440
rect 10509 14376 10525 14440
rect 10589 14376 10597 14440
rect 10277 13352 10597 14376
rect 10277 13288 10285 13352
rect 10349 13288 10365 13352
rect 10429 13288 10445 13352
rect 10509 13288 10525 13352
rect 10589 13288 10597 13352
rect 10277 12264 10597 13288
rect 10277 12200 10285 12264
rect 10349 12200 10365 12264
rect 10429 12200 10445 12264
rect 10509 12200 10525 12264
rect 10589 12200 10597 12264
rect 10277 11176 10597 12200
rect 10277 11112 10285 11176
rect 10349 11112 10365 11176
rect 10429 11112 10445 11176
rect 10509 11112 10525 11176
rect 10589 11112 10597 11176
rect 10277 10088 10597 11112
rect 10277 10024 10285 10088
rect 10349 10024 10365 10088
rect 10429 10024 10445 10088
rect 10509 10024 10525 10088
rect 10589 10024 10597 10088
rect 10277 9000 10597 10024
rect 10277 8936 10285 9000
rect 10349 8936 10365 9000
rect 10429 8936 10445 9000
rect 10509 8936 10525 9000
rect 10589 8936 10597 9000
rect 10277 7912 10597 8936
rect 10277 7848 10285 7912
rect 10349 7848 10365 7912
rect 10429 7848 10445 7912
rect 10509 7848 10525 7912
rect 10589 7848 10597 7912
rect 10277 6824 10597 7848
rect 10277 6760 10285 6824
rect 10349 6760 10365 6824
rect 10429 6760 10445 6824
rect 10509 6760 10525 6824
rect 10589 6760 10597 6824
rect 10277 5736 10597 6760
rect 10277 5672 10285 5736
rect 10349 5672 10365 5736
rect 10429 5672 10445 5736
rect 10509 5672 10525 5736
rect 10589 5672 10597 5736
rect 10277 4648 10597 5672
rect 10277 4584 10285 4648
rect 10349 4584 10365 4648
rect 10429 4584 10445 4648
rect 10509 4584 10525 4648
rect 10589 4584 10597 4648
rect 10277 3560 10597 4584
rect 10277 3496 10285 3560
rect 10349 3496 10365 3560
rect 10429 3496 10445 3560
rect 10509 3496 10525 3560
rect 10589 3496 10597 3560
rect 10277 2472 10597 3496
rect 10277 2408 10285 2472
rect 10349 2408 10365 2472
rect 10429 2408 10445 2472
rect 10509 2408 10525 2472
rect 10589 2408 10597 2472
rect 10277 1848 10597 2408
rect 14944 19336 15264 20360
rect 14944 19272 14952 19336
rect 15016 19272 15032 19336
rect 15096 19272 15112 19336
rect 15176 19272 15192 19336
rect 15256 19272 15264 19336
rect 14944 18248 15264 19272
rect 14944 18184 14952 18248
rect 15016 18184 15032 18248
rect 15096 18184 15112 18248
rect 15176 18184 15192 18248
rect 15256 18184 15264 18248
rect 14944 17160 15264 18184
rect 14944 17096 14952 17160
rect 15016 17096 15032 17160
rect 15096 17096 15112 17160
rect 15176 17096 15192 17160
rect 15256 17096 15264 17160
rect 14944 16072 15264 17096
rect 14944 16008 14952 16072
rect 15016 16008 15032 16072
rect 15096 16008 15112 16072
rect 15176 16008 15192 16072
rect 15256 16008 15264 16072
rect 14944 14984 15264 16008
rect 14944 14920 14952 14984
rect 15016 14920 15032 14984
rect 15096 14920 15112 14984
rect 15176 14920 15192 14984
rect 15256 14920 15264 14984
rect 14944 13896 15264 14920
rect 14944 13832 14952 13896
rect 15016 13832 15032 13896
rect 15096 13832 15112 13896
rect 15176 13832 15192 13896
rect 15256 13832 15264 13896
rect 14944 12808 15264 13832
rect 14944 12744 14952 12808
rect 15016 12744 15032 12808
rect 15096 12744 15112 12808
rect 15176 12744 15192 12808
rect 15256 12744 15264 12808
rect 14944 11720 15264 12744
rect 14944 11656 14952 11720
rect 15016 11656 15032 11720
rect 15096 11656 15112 11720
rect 15176 11656 15192 11720
rect 15256 11656 15264 11720
rect 14944 10632 15264 11656
rect 14944 10568 14952 10632
rect 15016 10568 15032 10632
rect 15096 10568 15112 10632
rect 15176 10568 15192 10632
rect 15256 10568 15264 10632
rect 14944 9544 15264 10568
rect 14944 9480 14952 9544
rect 15016 9480 15032 9544
rect 15096 9480 15112 9544
rect 15176 9480 15192 9544
rect 15256 9480 15264 9544
rect 14944 8456 15264 9480
rect 14944 8392 14952 8456
rect 15016 8392 15032 8456
rect 15096 8392 15112 8456
rect 15176 8392 15192 8456
rect 15256 8392 15264 8456
rect 14944 7368 15264 8392
rect 14944 7304 14952 7368
rect 15016 7304 15032 7368
rect 15096 7304 15112 7368
rect 15176 7304 15192 7368
rect 15256 7304 15264 7368
rect 14944 6280 15264 7304
rect 14944 6216 14952 6280
rect 15016 6216 15032 6280
rect 15096 6216 15112 6280
rect 15176 6216 15192 6280
rect 15256 6216 15264 6280
rect 14944 5192 15264 6216
rect 14944 5128 14952 5192
rect 15016 5128 15032 5192
rect 15096 5128 15112 5192
rect 15176 5128 15192 5192
rect 15256 5128 15264 5192
rect 14944 4104 15264 5128
rect 14944 4040 14952 4104
rect 15016 4040 15032 4104
rect 15096 4040 15112 4104
rect 15176 4040 15192 4104
rect 15256 4040 15264 4104
rect 14944 3016 15264 4040
rect 14944 2952 14952 3016
rect 15016 2952 15032 3016
rect 15096 2952 15112 3016
rect 15176 2952 15192 3016
rect 15256 2952 15264 3016
rect 14944 1928 15264 2952
rect 14944 1864 14952 1928
rect 15016 1864 15032 1928
rect 15096 1864 15112 1928
rect 15176 1864 15192 1928
rect 15256 1864 15264 1928
rect 14944 1848 15264 1864
rect 19610 25320 19930 25336
rect 19610 25256 19618 25320
rect 19682 25256 19698 25320
rect 19762 25256 19778 25320
rect 19842 25256 19858 25320
rect 19922 25256 19930 25320
rect 19610 24232 19930 25256
rect 19610 24168 19618 24232
rect 19682 24168 19698 24232
rect 19762 24168 19778 24232
rect 19842 24168 19858 24232
rect 19922 24168 19930 24232
rect 19610 23144 19930 24168
rect 19610 23080 19618 23144
rect 19682 23080 19698 23144
rect 19762 23080 19778 23144
rect 19842 23080 19858 23144
rect 19922 23080 19930 23144
rect 19610 22056 19930 23080
rect 19610 21992 19618 22056
rect 19682 21992 19698 22056
rect 19762 21992 19778 22056
rect 19842 21992 19858 22056
rect 19922 21992 19930 22056
rect 19610 20968 19930 21992
rect 24277 24776 24597 25336
rect 24277 24712 24285 24776
rect 24349 24712 24365 24776
rect 24429 24712 24445 24776
rect 24509 24712 24525 24776
rect 24589 24712 24597 24776
rect 24277 23688 24597 24712
rect 24277 23624 24285 23688
rect 24349 23624 24365 23688
rect 24429 23624 24445 23688
rect 24509 23624 24525 23688
rect 24589 23624 24597 23688
rect 24277 22600 24597 23624
rect 24277 22536 24285 22600
rect 24349 22536 24365 22600
rect 24429 22536 24445 22600
rect 24509 22536 24525 22600
rect 24589 22536 24597 22600
rect 24277 21512 24597 22536
rect 24277 21448 24285 21512
rect 24349 21448 24365 21512
rect 24429 21448 24445 21512
rect 24509 21448 24525 21512
rect 24589 21448 24597 21512
rect 19610 20904 19618 20968
rect 19682 20904 19698 20968
rect 19762 20904 19778 20968
rect 19842 20904 19858 20968
rect 19922 20904 19930 20968
rect 19610 19880 19930 20904
rect 21222 20901 21282 21022
rect 21219 20900 21285 20901
rect 21219 20836 21220 20900
rect 21284 20836 21285 20900
rect 21219 20835 21285 20836
rect 23979 20628 24045 20629
rect 23979 20578 23980 20628
rect 24044 20578 24045 20628
rect 24277 20424 24597 21448
rect 24277 20360 24285 20424
rect 24349 20360 24365 20424
rect 24429 20360 24445 20424
rect 24509 20360 24525 20424
rect 24589 20360 24597 20424
rect 19610 19816 19618 19880
rect 19682 19816 19698 19880
rect 19762 19816 19778 19880
rect 19842 19816 19858 19880
rect 19922 19816 19930 19880
rect 19610 18792 19930 19816
rect 19610 18728 19618 18792
rect 19682 18728 19698 18792
rect 19762 18728 19778 18792
rect 19842 18728 19858 18792
rect 19922 18728 19930 18792
rect 19610 17704 19930 18728
rect 19610 17640 19618 17704
rect 19682 17640 19698 17704
rect 19762 17640 19778 17704
rect 19842 17640 19858 17704
rect 19922 17640 19930 17704
rect 19610 16616 19930 17640
rect 19610 16552 19618 16616
rect 19682 16552 19698 16616
rect 19762 16552 19778 16616
rect 19842 16552 19858 16616
rect 19922 16552 19930 16616
rect 19610 15528 19930 16552
rect 19610 15464 19618 15528
rect 19682 15464 19698 15528
rect 19762 15464 19778 15528
rect 19842 15464 19858 15528
rect 19922 15464 19930 15528
rect 19610 14440 19930 15464
rect 19610 14376 19618 14440
rect 19682 14376 19698 14440
rect 19762 14376 19778 14440
rect 19842 14376 19858 14440
rect 19922 14376 19930 14440
rect 19610 13352 19930 14376
rect 19610 13288 19618 13352
rect 19682 13288 19698 13352
rect 19762 13288 19778 13352
rect 19842 13288 19858 13352
rect 19922 13288 19930 13352
rect 19610 12264 19930 13288
rect 19610 12200 19618 12264
rect 19682 12200 19698 12264
rect 19762 12200 19778 12264
rect 19842 12200 19858 12264
rect 19922 12200 19930 12264
rect 19610 11176 19930 12200
rect 19610 11112 19618 11176
rect 19682 11112 19698 11176
rect 19762 11112 19778 11176
rect 19842 11112 19858 11176
rect 19922 11112 19930 11176
rect 19610 10088 19930 11112
rect 19610 10024 19618 10088
rect 19682 10024 19698 10088
rect 19762 10024 19778 10088
rect 19842 10024 19858 10088
rect 19922 10024 19930 10088
rect 19610 9000 19930 10024
rect 19610 8936 19618 9000
rect 19682 8936 19698 9000
rect 19762 8936 19778 9000
rect 19842 8936 19858 9000
rect 19922 8936 19930 9000
rect 19610 7912 19930 8936
rect 19610 7848 19618 7912
rect 19682 7848 19698 7912
rect 19762 7848 19778 7912
rect 19842 7848 19858 7912
rect 19922 7848 19930 7912
rect 19610 6824 19930 7848
rect 19610 6760 19618 6824
rect 19682 6760 19698 6824
rect 19762 6760 19778 6824
rect 19842 6760 19858 6824
rect 19922 6760 19930 6824
rect 19610 5736 19930 6760
rect 19610 5672 19618 5736
rect 19682 5672 19698 5736
rect 19762 5672 19778 5736
rect 19842 5672 19858 5736
rect 19922 5672 19930 5736
rect 19610 4648 19930 5672
rect 19610 4584 19618 4648
rect 19682 4584 19698 4648
rect 19762 4584 19778 4648
rect 19842 4584 19858 4648
rect 19922 4584 19930 4648
rect 19610 3560 19930 4584
rect 19610 3496 19618 3560
rect 19682 3496 19698 3560
rect 19762 3496 19778 3560
rect 19842 3496 19858 3560
rect 19922 3496 19930 3560
rect 19610 2472 19930 3496
rect 19610 2408 19618 2472
rect 19682 2408 19698 2472
rect 19762 2408 19778 2472
rect 19842 2408 19858 2472
rect 19922 2408 19930 2472
rect 19610 1848 19930 2408
rect 24277 19336 24597 20360
rect 24277 19272 24285 19336
rect 24349 19272 24365 19336
rect 24429 19272 24445 19336
rect 24509 19272 24525 19336
rect 24589 19272 24597 19336
rect 24277 18248 24597 19272
rect 24277 18184 24285 18248
rect 24349 18184 24365 18248
rect 24429 18184 24445 18248
rect 24509 18184 24525 18248
rect 24589 18184 24597 18248
rect 24277 17160 24597 18184
rect 24277 17096 24285 17160
rect 24349 17096 24365 17160
rect 24429 17096 24445 17160
rect 24509 17096 24525 17160
rect 24589 17096 24597 17160
rect 24277 16072 24597 17096
rect 24277 16008 24285 16072
rect 24349 16008 24365 16072
rect 24429 16008 24445 16072
rect 24509 16008 24525 16072
rect 24589 16008 24597 16072
rect 24277 14984 24597 16008
rect 24277 14920 24285 14984
rect 24349 14920 24365 14984
rect 24429 14920 24445 14984
rect 24509 14920 24525 14984
rect 24589 14920 24597 14984
rect 24277 13896 24597 14920
rect 24277 13832 24285 13896
rect 24349 13832 24365 13896
rect 24429 13832 24445 13896
rect 24509 13832 24525 13896
rect 24589 13832 24597 13896
rect 24277 12808 24597 13832
rect 24277 12744 24285 12808
rect 24349 12744 24365 12808
rect 24429 12744 24445 12808
rect 24509 12744 24525 12808
rect 24589 12744 24597 12808
rect 24277 11720 24597 12744
rect 24277 11656 24285 11720
rect 24349 11656 24365 11720
rect 24429 11656 24445 11720
rect 24509 11656 24525 11720
rect 24589 11656 24597 11720
rect 24277 10632 24597 11656
rect 24277 10568 24285 10632
rect 24349 10568 24365 10632
rect 24429 10568 24445 10632
rect 24509 10568 24525 10632
rect 24589 10568 24597 10632
rect 24277 9544 24597 10568
rect 24277 9480 24285 9544
rect 24349 9480 24365 9544
rect 24429 9480 24445 9544
rect 24509 9480 24525 9544
rect 24589 9480 24597 9544
rect 24277 8456 24597 9480
rect 24277 8392 24285 8456
rect 24349 8392 24365 8456
rect 24429 8392 24445 8456
rect 24509 8392 24525 8456
rect 24589 8392 24597 8456
rect 24277 7368 24597 8392
rect 24277 7304 24285 7368
rect 24349 7304 24365 7368
rect 24429 7304 24445 7368
rect 24509 7304 24525 7368
rect 24589 7304 24597 7368
rect 24277 6280 24597 7304
rect 24277 6216 24285 6280
rect 24349 6216 24365 6280
rect 24429 6216 24445 6280
rect 24509 6216 24525 6280
rect 24589 6216 24597 6280
rect 24277 5192 24597 6216
rect 24277 5128 24285 5192
rect 24349 5128 24365 5192
rect 24429 5128 24445 5192
rect 24509 5128 24525 5192
rect 24589 5128 24597 5192
rect 24277 4104 24597 5128
rect 24277 4040 24285 4104
rect 24349 4040 24365 4104
rect 24429 4040 24445 4104
rect 24509 4040 24525 4104
rect 24589 4040 24597 4104
rect 24277 3016 24597 4040
rect 24277 2952 24285 3016
rect 24349 2952 24365 3016
rect 24429 2952 24445 3016
rect 24509 2952 24525 3016
rect 24589 2952 24597 3016
rect 24277 1928 24597 2952
rect 24277 1864 24285 1928
rect 24349 1864 24365 1928
rect 24429 1864 24445 1928
rect 24509 1864 24525 1928
rect 24589 1864 24597 1928
rect 24277 1848 24597 1864
<< via4 >>
rect 6046 21022 6282 21258
rect 10830 20342 11066 20578
rect 21134 21022 21370 21258
rect 23894 20564 23980 20578
rect 23980 20564 24044 20578
rect 24044 20564 24130 20578
rect 23894 20342 24130 20564
<< metal5 >>
rect 6004 21258 21412 21300
rect 6004 21022 6046 21258
rect 6282 21022 21134 21258
rect 21370 21022 21412 21258
rect 6004 20980 21412 21022
rect 10788 20578 24172 20620
rect 10788 20342 10830 20578
rect 11066 20342 23894 20578
rect 24130 20342 24172 20578
rect 10788 20300 24172 20342
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2440
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2440
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2440
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 3956 0 1 2440
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2440
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2440
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_32
timestamp 1586364061
transform 1 0 4048 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2440
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_44
timestamp 1586364061
transform 1 0 5152 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_56
timestamp 1586364061
transform 1 0 6256 0 1 2440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2440
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_68
timestamp 1586364061
transform 1 0 7360 0 1 2440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2440
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 9568 0 1 2440
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2440
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_93
timestamp 1586364061
transform 1 0 9660 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2440
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2440
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_129
timestamp 1586364061
transform 1 0 12972 0 1 2440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2440
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 15180 0 1 2440
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2440
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_141
timestamp 1586364061
transform 1 0 14076 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_154 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 1 2440
box -38 -48 774 592
use scs8hd_buf_2  _72_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16100 0 1 2440
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__72__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16652 0 1 2440
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2440
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_162 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16008 0 1 2440
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_167 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16468 0 1 2440
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2440
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2440
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_183
timestamp 1586364061
transform 1 0 17940 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_195
timestamp 1586364061
transform 1 0 19044 0 1 2440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2440
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 20792 0 1 2440
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2440
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_207
timestamp 1586364061
transform 1 0 20148 0 1 2440
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_213
timestamp 1586364061
transform 1 0 20700 0 1 2440
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_215
timestamp 1586364061
transform 1 0 20884 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_227
timestamp 1586364061
transform 1 0 21988 0 1 2440
box -38 -48 1142 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 24564 0 1 2440
box -38 -48 406 592
use scs8hd_buf_2  _74_
timestamp 1586364061
transform 1 0 24564 0 -1 2440
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2440
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2440
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2440
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_239
timestamp 1586364061
transform 1 0 23092 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_251
timestamp 1586364061
transform 1 0 24196 0 1 2440
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_259
timestamp 1586364061
transform 1 0 24932 0 1 2440
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2440
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__74__A
timestamp 1586364061
transform 1 0 25116 0 -1 2440
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 25116 0 1 2440
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2440
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2440
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 26404 0 1 2440
box -38 -48 130 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2440
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2440
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_263
timestamp 1586364061
transform 1 0 25300 0 1 2440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2440
box -38 -48 1142 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3528
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_39
timestamp 1586364061
transform 1 0 4692 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_51
timestamp 1586364061
transform 1 0 5796 0 -1 3528
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_59
timestamp 1586364061
transform 1 0 6532 0 -1 3528
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 6716 0 -1 3528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_62
timestamp 1586364061
transform 1 0 6808 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_74
timestamp 1586364061
transform 1 0 7912 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_86
timestamp 1586364061
transform 1 0 9016 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_98
timestamp 1586364061
transform 1 0 10120 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 12328 0 -1 3528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_123
timestamp 1586364061
transform 1 0 12420 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_147
timestamp 1586364061
transform 1 0 14628 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_159
timestamp 1586364061
transform 1 0 15732 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 17940 0 -1 3528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_196
timestamp 1586364061
transform 1 0 19136 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_208
timestamp 1586364061
transform 1 0 20240 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_220
timestamp 1586364061
transform 1 0 21344 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 23552 0 -1 3528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_245
timestamp 1586364061
transform 1 0 23644 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_257
timestamp 1586364061
transform 1 0 24748 0 -1 3528
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3528
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_269
timestamp 1586364061
transform 1 0 25852 0 -1 3528
box -38 -48 774 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3528
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 1 3528
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3528
box -38 -48 406 592
use scs8hd_decap_12  FILLER_3_32
timestamp 1586364061
transform 1 0 4048 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_44
timestamp 1586364061
transform 1 0 5152 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_68
timestamp 1586364061
transform 1 0 7360 0 1 3528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 1 3528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_129
timestamp 1586364061
transform 1 0 12972 0 1 3528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 1 3528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_141
timestamp 1586364061
transform 1 0 14076 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_154
timestamp 1586364061
transform 1 0 15272 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_166
timestamp 1586364061
transform 1 0 16376 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_190
timestamp 1586364061
transform 1 0 18584 0 1 3528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 1 3528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_202
timestamp 1586364061
transform 1 0 19688 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_215
timestamp 1586364061
transform 1 0 20884 0 1 3528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3528
box -38 -48 1142 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 24564 0 1 3528
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 24380 0 1 3528
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3528
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_3_251
timestamp 1586364061
transform 1 0 24196 0 1 3528
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3528
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 26404 0 1 3528
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 25116 0 1 3528
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_259
timestamp 1586364061
transform 1 0 24932 0 1 3528
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_263
timestamp 1586364061
transform 1 0 25300 0 1 3528
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3528
box -38 -48 130 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4616
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_39
timestamp 1586364061
transform 1 0 4692 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4616
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4616
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 6716 0 -1 4616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_62
timestamp 1586364061
transform 1 0 6808 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_74
timestamp 1586364061
transform 1 0 7912 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_86
timestamp 1586364061
transform 1 0 9016 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_98
timestamp 1586364061
transform 1 0 10120 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 12328 0 -1 4616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_135
timestamp 1586364061
transform 1 0 13524 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_159
timestamp 1586364061
transform 1 0 15732 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_171
timestamp 1586364061
transform 1 0 16836 0 -1 4616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 17940 0 -1 4616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_184
timestamp 1586364061
transform 1 0 18032 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_196
timestamp 1586364061
transform 1 0 19136 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_208
timestamp 1586364061
transform 1 0 20240 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_220
timestamp 1586364061
transform 1 0 21344 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4616
box -38 -48 1142 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 24564 0 -1 4616
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 23552 0 -1 4616
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_245
timestamp 1586364061
transform 1 0 23644 0 -1 4616
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_253
timestamp 1586364061
transform 1 0 24380 0 -1 4616
box -38 -48 222 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4616
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4616
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_271
timestamp 1586364061
transform 1 0 26036 0 -1 4616
box -38 -48 590 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4616
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 3956 0 1 4616
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4616
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_44
timestamp 1586364061
transform 1 0 5152 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_56
timestamp 1586364061
transform 1 0 6256 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_68
timestamp 1586364061
transform 1 0 7360 0 1 4616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 9568 0 1 4616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_80
timestamp 1586364061
transform 1 0 8464 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_93
timestamp 1586364061
transform 1 0 9660 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_129
timestamp 1586364061
transform 1 0 12972 0 1 4616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 15180 0 1 4616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_141
timestamp 1586364061
transform 1 0 14076 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_190
timestamp 1586364061
transform 1 0 18584 0 1 4616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 20792 0 1 4616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_202
timestamp 1586364061
transform 1 0 19688 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_215
timestamp 1586364061
transform 1 0 20884 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_227
timestamp 1586364061
transform 1 0 21988 0 1 4616
box -38 -48 1142 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 24564 0 1 4616
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_239
timestamp 1586364061
transform 1 0 23092 0 1 4616
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_251
timestamp 1586364061
transform 1 0 24196 0 1 4616
box -38 -48 406 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4616
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 26404 0 1 4616
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 25116 0 1 4616
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_259
timestamp 1586364061
transform 1 0 24932 0 1 4616
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_263
timestamp 1586364061
transform 1 0 25300 0 1 4616
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4616
box -38 -48 130 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5704
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5704
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 3956 0 1 5704
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_39
timestamp 1586364061
transform 1 0 4692 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5704
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5704
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5704
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_44
timestamp 1586364061
transform 1 0 5152 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 6716 0 -1 5704
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_74
timestamp 1586364061
transform 1 0 7912 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_68
timestamp 1586364061
transform 1 0 7360 0 1 5704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 9568 0 1 5704
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_98
timestamp 1586364061
transform 1 0 10120 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_93
timestamp 1586364061
transform 1 0 9660 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 12328 0 -1 5704
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_135
timestamp 1586364061
transform 1 0 13524 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_129
timestamp 1586364061
transform 1 0 12972 0 1 5704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 15180 0 1 5704
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_147
timestamp 1586364061
transform 1 0 14628 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_141
timestamp 1586364061
transform 1 0 14076 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_154
timestamp 1586364061
transform 1 0 15272 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_159
timestamp 1586364061
transform 1 0 15732 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_171
timestamp 1586364061
transform 1 0 16836 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 17940 0 -1 5704
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_184
timestamp 1586364061
transform 1 0 18032 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_196
timestamp 1586364061
transform 1 0 19136 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_190
timestamp 1586364061
transform 1 0 18584 0 1 5704
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_198
timestamp 1586364061
transform 1 0 19320 0 1 5704
box -38 -48 130 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 19596 0 1 5704
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 20792 0 1 5704
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 20332 0 1 5704
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 19412 0 1 5704
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_208
timestamp 1586364061
transform 1 0 20240 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_205
timestamp 1586364061
transform 1 0 19964 0 1 5704
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_211
timestamp 1586364061
transform 1 0 20516 0 1 5704
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_215
timestamp 1586364061
transform 1 0 20884 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_220
timestamp 1586364061
transform 1 0 21344 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 23552 0 -1 5704
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_245
timestamp 1586364061
transform 1 0 23644 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_257
timestamp 1586364061
transform 1 0 24748 0 -1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_239
timestamp 1586364061
transform 1 0 23092 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_251
timestamp 1586364061
transform 1 0 24196 0 1 5704
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5704
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5704
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 26404 0 1 5704
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_269
timestamp 1586364061
transform 1 0 25852 0 -1 5704
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5704
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_276
timestamp 1586364061
transform 1 0 26496 0 1 5704
box -38 -48 130 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 6792
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_39
timestamp 1586364061
transform 1 0 4692 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 6792
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_59
timestamp 1586364061
transform 1 0 6532 0 -1 6792
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 6716 0 -1 6792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_98
timestamp 1586364061
transform 1 0 10120 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 6792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 12328 0 -1 6792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_147
timestamp 1586364061
transform 1 0 14628 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_159
timestamp 1586364061
transform 1 0 15732 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_171
timestamp 1586364061
transform 1 0 16836 0 -1 6792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 17940 0 -1 6792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_184
timestamp 1586364061
transform 1 0 18032 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 6792
box -38 -48 1142 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 20332 0 -1 6792
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_208
timestamp 1586364061
transform 1 0 20240 0 -1 6792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_225
timestamp 1586364061
transform 1 0 21804 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_237
timestamp 1586364061
transform 1 0 22908 0 -1 6792
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 23552 0 -1 6792
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_243
timestamp 1586364061
transform 1 0 23460 0 -1 6792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_245
timestamp 1586364061
transform 1 0 23644 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_257
timestamp 1586364061
transform 1 0 24748 0 -1 6792
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 6792
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_269
timestamp 1586364061
transform 1 0 25852 0 -1 6792
box -38 -48 774 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 6792
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 6792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 3956 0 1 6792
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 6792
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_32
timestamp 1586364061
transform 1 0 4048 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_68
timestamp 1586364061
transform 1 0 7360 0 1 6792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 9568 0 1 6792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_80
timestamp 1586364061
transform 1 0 8464 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_93
timestamp 1586364061
transform 1 0 9660 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_105
timestamp 1586364061
transform 1 0 10764 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_129
timestamp 1586364061
transform 1 0 12972 0 1 6792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 15180 0 1 6792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_141
timestamp 1586364061
transform 1 0 14076 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_166
timestamp 1586364061
transform 1 0 16376 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_190
timestamp 1586364061
transform 1 0 18584 0 1 6792
box -38 -48 1142 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 20976 0 1 6792
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 20792 0 1 6792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_202
timestamp 1586364061
transform 1 0 19688 0 1 6792
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 6792
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 21528 0 1 6792
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 6792
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_224
timestamp 1586364061
transform 1 0 21712 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 6792
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 24564 0 1 6792
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_248
timestamp 1586364061
transform 1 0 23920 0 1 6792
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 6792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 6792
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 6792
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 26404 0 1 6792
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 6792
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26496 0 1 6792
box -38 -48 130 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 7880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_39
timestamp 1586364061
transform 1 0 4692 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_51
timestamp 1586364061
transform 1 0 5796 0 -1 7880
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 7880
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 -1 7880
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_62
timestamp 1586364061
transform 1 0 6808 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_86
timestamp 1586364061
transform 1 0 9016 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_98
timestamp 1586364061
transform 1 0 10120 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 7880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 -1 7880
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_135
timestamp 1586364061
transform 1 0 13524 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_159
timestamp 1586364061
transform 1 0 15732 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_171
timestamp 1586364061
transform 1 0 16836 0 -1 7880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 -1 7880
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_184
timestamp 1586364061
transform 1 0 18032 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_220
timestamp 1586364061
transform 1 0 21344 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_232
timestamp 1586364061
transform 1 0 22448 0 -1 7880
box -38 -48 1142 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 24564 0 -1 7880
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 23552 0 -1 7880
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_245
timestamp 1586364061
transform 1 0 23644 0 -1 7880
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 7880
box -38 -48 222 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 7880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_259
timestamp 1586364061
transform 1 0 24932 0 -1 7880
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 7880
box -38 -48 590 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 7880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 7880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 1 7880
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 7880
box -38 -48 406 592
use scs8hd_decap_12  FILLER_11_32
timestamp 1586364061
transform 1 0 4048 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_44
timestamp 1586364061
transform 1 0 5152 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_68
timestamp 1586364061
transform 1 0 7360 0 1 7880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 1 7880
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_129
timestamp 1586364061
transform 1 0 12972 0 1 7880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 1 7880
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_141
timestamp 1586364061
transform 1 0 14076 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_166
timestamp 1586364061
transform 1 0 16376 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_190
timestamp 1586364061
transform 1 0 18584 0 1 7880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 1 7880
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_202
timestamp 1586364061
transform 1 0 19688 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_215
timestamp 1586364061
transform 1 0 20884 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 7880
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 24380 0 1 7880
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_239
timestamp 1586364061
transform 1 0 23092 0 1 7880
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_11_251
timestamp 1586364061
transform 1 0 24196 0 1 7880
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_255
timestamp 1586364061
transform 1 0 24564 0 1 7880
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 7880
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 1 7880
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_267
timestamp 1586364061
transform 1 0 25668 0 1 7880
box -38 -48 774 592
use scs8hd_fill_1  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 7880
box -38 -48 130 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 8968
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_39
timestamp 1586364061
transform 1 0 4692 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 8968
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 8968
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 6716 0 -1 8968
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_98
timestamp 1586364061
transform 1 0 10120 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 8968
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 12328 0 -1 8968
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_123
timestamp 1586364061
transform 1 0 12420 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_135
timestamp 1586364061
transform 1 0 13524 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_159
timestamp 1586364061
transform 1 0 15732 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_171
timestamp 1586364061
transform 1 0 16836 0 -1 8968
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 17940 0 -1 8968
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_184
timestamp 1586364061
transform 1 0 18032 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_196
timestamp 1586364061
transform 1 0 19136 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_208
timestamp 1586364061
transform 1 0 20240 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_220
timestamp 1586364061
transform 1 0 21344 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_232
timestamp 1586364061
transform 1 0 22448 0 -1 8968
box -38 -48 1142 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 24380 0 -1 8968
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 23552 0 -1 8968
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_245
timestamp 1586364061
transform 1 0 23644 0 -1 8968
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_257
timestamp 1586364061
transform 1 0 24748 0 -1 8968
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 8968
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_269
timestamp 1586364061
transform 1 0 25852 0 -1 8968
box -38 -48 774 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 8968
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10056
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 1 8968
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 8968
box -38 -48 406 592
use scs8hd_decap_12  FILLER_13_32
timestamp 1586364061
transform 1 0 4048 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_39
timestamp 1586364061
transform 1 0 4692 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_51
timestamp 1586364061
transform 1 0 5796 0 -1 10056
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10056
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 6716 0 -1 10056
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_68
timestamp 1586364061
transform 1 0 7360 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_74
timestamp 1586364061
transform 1 0 7912 0 -1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 1 8968
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_86
timestamp 1586364061
transform 1 0 9016 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_98
timestamp 1586364061
transform 1 0 10120 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_110
timestamp 1586364061
transform 1 0 11224 0 -1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 12328 0 -1 10056
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_123
timestamp 1586364061
transform 1 0 12420 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 15180 0 1 8968
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_159
timestamp 1586364061
transform 1 0 15732 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_171
timestamp 1586364061
transform 1 0 16836 0 -1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 17940 0 -1 10056
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_190
timestamp 1586364061
transform 1 0 18584 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_184
timestamp 1586364061
transform 1 0 18032 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_196
timestamp 1586364061
transform 1 0 19136 0 -1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 20792 0 1 8968
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_202
timestamp 1586364061
transform 1 0 19688 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_215
timestamp 1586364061
transform 1 0 20884 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_220
timestamp 1586364061
transform 1 0 21344 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_245
timestamp 1586364061
transform 1 0 23644 0 -1 10056
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 8968
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 8968
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 23552 0 -1 10056
box -38 -48 130 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 23736 0 1 8968
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_253
timestamp 1586364061
transform 1 0 24380 0 -1 10056
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 8968
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_250
timestamp 1586364061
transform 1 0 24104 0 1 8968
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 24288 0 1 8968
box -38 -48 222 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 24564 0 -1 10056
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 24656 0 1 8968
box -38 -48 222 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 8968
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10056
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 26404 0 1 8968
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 8968
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_13_270
timestamp 1586364061
transform 1 0 25944 0 1 8968
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_274
timestamp 1586364061
transform 1 0 26312 0 1 8968
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 8968
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10056
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10056
box -38 -48 590 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10056
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 3956 0 1 10056
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10056
box -38 -48 406 592
use scs8hd_decap_12  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_44
timestamp 1586364061
transform 1 0 5152 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_68
timestamp 1586364061
transform 1 0 7360 0 1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 9568 0 1 10056
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_129
timestamp 1586364061
transform 1 0 12972 0 1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 15180 0 1 10056
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_141
timestamp 1586364061
transform 1 0 14076 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_190
timestamp 1586364061
transform 1 0 18584 0 1 10056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 20792 0 1 10056
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_215
timestamp 1586364061
transform 1 0 20884 0 1 10056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_227
timestamp 1586364061
transform 1 0 21988 0 1 10056
box -38 -48 1142 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 24564 0 1 10056
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 24380 0 1 10056
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_239
timestamp 1586364061
transform 1 0 23092 0 1 10056
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_15_251
timestamp 1586364061
transform 1 0 24196 0 1 10056
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10056
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 26404 0 1 10056
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 25116 0 1 10056
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10056
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10056
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10056
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11144
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_39
timestamp 1586364061
transform 1 0 4692 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_51
timestamp 1586364061
transform 1 0 5796 0 -1 11144
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11144
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 -1 11144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_98
timestamp 1586364061
transform 1 0 10120 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_110
timestamp 1586364061
transform 1 0 11224 0 -1 11144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 -1 11144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_123
timestamp 1586364061
transform 1 0 12420 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_135
timestamp 1586364061
transform 1 0 13524 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_147
timestamp 1586364061
transform 1 0 14628 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_159
timestamp 1586364061
transform 1 0 15732 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 17940 0 -1 11144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_184
timestamp 1586364061
transform 1 0 18032 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_196
timestamp 1586364061
transform 1 0 19136 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_208
timestamp 1586364061
transform 1 0 20240 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_220
timestamp 1586364061
transform 1 0 21344 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_232
timestamp 1586364061
transform 1 0 22448 0 -1 11144
box -38 -48 1142 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 24564 0 -1 11144
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 23552 0 -1 11144
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_245
timestamp 1586364061
transform 1 0 23644 0 -1 11144
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_253
timestamp 1586364061
transform 1 0 24380 0 -1 11144
box -38 -48 222 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11144
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_259
timestamp 1586364061
transform 1 0 24932 0 -1 11144
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11144
box -38 -48 590 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11144
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 1 11144
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11144
box -38 -48 406 592
use scs8hd_decap_12  FILLER_17_32
timestamp 1586364061
transform 1 0 4048 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_44
timestamp 1586364061
transform 1 0 5152 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 1 11144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_129
timestamp 1586364061
transform 1 0 12972 0 1 11144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 1 11144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_154
timestamp 1586364061
transform 1 0 15272 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11144
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11144
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 1 11144
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18584 0 1 11144
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18952 0 1 11144
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_188
timestamp 1586364061
transform 1 0 18400 0 1 11144
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_192
timestamp 1586364061
transform 1 0 18768 0 1 11144
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 1 11144
box -38 -48 130 592
use scs8hd_decap_6  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11144
box -38 -48 590 592
use scs8hd_decap_12  FILLER_17_215
timestamp 1586364061
transform 1 0 20884 0 1 11144
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22540 0 1 11144
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_227
timestamp 1586364061
transform 1 0 21988 0 1 11144
box -38 -48 590 592
use scs8hd_decap_8  FILLER_17_235
timestamp 1586364061
transform 1 0 22724 0 1 11144
box -38 -48 774 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 24564 0 1 11144
box -38 -48 406 592
use scs8hd_buf_1  mux_right_track_0.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23552 0 1 11144
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 24380 0 1 11144
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24012 0 1 11144
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_243
timestamp 1586364061
transform 1 0 23460 0 1 11144
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_247
timestamp 1586364061
transform 1 0 23828 0 1 11144
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_251
timestamp 1586364061
transform 1 0 24196 0 1 11144
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11144
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 26404 0 1 11144
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 25116 0 1 11144
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24932 0 1 11144
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_263
timestamp 1586364061
transform 1 0 25300 0 1 11144
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11144
box -38 -48 130 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12232
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_39
timestamp 1586364061
transform 1 0 4692 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_51
timestamp 1586364061
transform 1 0 5796 0 -1 12232
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_59
timestamp 1586364061
transform 1 0 6532 0 -1 12232
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 6716 0 -1 12232
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_86
timestamp 1586364061
transform 1 0 9016 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_98
timestamp 1586364061
transform 1 0 10120 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12232
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 12328 0 -1 12232
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_147
timestamp 1586364061
transform 1 0 14628 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_159
timestamp 1586364061
transform 1 0 15732 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12232
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18216 0 -1 12232
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 17940 0 -1 12232
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12232
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_195
timestamp 1586364061
transform 1 0 19044 0 -1 12232
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19412 0 -1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20884 0 -1 12232
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_201
timestamp 1586364061
transform 1 0 19596 0 -1 12232
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12232
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_217
timestamp 1586364061
transform 1 0 21068 0 -1 12232
box -38 -48 774 592
use scs8hd_buf_1  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22540 0 -1 12232
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 -1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22264 0 -1 12232
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_225
timestamp 1586364061
transform 1 0 21804 0 -1 12232
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12232
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_232
timestamp 1586364061
transform 1 0 22448 0 -1 12232
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_236
timestamp 1586364061
transform 1 0 22816 0 -1 12232
box -38 -48 774 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 24564 0 -1 12232
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 23552 0 -1 12232
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_245
timestamp 1586364061
transform 1 0 23644 0 -1 12232
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_253
timestamp 1586364061
transform 1 0 24380 0 -1 12232
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12232
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12232
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12232
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 13320
box -38 -48 1786 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12232
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13320
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 1564 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1932 0 1 12232
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12232
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12232
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12232
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 3956 0 1 12232
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12232
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_22
timestamp 1586364061
transform 1 0 3128 0 -1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_34
timestamp 1586364061
transform 1 0 4232 0 -1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_44
timestamp 1586364061
transform 1 0 5152 0 1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13320
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_58
timestamp 1586364061
transform 1 0 6440 0 -1 13320
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 6716 0 -1 13320
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_68
timestamp 1586364061
transform 1 0 7360 0 1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13320
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 9568 0 1 12232
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_80
timestamp 1586364061
transform 1 0 8464 0 1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_98
timestamp 1586364061
transform 1 0 10120 0 -1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_105
timestamp 1586364061
transform 1 0 10764 0 1 12232
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12232
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_110
timestamp 1586364061
transform 1 0 11224 0 -1 13320
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_127
timestamp 1586364061
transform 1 0 12788 0 -1 13320
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_123
timestamp 1586364061
transform 1 0 12420 0 -1 13320
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_125
timestamp 1586364061
transform 1 0 12604 0 1 12232
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12880 0 1 12232
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12328 0 -1 13320
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 13320
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12232
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13616 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13248 0 1 12232
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12232
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15456 0 -1 13320
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 15180 0 1 12232
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 15272 0 -1 13320
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_150
timestamp 1586364061
transform 1 0 14904 0 1 12232
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12232
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12232
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13320
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_153
timestamp 1586364061
transform 1 0 15180 0 -1 13320
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15824 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16192 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17480 0 1 12232
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12232
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_166
timestamp 1586364061
transform 1 0 16376 0 1 12232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13320
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_177
timestamp 1586364061
transform 1 0 17388 0 -1 13320
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 -1 13320
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17848 0 1 12232
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 17940 0 -1 13320
box -38 -48 130 592
use scs8hd_conb_1  _22_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18032 0 -1 13320
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_195
timestamp 1586364061
transform 1 0 19044 0 -1 13320
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_191
timestamp 1586364061
transform 1 0 18676 0 -1 13320
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18860 0 -1 13320
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18492 0 -1 13320
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 12232
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19412 0 -1 13320
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 1 12232
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 20792 0 1 12232
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20608 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19964 0 1 12232
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12232
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12232
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_211
timestamp 1586364061
transform 1 0 20516 0 1 12232
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13320
box -38 -48 774 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21896 0 -1 13320
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22816 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22908 0 -1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12232
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_238
timestamp 1586364061
transform 1 0 23000 0 1 12232
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_235
timestamp 1586364061
transform 1 0 22724 0 -1 13320
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_245
timestamp 1586364061
transform 1 0 23644 0 -1 13320
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_243
timestamp 1586364061
transform 1 0 23460 0 -1 13320
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13320
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_242
timestamp 1586364061
transform 1 0 23368 0 1 12232
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 23552 0 -1 13320
box -38 -48 130 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 23460 0 1 12232
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_253
timestamp 1586364061
transform 1 0 24380 0 -1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_251
timestamp 1586364061
transform 1 0 24196 0 1 12232
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_247
timestamp 1586364061
transform 1 0 23828 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 24380 0 1 12232
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 24012 0 1 12232
box -38 -48 222 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 24564 0 1 12232
box -38 -48 406 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 24564 0 -1 13320
box -38 -48 406 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12232
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13320
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 26404 0 1 12232
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 25116 0 1 12232
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12232
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12232
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_19_276
timestamp 1586364061
transform 1 0 26496 0 1 12232
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13320
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13320
box -38 -48 590 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13320
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13320
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 1 13320
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13320
box -38 -48 406 592
use scs8hd_decap_12  FILLER_21_32
timestamp 1586364061
transform 1 0 4048 0 1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_44
timestamp 1586364061
transform 1 0 5152 0 1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_56
timestamp 1586364061
transform 1 0 6256 0 1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_68
timestamp 1586364061
transform 1 0 7360 0 1 13320
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 1 13320
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13320
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12052 0 1 13320
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11684 0 1 13320
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_105
timestamp 1586364061
transform 1 0 10764 0 1 13320
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_117
timestamp 1586364061
transform 1 0 11868 0 1 13320
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12236 0 1 13320
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 1 13320
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 15180 0 1 13320
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14996 0 1 13320
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14168 0 1 13320
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14536 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_140
timestamp 1586364061
transform 1 0 13984 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_144
timestamp 1586364061
transform 1 0 14352 0 1 13320
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_148
timestamp 1586364061
transform 1 0 14720 0 1 13320
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17204 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_173
timestamp 1586364061
transform 1 0 17020 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_177
timestamp 1586364061
transform 1 0 17388 0 1 13320
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17756 0 1 13320
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17572 0 1 13320
box -38 -48 222 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 21160 0 1 13320
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 20792 0 1 13320
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20608 0 1 13320
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 1 13320
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_200
timestamp 1586364061
transform 1 0 19504 0 1 13320
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_210
timestamp 1586364061
transform 1 0 20424 0 1 13320
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_215
timestamp 1586364061
transform 1 0 20884 0 1 13320
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22172 0 1 13320
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21988 0 1 13320
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21620 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_221
timestamp 1586364061
transform 1 0 21436 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_225
timestamp 1586364061
transform 1 0 21804 0 1 13320
box -38 -48 222 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 24656 0 1 13320
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 24104 0 1 13320
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24472 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_248
timestamp 1586364061
transform 1 0 23920 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_252
timestamp 1586364061
transform 1 0 24288 0 1 13320
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13320
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 26404 0 1 13320
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 25208 0 1 13320
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_260
timestamp 1586364061
transform 1 0 25024 0 1 13320
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_264
timestamp 1586364061
transform 1 0 25392 0 1 13320
box -38 -48 774 592
use scs8hd_decap_3  FILLER_21_272
timestamp 1586364061
transform 1 0 26128 0 1 13320
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13320
box -38 -48 130 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_39
timestamp 1586364061
transform 1 0 4692 0 -1 14408
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14408
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_59
timestamp 1586364061
transform 1 0 6532 0 -1 14408
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 6716 0 -1 14408
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_62
timestamp 1586364061
transform 1 0 6808 0 -1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_74
timestamp 1586364061
transform 1 0 7912 0 -1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_98
timestamp 1586364061
transform 1 0 10120 0 -1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14408
box -38 -48 1142 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 12696 0 -1 14408
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13708 0 -1 14408
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 12328 0 -1 14408
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14408
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14408
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_156
timestamp 1586364061
transform 1 0 15456 0 -1 14408
box -38 -48 774 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 16192 0 -1 14408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_167
timestamp 1586364061
transform 1 0 16468 0 -1 14408
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 -1 14408
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 17940 0 -1 14408
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_179
timestamp 1586364061
transform 1 0 17572 0 -1 14408
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_193
timestamp 1586364061
transform 1 0 18860 0 -1 14408
box -38 -48 1142 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20976 0 -1 14408
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_205
timestamp 1586364061
transform 1 0 19964 0 -1 14408
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14408
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22540 0 -1 14408
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22172 0 -1 14408
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_225
timestamp 1586364061
transform 1 0 21804 0 -1 14408
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_231
timestamp 1586364061
transform 1 0 22356 0 -1 14408
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_236
timestamp 1586364061
transform 1 0 22816 0 -1 14408
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 -1 14408
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 23552 0 -1 14408
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_264
timestamp 1586364061
transform 1 0 25392 0 -1 14408
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14408
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14408
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 3956 0 1 14408
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14408
box -38 -48 406 592
use scs8hd_decap_12  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_44
timestamp 1586364061
transform 1 0 5152 0 1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_68
timestamp 1586364061
transform 1 0 7360 0 1 14408
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 9568 0 1 14408
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14408
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11960 0 1 14408
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_105
timestamp 1586364061
transform 1 0 10764 0 1 14408
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14408
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12880 0 1 14408
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12696 0 1 14408
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12328 0 1 14408
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_120
timestamp 1586364061
transform 1 0 12144 0 1 14408
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_124
timestamp 1586364061
transform 1 0 12512 0 1 14408
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_137
timestamp 1586364061
transform 1 0 13708 0 1 14408
box -38 -48 590 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 1 14408
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 15180 0 1 14408
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 1 14408
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 1 14408
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14260 0 1 14408
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_145
timestamp 1586364061
transform 1 0 14444 0 1 14408
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14408
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 17020 0 1 14408
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17480 0 1 14408
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14408
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14408
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_176
timestamp 1586364061
transform 1 0 17296 0 1 14408
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 14408
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19136 0 1 14408
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18492 0 1 14408
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14408
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14408
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14408
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_195
timestamp 1586364061
transform 1 0 19044 0 1 14408
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14408
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 20792 0 1 14408
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19504 0 1 14408
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_202
timestamp 1586364061
transform 1 0 19688 0 1 14408
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_23_215
timestamp 1586364061
transform 1 0 20884 0 1 14408
box -38 -48 406 592
use scs8hd_buf_1  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21252 0 1 14408
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 22908 0 1 14408
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21712 0 1 14408
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_222
timestamp 1586364061
transform 1 0 21528 0 1 14408
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_226
timestamp 1586364061
transform 1 0 21896 0 1 14408
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14408
box -38 -48 314 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 24564 0 1 14408
box -38 -48 406 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 23460 0 1 14408
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 24012 0 1 14408
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24380 0 1 14408
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 23276 0 1 14408
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_239
timestamp 1586364061
transform 1 0 23092 0 1 14408
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_247
timestamp 1586364061
transform 1 0 23828 0 1 14408
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_251
timestamp 1586364061
transform 1 0 24196 0 1 14408
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14408
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 26404 0 1 14408
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 25208 0 1 14408
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_259
timestamp 1586364061
transform 1 0 24932 0 1 14408
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_264
timestamp 1586364061
transform 1 0 25392 0 1 14408
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_272
timestamp 1586364061
transform 1 0 26128 0 1 14408
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14408
box -38 -48 130 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15496
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_39
timestamp 1586364061
transform 1 0 4692 0 -1 15496
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_51
timestamp 1586364061
transform 1 0 5796 0 -1 15496
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15496
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 -1 15496
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_86
timestamp 1586364061
transform 1 0 9016 0 -1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_98
timestamp 1586364061
transform 1 0 10120 0 -1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15496
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12420 0 -1 15496
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 -1 15496
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12880 0 -1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15496
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15496
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14628 0 -1 15496
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15272 0 -1 15496
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15496
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_146
timestamp 1586364061
transform 1 0 14536 0 -1 15496
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15496
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_156
timestamp 1586364061
transform 1 0 15456 0 -1 15496
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17020 0 -1 15496
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15496
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_172
timestamp 1586364061
transform 1 0 16928 0 -1 15496
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_175
timestamp 1586364061
transform 1 0 17204 0 -1 15496
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19136 0 -1 15496
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 17940 0 -1 15496
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_184
timestamp 1586364061
transform 1 0 18032 0 -1 15496
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21068 0 -1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15496
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_219
timestamp 1586364061
transform 1 0 21252 0 -1 15496
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_231
timestamp 1586364061
transform 1 0 22356 0 -1 15496
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 -1 15496
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 23552 0 -1 15496
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 23368 0 -1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 24656 0 -1 15496
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15496
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_254
timestamp 1586364061
transform 1 0 24472 0 -1 15496
box -38 -48 222 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 25208 0 -1 15496
box -38 -48 406 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15496
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_258
timestamp 1586364061
transform 1 0 24840 0 -1 15496
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_266
timestamp 1586364061
transform 1 0 25576 0 -1 15496
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15496
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15496
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15496
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 3956 0 1 15496
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15496
box -38 -48 406 592
use scs8hd_decap_12  FILLER_25_32
timestamp 1586364061
transform 1 0 4048 0 1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_44
timestamp 1586364061
transform 1 0 5152 0 1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_68
timestamp 1586364061
transform 1 0 7360 0 1 15496
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 9568 0 1 15496
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_93
timestamp 1586364061
transform 1 0 9660 0 1 15496
box -38 -48 1142 592
use scs8hd_buf_1  mux_right_track_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12052 0 1 15496
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_105
timestamp 1586364061
transform 1 0 10764 0 1 15496
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12512 0 1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_122
timestamp 1586364061
transform 1 0 12328 0 1 15496
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15496
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15496
box -38 -48 222 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 15272 0 1 15496
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 1 15496
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 15180 0 1 15496
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14628 0 1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13984 0 1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14996 0 1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15496
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_157
timestamp 1586364061
transform 1 0 15548 0 1 15496
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17020 0 1 15496
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16836 0 1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_169
timestamp 1586364061
transform 1 0 16652 0 1 15496
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_192
timestamp 1586364061
transform 1 0 18768 0 1 15496
box -38 -48 774 592
use scs8hd_conb_1  _34_
timestamp 1586364061
transform 1 0 19780 0 1 15496
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 20884 0 1 15496
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 20792 0 1 15496
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19596 0 1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 20608 0 1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20240 0 1 15496
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_200
timestamp 1586364061
transform 1 0 19504 0 1 15496
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_206
timestamp 1586364061
transform 1 0 20056 0 1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 22908 0 1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_224
timestamp 1586364061
transform 1 0 21712 0 1 15496
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_228
timestamp 1586364061
transform 1 0 22080 0 1 15496
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15496
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23092 0 1 15496
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_25_262
timestamp 1586364061
transform 1 0 25208 0 1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 25024 0 1 15496
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_266
timestamp 1586364061
transform 1 0 25576 0 1 15496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 25392 0 1 15496
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_270
timestamp 1586364061
transform 1 0 25944 0 1 15496
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 25760 0 1 15496
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15496
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_274
timestamp 1586364061
transform 1 0 26312 0 1 15496
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 26404 0 1 15496
box -38 -48 130 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15496
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16584
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16584
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16584
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 3956 0 1 16584
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_39
timestamp 1586364061
transform 1 0 4692 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16584
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_32
timestamp 1586364061
transform 1 0 4048 0 1 16584
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16584
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_59
timestamp 1586364061
transform 1 0 6532 0 -1 16584
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16584
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 6716 0 -1 16584
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_68
timestamp 1586364061
transform 1 0 7360 0 1 16584
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 9568 0 1 16584
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_86
timestamp 1586364061
transform 1 0 9016 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_98
timestamp 1586364061
transform 1 0 10120 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_110
timestamp 1586364061
transform 1 0 11224 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16584
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 12328 0 -1 16584
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16584
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_129
timestamp 1586364061
transform 1 0 12972 0 1 16584
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16584
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_135
timestamp 1586364061
transform 1 0 13524 0 -1 16584
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13064 0 1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13616 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 16584
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 1 16584
box -38 -48 866 592
use scs8hd_decap_12  FILLER_26_123
timestamp 1586364061
transform 1 0 12420 0 -1 16584
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14076 0 -1 16584
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15272 0 1 16584
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 15180 0 1 16584
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14628 0 1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 1 16584
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_145
timestamp 1586364061
transform 1 0 14444 0 1 16584
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16584
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_167
timestamp 1586364061
transform 1 0 16468 0 1 16584
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_163
timestamp 1586364061
transform 1 0 16100 0 1 16584
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_164
timestamp 1586364061
transform 1 0 16192 0 -1 16584
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_160
timestamp 1586364061
transform 1 0 15824 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16008 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16284 0 1 16584
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16584
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_172
timestamp 1586364061
transform 1 0 16928 0 -1 16584
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17020 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16836 0 1 16584
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17020 0 1 16584
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 17940 0 -1 16584
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19044 0 1 16584
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_184
timestamp 1586364061
transform 1 0 18032 0 -1 16584
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_196
timestamp 1586364061
transform 1 0 19136 0 -1 16584
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_192
timestamp 1586364061
transform 1 0 18768 0 1 16584
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16584
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_205
timestamp 1586364061
transform 1 0 19964 0 1 16584
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_201
timestamp 1586364061
transform 1 0 19596 0 1 16584
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_200
timestamp 1586364061
transform 1 0 19504 0 -1 16584
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19412 0 1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20240 0 1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19780 0 1 16584
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20608 0 1 16584
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 20792 0 1 16584
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20884 0 1 16584
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19596 0 -1 16584
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_27_228
timestamp 1586364061
transform 1 0 22080 0 1 16584
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_224
timestamp 1586364061
transform 1 0 21712 0 1 16584
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_228
timestamp 1586364061
transform 1 0 22080 0 -1 16584
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16584
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_220
timestamp 1586364061
transform 1 0 21344 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21528 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21896 0 1 16584
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_236
timestamp 1586364061
transform 1 0 22816 0 -1 16584
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_232
timestamp 1586364061
transform 1 0 22448 0 -1 16584
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22448 0 1 16584
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 22632 0 1 16584
box -38 -48 866 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 22540 0 -1 16584
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_247
timestamp 1586364061
transform 1 0 23828 0 1 16584
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_243
timestamp 1586364061
transform 1 0 23460 0 1 16584
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_241
timestamp 1586364061
transform 1 0 23276 0 -1 16584
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23092 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23644 0 1 16584
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 23552 0 -1 16584
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 23644 0 -1 16584
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_254
timestamp 1586364061
transform 1 0 24472 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24656 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 24012 0 1 16584
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24196 0 1 16584
box -38 -48 866 592
use scs8hd_decap_8  FILLER_27_264
timestamp 1586364061
transform 1 0 25392 0 1 16584
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_260
timestamp 1586364061
transform 1 0 25024 0 1 16584
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_266
timestamp 1586364061
transform 1 0 25576 0 -1 16584
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_258
timestamp 1586364061
transform 1 0 24840 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 -1 16584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 25208 0 1 16584
box -38 -48 222 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 25208 0 -1 16584
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_272
timestamp 1586364061
transform 1 0 26128 0 1 16584
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16584
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 26404 0 1 16584
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16584
box -38 -48 130 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16584
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16584
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17672
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_39
timestamp 1586364061
transform 1 0 4692 0 -1 17672
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_51
timestamp 1586364061
transform 1 0 5796 0 -1 17672
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17672
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 6716 0 -1 17672
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_62
timestamp 1586364061
transform 1 0 6808 0 -1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17672
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_98
timestamp 1586364061
transform 1 0 10120 0 -1 17672
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11040 0 -1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17672
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17672
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 12328 0 -1 17672
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13616 0 -1 17672
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_123
timestamp 1586364061
transform 1 0 12420 0 -1 17672
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17672
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_138
timestamp 1586364061
transform 1 0 13800 0 -1 17672
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14260 0 -1 17672
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14076 0 -1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17112 0 -1 17672
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_162
timestamp 1586364061
transform 1 0 16008 0 -1 17672
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_176
timestamp 1586364061
transform 1 0 17296 0 -1 17672
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 17940 0 -1 17672
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18216 0 -1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 18584 0 -1 17672
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_182
timestamp 1586364061
transform 1 0 17848 0 -1 17672
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17672
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17672
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19780 0 -1 17672
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20884 0 -1 17672
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_200
timestamp 1586364061
transform 1 0 19504 0 -1 17672
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17672
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_217
timestamp 1586364061
transform 1 0 21068 0 -1 17672
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21344 0 -1 17672
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22356 0 -1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22724 0 -1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_229
timestamp 1586364061
transform 1 0 22172 0 -1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_233
timestamp 1586364061
transform 1 0 22540 0 -1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_237
timestamp 1586364061
transform 1 0 22908 0 -1 17672
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24104 0 -1 17672
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 23552 0 -1 17672
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23920 0 -1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23092 0 -1 17672
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_241
timestamp 1586364061
transform 1 0 23276 0 -1 17672
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_245
timestamp 1586364061
transform 1 0 23644 0 -1 17672
box -38 -48 314 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17672
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_269
timestamp 1586364061
transform 1 0 25852 0 -1 17672
box -38 -48 774 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17672
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17672
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 1 17672
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17672
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_44
timestamp 1586364061
transform 1 0 5152 0 1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_56
timestamp 1586364061
transform 1 0 6256 0 1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_68
timestamp 1586364061
transform 1 0 7360 0 1 17672
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 1 17672
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17672
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11040 0 1 17672
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10856 0 1 17672
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17672
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 1 17672
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 17672
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_127
timestamp 1586364061
transform 1 0 12788 0 1 17672
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_133
timestamp 1586364061
transform 1 0 13340 0 1 17672
box -38 -48 130 592
use scs8hd_buf_1  mux_right_track_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 1 17672
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 15180 0 1 17672
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 1 17672
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_145
timestamp 1586364061
transform 1 0 14444 0 1 17672
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_149
timestamp 1586364061
transform 1 0 14812 0 1 17672
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_152
timestamp 1586364061
transform 1 0 15088 0 1 17672
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_157
timestamp 1586364061
transform 1 0 15548 0 1 17672
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 17112 0 1 17672
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16928 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15732 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16100 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16468 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_161
timestamp 1586364061
transform 1 0 15916 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_165
timestamp 1586364061
transform 1 0 16284 0 1 17672
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_169
timestamp 1586364061
transform 1 0 16652 0 1 17672
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17672
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17672
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 20792 0 1 17672
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 20424 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21068 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20056 0 1 17672
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_205
timestamp 1586364061
transform 1 0 19964 0 1 17672
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_212
timestamp 1586364061
transform 1 0 20608 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_215
timestamp 1586364061
transform 1 0 20884 0 1 17672
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 22356 0 1 17672
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22172 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21436 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_219
timestamp 1586364061
transform 1 0 21252 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_223
timestamp 1586364061
transform 1 0 21620 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_227
timestamp 1586364061
transform 1 0 21988 0 1 17672
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23920 0 1 17672
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23736 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_244
timestamp 1586364061
transform 1 0 23552 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17672
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17672
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 26404 0 1 17672
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 24932 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 25300 0 1 17672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 25668 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_261
timestamp 1586364061
transform 1 0 25116 0 1 17672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_265
timestamp 1586364061
transform 1 0 25484 0 1 17672
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17672
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_276
timestamp 1586364061
transform 1 0 26496 0 1 17672
box -38 -48 130 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 18760
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 18760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 18760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 18760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_39
timestamp 1586364061
transform 1 0 4692 0 -1 18760
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_51
timestamp 1586364061
transform 1 0 5796 0 -1 18760
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_59
timestamp 1586364061
transform 1 0 6532 0 -1 18760
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 6716 0 -1 18760
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_62
timestamp 1586364061
transform 1 0 6808 0 -1 18760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_74
timestamp 1586364061
transform 1 0 7912 0 -1 18760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_86
timestamp 1586364061
transform 1 0 9016 0 -1 18760
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_98
timestamp 1586364061
transform 1 0 10120 0 -1 18760
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11132 0 -1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11500 0 -1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_104
timestamp 1586364061
transform 1 0 10672 0 -1 18760
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_111
timestamp 1586364061
transform 1 0 11316 0 -1 18760
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_115
timestamp 1586364061
transform 1 0 11684 0 -1 18760
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 12328 0 -1 18760
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12696 0 -1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13616 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 18760
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_123
timestamp 1586364061
transform 1 0 12420 0 -1 18760
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 18760
box -38 -48 774 592
use scs8hd_decap_6  FILLER_30_138
timestamp 1586364061
transform 1 0 13800 0 -1 18760
box -38 -48 590 592
use scs8hd_mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14904 0 -1 18760
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14444 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_144
timestamp 1586364061
transform 1 0 14352 0 -1 18760
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_147
timestamp 1586364061
transform 1 0 14628 0 -1 18760
box -38 -48 314 592
use scs8hd_conb_1  _35_
timestamp 1586364061
transform 1 0 16928 0 -1 18760
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15916 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_159
timestamp 1586364061
transform 1 0 15732 0 -1 18760
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 18760
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_171
timestamp 1586364061
transform 1 0 16836 0 -1 18760
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_175
timestamp 1586364061
transform 1 0 17204 0 -1 18760
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18032 0 -1 18760
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 17940 0 -1 18760
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19228 0 -1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17572 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_181
timestamp 1586364061
transform 1 0 17756 0 -1 18760
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 18760
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20424 0 -1 18760
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_199
timestamp 1586364061
transform 1 0 19412 0 -1 18760
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_207
timestamp 1586364061
transform 1 0 20148 0 -1 18760
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21988 0 -1 18760
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21436 0 -1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21804 0 -1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_219
timestamp 1586364061
transform 1 0 21252 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_223
timestamp 1586364061
transform 1 0 21620 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_236
timestamp 1586364061
transform 1 0 22816 0 -1 18760
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 -1 18760
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 23552 0 -1 18760
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24656 0 -1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_240
timestamp 1586364061
transform 1 0 23184 0 -1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_254
timestamp 1586364061
transform 1 0 24472 0 -1 18760
box -38 -48 222 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 25208 0 -1 18760
box -38 -48 406 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 18760
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_258
timestamp 1586364061
transform 1 0 24840 0 -1 18760
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_266
timestamp 1586364061
transform 1 0 25576 0 -1 18760
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 18760
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 18760
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 18760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 18760
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 3956 0 1 18760
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 18760
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 18760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 18760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 18760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_68
timestamp 1586364061
transform 1 0 7360 0 1 18760
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 9568 0 1 18760
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 18760
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 18760
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11132 0 1 18760
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_103
timestamp 1586364061
transform 1 0 10580 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_107
timestamp 1586364061
transform 1 0 10948 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 18760
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12696 0 1 18760
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12512 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_122
timestamp 1586364061
transform 1 0 12328 0 1 18760
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 1 18760
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 15180 0 1 18760
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14628 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_145
timestamp 1586364061
transform 1 0 14444 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17388 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 17020 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_167
timestamp 1586364061
transform 1 0 16468 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 18760
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 1 18760
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 17572 0 1 18760
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18676 0 1 18760
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_188
timestamp 1586364061
transform 1 0 18400 0 1 18760
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 18760
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 1 18760
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 20792 0 1 18760
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20608 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 20240 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_206
timestamp 1586364061
transform 1 0 20056 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 18760
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_234
timestamp 1586364061
transform 1 0 22632 0 1 18760
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23552 0 1 18760
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 24564 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23368 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 18760
box -38 -48 222 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 25116 0 1 18760
box -38 -48 406 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 18760
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 26404 0 1 18760
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24932 0 1 18760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 25668 0 1 18760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_265
timestamp 1586364061
transform 1 0 25484 0 1 18760
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 18760
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 18760
box -38 -48 130 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 19848
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_39
timestamp 1586364061
transform 1 0 4692 0 -1 19848
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_51
timestamp 1586364061
transform 1 0 5796 0 -1 19848
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 19848
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 -1 19848
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_62
timestamp 1586364061
transform 1 0 6808 0 -1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_86
timestamp 1586364061
transform 1 0 9016 0 -1 19848
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_98
timestamp 1586364061
transform 1 0 10120 0 -1 19848
box -38 -48 590 592
use scs8hd_mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 -1 19848
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11776 0 -1 19848
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 19848
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_114
timestamp 1586364061
transform 1 0 11592 0 -1 19848
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_118
timestamp 1586364061
transform 1 0 11960 0 -1 19848
box -38 -48 406 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 12420 0 -1 19848
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13432 0 -1 19848
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 -1 19848
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 19848
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_137
timestamp 1586364061
transform 1 0 13708 0 -1 19848
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14444 0 -1 19848
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13892 0 -1 19848
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 19848
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16744 0 -1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17388 0 -1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_164
timestamp 1586364061
transform 1 0 16192 0 -1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_168
timestamp 1586364061
transform 1 0 16560 0 -1 19848
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_172
timestamp 1586364061
transform 1 0 16928 0 -1 19848
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_176
timestamp 1586364061
transform 1 0 17296 0 -1 19848
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 -1 19848
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 17940 0 -1 19848
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19044 0 -1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17756 0 -1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_179
timestamp 1586364061
transform 1 0 17572 0 -1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_193
timestamp 1586364061
transform 1 0 18860 0 -1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_197
timestamp 1586364061
transform 1 0 19228 0 -1 19848
box -38 -48 222 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 19596 0 -1 19848
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21068 0 -1 19848
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20884 0 -1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20056 0 -1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 -1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_204
timestamp 1586364061
transform 1 0 19872 0 -1 19848
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_208
timestamp 1586364061
transform 1 0 20240 0 -1 19848
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_214
timestamp 1586364061
transform 1 0 20792 0 -1 19848
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_236
timestamp 1586364061
transform 1 0 22816 0 -1 19848
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 24012 0 -1 19848
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 23552 0 -1 19848
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23828 0 -1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_245
timestamp 1586364061
transform 1 0 23644 0 -1 19848
box -38 -48 222 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 19848
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_268
timestamp 1586364061
transform 1 0 25760 0 -1 19848
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 19848
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 19848
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 20936
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 20936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 20936
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 3956 0 1 19848
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 19848
box -38 -48 406 592
use scs8hd_decap_12  FILLER_33_32
timestamp 1586364061
transform 1 0 4048 0 1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 20936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_39
timestamp 1586364061
transform 1 0 4692 0 -1 20936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_44
timestamp 1586364061
transform 1 0 5152 0 1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 19848
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_51
timestamp 1586364061
transform 1 0 5796 0 -1 20936
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_59
timestamp 1586364061
transform 1 0 6532 0 -1 20936
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 6716 0 -1 20936
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_68
timestamp 1586364061
transform 1 0 7360 0 1 19848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_62
timestamp 1586364061
transform 1 0 6808 0 -1 20936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_74
timestamp 1586364061
transform 1 0 7912 0 -1 20936
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 9568 0 1 19848
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10212 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 1 19848
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_80
timestamp 1586364061
transform 1 0 8464 0 1 19848
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_33_93
timestamp 1586364061
transform 1 0 9660 0 1 19848
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_99
timestamp 1586364061
transform 1 0 10212 0 1 19848
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_86
timestamp 1586364061
transform 1 0 9016 0 -1 20936
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_98
timestamp 1586364061
transform 1 0 10120 0 -1 20936
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_101
timestamp 1586364061
transform 1 0 10396 0 -1 20936
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_107
timestamp 1586364061
transform 1 0 10948 0 1 19848
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_103
timestamp 1586364061
transform 1 0 10580 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 1 19848
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 -1 20936
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_114
timestamp 1586364061
transform 1 0 11592 0 -1 20936
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11224 0 1 19848
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11408 0 1 19848
box -38 -48 1786 592
use scs8hd_buf_1  mux_right_track_26.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12420 0 -1 20936
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 12328 0 -1 20936
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13340 0 1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_131
timestamp 1586364061
transform 1 0 13156 0 1 19848
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 19848
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_126
timestamp 1586364061
transform 1 0 12696 0 -1 20936
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_138
timestamp 1586364061
transform 1 0 13800 0 -1 20936
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_145
timestamp 1586364061
transform 1 0 14444 0 1 19848
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_139
timestamp 1586364061
transform 1 0 13892 0 1 19848
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13984 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14628 0 1 19848
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 14168 0 -1 20936
box -38 -48 866 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 14168 0 1 19848
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 19848
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_149
timestamp 1586364061
transform 1 0 14812 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15640 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14996 0 1 19848
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 15180 0 1 19848
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_151
timestamp 1586364061
transform 1 0 14996 0 -1 20936
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16192 0 1 19848
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 -1 20936
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16008 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16192 0 -1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 19848
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 20936
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_175
timestamp 1586364061
transform 1 0 17204 0 -1 20936
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_187
timestamp 1586364061
transform 1 0 18308 0 1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_183
timestamp 1586364061
transform 1 0 17940 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18124 0 1 19848
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 17940 0 -1 20936
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 -1 20936
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_197
timestamp 1586364061
transform 1 0 19228 0 -1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_193
timestamp 1586364061
transform 1 0 18860 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19044 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18492 0 1 19848
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18676 0 1 19848
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_204
timestamp 1586364061
transform 1 0 19872 0 1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_200
timestamp 1586364061
transform 1 0 19504 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19412 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20056 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19688 0 1 19848
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19596 0 -1 20936
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_217
timestamp 1586364061
transform 1 0 21068 0 -1 20936
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_214
timestamp 1586364061
transform 1 0 20792 0 -1 20936
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_210
timestamp 1586364061
transform 1 0 20424 0 -1 20936
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_218
timestamp 1586364061
transform 1 0 21160 0 1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_212
timestamp 1586364061
transform 1 0 20608 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20884 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20424 0 1 19848
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 20792 0 1 19848
box -38 -48 130 592
use scs8hd_buf_1  mux_right_track_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 1 19848
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_226
timestamp 1586364061
transform 1 0 21896 0 -1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_222
timestamp 1586364061
transform 1 0 21528 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21344 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22080 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21712 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21344 0 -1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_237
timestamp 1586364061
transform 1 0 22908 0 1 19848
box -38 -48 222 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 22632 0 1 19848
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_230
timestamp 1586364061
transform 1 0 22264 0 -1 20936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_222
timestamp 1586364061
transform 1 0 21528 0 1 19848
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_245
timestamp 1586364061
transform 1 0 23644 0 -1 20936
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_242
timestamp 1586364061
transform 1 0 23368 0 -1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_241
timestamp 1586364061
transform 1 0 23276 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23092 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23460 0 1 19848
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 23552 0 -1 20936
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 19848
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 20936
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_254
timestamp 1586364061
transform 1 0 24472 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 19848
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24288 0 -1 20936
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_261
timestamp 1586364061
transform 1 0 25116 0 -1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_266
timestamp 1586364061
transform 1 0 25576 0 1 19848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_258
timestamp 1586364061
transform 1 0 24840 0 1 19848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 25300 0 -1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 19848
box -38 -48 222 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 25208 0 1 19848
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_276
timestamp 1586364061
transform 1 0 26496 0 1 19848
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_274
timestamp 1586364061
transform 1 0 26312 0 1 19848
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_270
timestamp 1586364061
transform 1 0 25944 0 1 19848
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 25760 0 1 19848
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 26404 0 1 19848
box -38 -48 130 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 20936
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 19848
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_265
timestamp 1586364061
transform 1 0 25484 0 -1 20936
box -38 -48 1142 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 20936
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 20936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 20936
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 3956 0 1 20936
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 20936
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 20936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 20936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 20936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_68
timestamp 1586364061
transform 1 0 7360 0 1 20936
box -38 -48 1142 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 9660 0 1 20936
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 9568 0 1 20936
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10120 0 1 20936
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_80
timestamp 1586364061
transform 1 0 8464 0 1 20936
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_35_96
timestamp 1586364061
transform 1 0 9936 0 1 20936
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_26.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10672 0 1 20936
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10488 0 1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_100
timestamp 1586364061
transform 1 0 10304 0 1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13616 0 1 20936
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 20936
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 20936
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_138
timestamp 1586364061
transform 1 0 13800 0 1 20936
box -38 -48 222 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 14168 0 1 20936
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 15180 0 1 20936
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13984 0 1 20936
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_145
timestamp 1586364061
transform 1 0 14444 0 1 20936
box -38 -48 774 592
use scs8hd_decap_12  FILLER_35_154
timestamp 1586364061
transform 1 0 15272 0 1 20936
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17388 0 1 20936
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_166
timestamp 1586364061
transform 1 0 16376 0 1 20936
box -38 -48 774 592
use scs8hd_decap_3  FILLER_35_174
timestamp 1586364061
transform 1 0 17112 0 1 20936
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18308 0 1 20936
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18124 0 1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17756 0 1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_183
timestamp 1586364061
transform 1 0 17940 0 1 20936
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 1 20936
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 20792 0 1 20936
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20608 0 1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_206
timestamp 1586364061
transform 1 0 20056 0 1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_210
timestamp 1586364061
transform 1 0 20424 0 1 20936
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_234
timestamp 1586364061
transform 1 0 22632 0 1 20936
box -38 -48 590 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 23368 0 1 20936
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24380 0 1 20936
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23828 0 1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24196 0 1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_249
timestamp 1586364061
transform 1 0 24012 0 1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_256
timestamp 1586364061
transform 1 0 24656 0 1 20936
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 20936
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 26404 0 1 20936
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24840 0 1 20936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 25208 0 1 20936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_260
timestamp 1586364061
transform 1 0 25024 0 1 20936
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_264
timestamp 1586364061
transform 1 0 25392 0 1 20936
box -38 -48 774 592
use scs8hd_decap_3  FILLER_35_272
timestamp 1586364061
transform 1 0 26128 0 1 20936
box -38 -48 314 592
use scs8hd_fill_1  FILLER_35_276
timestamp 1586364061
transform 1 0 26496 0 1 20936
box -38 -48 130 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22024
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_39
timestamp 1586364061
transform 1 0 4692 0 -1 22024
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_51
timestamp 1586364061
transform 1 0 5796 0 -1 22024
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_59
timestamp 1586364061
transform 1 0 6532 0 -1 22024
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 6716 0 -1 22024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_62
timestamp 1586364061
transform 1 0 6808 0 -1 22024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_74
timestamp 1586364061
transform 1 0 7912 0 -1 22024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_86
timestamp 1586364061
transform 1 0 9016 0 -1 22024
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_98
timestamp 1586364061
transform 1 0 10120 0 -1 22024
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 -1 22024
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10580 0 -1 22024
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22024
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_114
timestamp 1586364061
transform 1 0 11592 0 -1 22024
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13616 0 -1 22024
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 12328 0 -1 22024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_123
timestamp 1586364061
transform 1 0 12420 0 -1 22024
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_135
timestamp 1586364061
transform 1 0 13524 0 -1 22024
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_155
timestamp 1586364061
transform 1 0 15364 0 -1 22024
box -38 -48 774 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 16744 0 -1 22024
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16284 0 -1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17204 0 -1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22024
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_167
timestamp 1586364061
transform 1 0 16468 0 -1 22024
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_173
timestamp 1586364061
transform 1 0 17020 0 -1 22024
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_177
timestamp 1586364061
transform 1 0 17388 0 -1 22024
box -38 -48 590 592
use scs8hd_buf_1  mux_right_track_22.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 -1 22024
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 17940 0 -1 22024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_187
timestamp 1586364061
transform 1 0 18308 0 -1 22024
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19780 0 -1 22024
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19596 0 -1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_199
timestamp 1586364061
transform 1 0 19412 0 -1 22024
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_212
timestamp 1586364061
transform 1 0 20608 0 -1 22024
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21344 0 -1 22024
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22540 0 -1 22024
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_229
timestamp 1586364061
transform 1 0 22172 0 -1 22024
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_235
timestamp 1586364061
transform 1 0 22724 0 -1 22024
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 -1 22024
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 23552 0 -1 22024
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_243
timestamp 1586364061
transform 1 0 23460 0 -1 22024
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_254
timestamp 1586364061
transform 1 0 24472 0 -1 22024
box -38 -48 774 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 25208 0 -1 22024
box -38 -48 406 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22024
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_266
timestamp 1586364061
transform 1 0 25576 0 -1 22024
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22024
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22024
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 1 22024
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22024
box -38 -48 406 592
use scs8hd_decap_12  FILLER_37_32
timestamp 1586364061
transform 1 0 4048 0 1 22024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_44
timestamp 1586364061
transform 1 0 5152 0 1 22024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_56
timestamp 1586364061
transform 1 0 6256 0 1 22024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_68
timestamp 1586364061
transform 1 0 7360 0 1 22024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 1 22024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22024
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_93
timestamp 1586364061
transform 1 0 9660 0 1 22024
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_26.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10764 0 1 22024
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10580 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_101
timestamp 1586364061
transform 1 0 10396 0 1 22024
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 1 22024
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13432 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13064 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12696 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_124
timestamp 1586364061
transform 1 0 12512 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_128
timestamp 1586364061
transform 1 0 12880 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22024
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 15180 0 1 22024
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_145
timestamp 1586364061
transform 1 0 14444 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_149
timestamp 1586364061
transform 1 0 14812 0 1 22024
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_154
timestamp 1586364061
transform 1 0 15272 0 1 22024
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_158
timestamp 1586364061
transform 1 0 15640 0 1 22024
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_22.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16284 0 1 22024
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16100 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_161
timestamp 1586364061
transform 1 0 15916 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18584 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18952 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_192
timestamp 1586364061
transform 1 0 18768 0 1 22024
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22024
box -38 -48 406 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 19780 0 1 22024
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_20.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 1 22024
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 20792 0 1 22024
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19596 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20240 0 1 22024
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_200
timestamp 1586364061
transform 1 0 19504 0 1 22024
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_206
timestamp 1586364061
transform 1 0 20056 0 1 22024
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_210
timestamp 1586364061
transform 1 0 20424 0 1 22024
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_218
timestamp 1586364061
transform 1 0 21160 0 1 22024
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21896 0 1 22024
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21712 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21344 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_222
timestamp 1586364061
transform 1 0 21528 0 1 22024
box -38 -48 222 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 24564 0 1 22024
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23828 0 1 22024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24196 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_249
timestamp 1586364061
transform 1 0 24012 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22024
box -38 -48 222 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22024
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 26404 0 1 22024
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 25116 0 1 22024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_259
timestamp 1586364061
transform 1 0 24932 0 1 22024
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_263
timestamp 1586364061
transform 1 0 25300 0 1 22024
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_37_276
timestamp 1586364061
transform 1 0 26496 0 1 22024
box -38 -48 130 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23112
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_39
timestamp 1586364061
transform 1 0 4692 0 -1 23112
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_51
timestamp 1586364061
transform 1 0 5796 0 -1 23112
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_59
timestamp 1586364061
transform 1 0 6532 0 -1 23112
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6716 0 -1 23112
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_62
timestamp 1586364061
transform 1 0 6808 0 -1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_74
timestamp 1586364061
transform 1 0 7912 0 -1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_86
timestamp 1586364061
transform 1 0 9016 0 -1 23112
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_38_98
timestamp 1586364061
transform 1 0 10120 0 -1 23112
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10764 0 -1 23112
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_104
timestamp 1586364061
transform 1 0 10672 0 -1 23112
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_107
timestamp 1586364061
transform 1 0 10948 0 -1 23112
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_38_119
timestamp 1586364061
transform 1 0 12052 0 -1 23112
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13800 0 -1 23112
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 12328 0 -1 23112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13616 0 -1 23112
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_123
timestamp 1586364061
transform 1 0 12420 0 -1 23112
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_135
timestamp 1586364061
transform 1 0 13524 0 -1 23112
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_147
timestamp 1586364061
transform 1 0 14628 0 -1 23112
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 -1 23112
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16192 0 -1 23112
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_159
timestamp 1586364061
transform 1 0 15732 0 -1 23112
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23112
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_175
timestamp 1586364061
transform 1 0 17204 0 -1 23112
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 -1 23112
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 17940 0 -1 23112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19228 0 -1 23112
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23112
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_20.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19596 0 -1 23112
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_38_199
timestamp 1586364061
transform 1 0 19412 0 -1 23112
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_18.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22540 0 -1 23112
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21896 0 -1 23112
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_220
timestamp 1586364061
transform 1 0 21344 0 -1 23112
box -38 -48 590 592
use scs8hd_decap_4  FILLER_38_228
timestamp 1586364061
transform 1 0 22080 0 -1 23112
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_232
timestamp 1586364061
transform 1 0 22448 0 -1 23112
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_236
timestamp 1586364061
transform 1 0 22816 0 -1 23112
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_track_18.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 -1 23112
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 23552 0 -1 23112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 -1 23112
box -38 -48 222 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23112
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_264
timestamp 1586364061
transform 1 0 25392 0 -1 23112
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23112
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23112
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24200
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24200
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 3956 0 1 23112
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23112
box -38 -48 406 592
use scs8hd_decap_12  FILLER_39_32
timestamp 1586364061
transform 1 0 4048 0 1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_39
timestamp 1586364061
transform 1 0 4692 0 -1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_44
timestamp 1586364061
transform 1 0 5152 0 1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_56
timestamp 1586364061
transform 1 0 6256 0 1 23112
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_51
timestamp 1586364061
transform 1 0 5796 0 -1 24200
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_59
timestamp 1586364061
transform 1 0 6532 0 -1 24200
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 6716 0 -1 24200
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_68
timestamp 1586364061
transform 1 0 7360 0 1 23112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_62
timestamp 1586364061
transform 1 0 6808 0 -1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_74
timestamp 1586364061
transform 1 0 7912 0 -1 24200
box -38 -48 1142 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 9660 0 1 23112
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 9568 0 1 23112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 10212 0 1 23112
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_80
timestamp 1586364061
transform 1 0 8464 0 1 23112
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_97
timestamp 1586364061
transform 1 0 10028 0 1 23112
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_86
timestamp 1586364061
transform 1 0 9016 0 -1 24200
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_98
timestamp 1586364061
transform 1 0 10120 0 -1 24200
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_106
timestamp 1586364061
transform 1 0 10856 0 -1 24200
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23112
box -38 -48 406 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 10764 0 1 23112
box -38 -48 406 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 10948 0 -1 24200
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_111
timestamp 1586364061
transform 1 0 11316 0 -1 24200
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_113
timestamp 1586364061
transform 1 0 11500 0 1 23112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_109
timestamp 1586364061
transform 1 0 11132 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 11684 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 11316 0 1 23112
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_119
timestamp 1586364061
transform 1 0 12052 0 -1 24200
box -38 -48 314 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 11868 0 1 23112
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_125
timestamp 1586364061
transform 1 0 12604 0 1 23112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12788 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 12420 0 1 23112
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 12328 0 -1 24200
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_135
timestamp 1586364061
transform 1 0 13524 0 -1 24200
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_137
timestamp 1586364061
transform 1 0 13708 0 1 23112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_133
timestamp 1586364061
transform 1 0 13340 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 13524 0 1 23112
box -38 -48 222 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 12972 0 1 23112
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_123
timestamp 1586364061
transform 1 0 12420 0 -1 24200
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13708 0 -1 24200
box -38 -48 1786 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 15272 0 1 23112
box -38 -48 406 592
use scs8hd_buf_2  _75_
timestamp 1586364061
transform 1 0 14076 0 1 23112
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 15180 0 1 23112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13892 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__75__A
timestamp 1586364061
transform 1 0 14628 0 1 23112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_145
timestamp 1586364061
transform 1 0 14444 0 1 23112
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_149
timestamp 1586364061
transform 1 0 14812 0 1 23112
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23112
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_156
timestamp 1586364061
transform 1 0 15456 0 -1 24200
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_164
timestamp 1586364061
transform 1 0 16192 0 -1 24200
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_162
timestamp 1586364061
transform 1 0 16008 0 1 23112
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 15824 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16468 0 -1 24200
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16284 0 1 23112
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_177
timestamp 1586364061
transform 1 0 17388 0 -1 24200
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_173
timestamp 1586364061
transform 1 0 17020 0 -1 24200
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 17204 0 -1 24200
box -38 -48 222 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 16652 0 -1 24200
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_22.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16468 0 1 23112
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_39_186
timestamp 1586364061
transform 1 0 18216 0 1 23112
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 17940 0 -1 24200
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_196
timestamp 1586364061
transform 1 0 19136 0 -1 24200
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23112
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_190
timestamp 1586364061
transform 1 0 18584 0 1 23112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19228 0 -1 24200
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18676 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 1 23112
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 1 23112
box -38 -48 866 592
use scs8hd_decap_12  FILLER_40_184
timestamp 1586364061
transform 1 0 18032 0 -1 24200
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_20.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19596 0 -1 24200
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 20792 0 1 23112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20240 0 1 23112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_206
timestamp 1586364061
transform 1 0 20056 0 1 23112
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_210
timestamp 1586364061
transform 1 0 20424 0 1 23112
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_215
timestamp 1586364061
transform 1 0 20884 0 1 23112
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_199
timestamp 1586364061
transform 1 0 19412 0 -1 24200
box -38 -48 222 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 22724 0 1 23112
box -38 -48 314 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 21252 0 1 23112
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 21804 0 1 23112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23112
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23112
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_238
timestamp 1586364061
transform 1 0 23000 0 1 23112
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_220
timestamp 1586364061
transform 1 0 21344 0 -1 24200
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_232
timestamp 1586364061
transform 1 0 22448 0 -1 24200
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_245
timestamp 1586364061
transform 1 0 23644 0 -1 24200
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_240
timestamp 1586364061
transform 1 0 23184 0 -1 24200
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_242
timestamp 1586364061
transform 1 0 23368 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23828 0 -1 24200
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23184 0 1 23112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 -1 24200
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23552 0 1 23112
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 23552 0 -1 24200
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_249
timestamp 1586364061
transform 1 0 24012 0 -1 24200
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24104 0 -1 24200
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_18.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23736 0 1 23112
box -38 -48 1786 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23112
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24200
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 26404 0 1 23112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 25668 0 1 23112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_265
timestamp 1586364061
transform 1 0 25484 0 1 23112
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23112
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_276
timestamp 1586364061
transform 1 0 26496 0 1 23112
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_259
timestamp 1586364061
transform 1 0 24932 0 -1 24200
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24200
box -38 -48 590 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24200
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24200
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 3956 0 1 24200
box -38 -48 130 592
use scs8hd_decap_4  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24200
box -38 -48 406 592
use scs8hd_decap_12  FILLER_41_32
timestamp 1586364061
transform 1 0 4048 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_44
timestamp 1586364061
transform 1 0 5152 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_56
timestamp 1586364061
transform 1 0 6256 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_68
timestamp 1586364061
transform 1 0 7360 0 1 24200
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 9568 0 1 24200
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_80
timestamp 1586364061
transform 1 0 8464 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_93
timestamp 1586364061
transform 1 0 9660 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_105
timestamp 1586364061
transform 1 0 10764 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_117
timestamp 1586364061
transform 1 0 11868 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_129
timestamp 1586364061
transform 1 0 12972 0 1 24200
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 15180 0 1 24200
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_141
timestamp 1586364061
transform 1 0 14076 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_154
timestamp 1586364061
transform 1 0 15272 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_166
timestamp 1586364061
transform 1 0 16376 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_178
timestamp 1586364061
transform 1 0 17480 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_190
timestamp 1586364061
transform 1 0 18584 0 1 24200
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 20792 0 1 24200
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_202
timestamp 1586364061
transform 1 0 19688 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_215
timestamp 1586364061
transform 1 0 20884 0 1 24200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_227
timestamp 1586364061
transform 1 0 21988 0 1 24200
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23368 0 1 24200
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 1 24200
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_239
timestamp 1586364061
transform 1 0 23092 0 1 24200
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_251
timestamp 1586364061
transform 1 0 24196 0 1 24200
box -38 -48 774 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 24932 0 1 24200
box -38 -48 406 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24200
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 26404 0 1 24200
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 25484 0 1 24200
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_263
timestamp 1586364061
transform 1 0 25300 0 1 24200
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_267
timestamp 1586364061
transform 1 0 25668 0 1 24200
box -38 -48 774 592
use scs8hd_fill_1  FILLER_41_276
timestamp 1586364061
transform 1 0 26496 0 1 24200
box -38 -48 130 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25288
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 3956 0 -1 25288
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25288
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25288
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 6808 0 -1 25288
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 9660 0 -1 25288
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25288
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25288
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 12512 0 -1 25288
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 15364 0 -1 25288
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25288
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 18216 0 -1 25288
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25288
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 21068 0 -1 25288
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25288
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 23920 0 -1 25288
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23368 0 -1 25288
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_244
timestamp 1586364061
transform 1 0 23552 0 -1 25288
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25288
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25288
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25288
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 13600 480 13720 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 22984 480 23104 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 27520 544 28000 664 6 chanx_right_in[0]
port 2 nsew default input
rlabel metal3 s 27520 6256 28000 6376 6 chanx_right_in[10]
port 3 nsew default input
rlabel metal3 s 27520 6800 28000 6920 6 chanx_right_in[11]
port 4 nsew default input
rlabel metal3 s 27520 7344 28000 7464 6 chanx_right_in[12]
port 5 nsew default input
rlabel metal3 s 27520 7888 28000 8008 6 chanx_right_in[13]
port 6 nsew default input
rlabel metal3 s 27520 8568 28000 8688 6 chanx_right_in[14]
port 7 nsew default input
rlabel metal3 s 27520 9112 28000 9232 6 chanx_right_in[15]
port 8 nsew default input
rlabel metal3 s 27520 9656 28000 9776 6 chanx_right_in[16]
port 9 nsew default input
rlabel metal3 s 27520 10200 28000 10320 6 chanx_right_in[17]
port 10 nsew default input
rlabel metal3 s 27520 10744 28000 10864 6 chanx_right_in[18]
port 11 nsew default input
rlabel metal3 s 27520 11424 28000 11544 6 chanx_right_in[19]
port 12 nsew default input
rlabel metal3 s 27520 1088 28000 1208 6 chanx_right_in[1]
port 13 nsew default input
rlabel metal3 s 27520 1632 28000 1752 6 chanx_right_in[2]
port 14 nsew default input
rlabel metal3 s 27520 2176 28000 2296 6 chanx_right_in[3]
port 15 nsew default input
rlabel metal3 s 27520 2856 28000 2976 6 chanx_right_in[4]
port 16 nsew default input
rlabel metal3 s 27520 3400 28000 3520 6 chanx_right_in[5]
port 17 nsew default input
rlabel metal3 s 27520 3944 28000 4064 6 chanx_right_in[6]
port 18 nsew default input
rlabel metal3 s 27520 4488 28000 4608 6 chanx_right_in[7]
port 19 nsew default input
rlabel metal3 s 27520 5032 28000 5152 6 chanx_right_in[8]
port 20 nsew default input
rlabel metal3 s 27520 5712 28000 5832 6 chanx_right_in[9]
port 21 nsew default input
rlabel metal3 s 27520 11968 28000 12088 6 chanx_right_out[0]
port 22 nsew default tristate
rlabel metal3 s 27520 17680 28000 17800 6 chanx_right_out[10]
port 23 nsew default tristate
rlabel metal3 s 27520 18224 28000 18344 6 chanx_right_out[11]
port 24 nsew default tristate
rlabel metal3 s 27520 18768 28000 18888 6 chanx_right_out[12]
port 25 nsew default tristate
rlabel metal3 s 27520 19312 28000 19432 6 chanx_right_out[13]
port 26 nsew default tristate
rlabel metal3 s 27520 19992 28000 20112 6 chanx_right_out[14]
port 27 nsew default tristate
rlabel metal3 s 27520 20536 28000 20656 6 chanx_right_out[15]
port 28 nsew default tristate
rlabel metal3 s 27520 21080 28000 21200 6 chanx_right_out[16]
port 29 nsew default tristate
rlabel metal3 s 27520 21624 28000 21744 6 chanx_right_out[17]
port 30 nsew default tristate
rlabel metal3 s 27520 22168 28000 22288 6 chanx_right_out[18]
port 31 nsew default tristate
rlabel metal3 s 27520 22848 28000 22968 6 chanx_right_out[19]
port 32 nsew default tristate
rlabel metal3 s 27520 12512 28000 12632 6 chanx_right_out[1]
port 33 nsew default tristate
rlabel metal3 s 27520 13056 28000 13176 6 chanx_right_out[2]
port 34 nsew default tristate
rlabel metal3 s 27520 13600 28000 13720 6 chanx_right_out[3]
port 35 nsew default tristate
rlabel metal3 s 27520 14280 28000 14400 6 chanx_right_out[4]
port 36 nsew default tristate
rlabel metal3 s 27520 14824 28000 14944 6 chanx_right_out[5]
port 37 nsew default tristate
rlabel metal3 s 27520 15368 28000 15488 6 chanx_right_out[6]
port 38 nsew default tristate
rlabel metal3 s 27520 15912 28000 16032 6 chanx_right_out[7]
port 39 nsew default tristate
rlabel metal3 s 27520 16456 28000 16576 6 chanx_right_out[8]
port 40 nsew default tristate
rlabel metal3 s 27520 17136 28000 17256 6 chanx_right_out[9]
port 41 nsew default tristate
rlabel metal2 s 938 27240 994 27720 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 7746 27240 7802 27720 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 8390 27240 8446 27720 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 9126 27240 9182 27720 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 9770 27240 9826 27720 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 10506 27240 10562 27720 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 11150 27240 11206 27720 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 11886 27240 11942 27720 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 12530 27240 12586 27720 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 13174 27240 13230 27720 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 13910 27240 13966 27720 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 1582 27240 1638 27720 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 2318 27240 2374 27720 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 2962 27240 3018 27720 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 3698 27240 3754 27720 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 4342 27240 4398 27720 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 4986 27240 5042 27720 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 5722 27240 5778 27720 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 6366 27240 6422 27720 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 7102 27240 7158 27720 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 14554 27240 14610 27720 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 21362 27240 21418 27720 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 22098 27240 22154 27720 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 22742 27240 22798 27720 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 23478 27240 23534 27720 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 24122 27240 24178 27720 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24766 27240 24822 27720 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 25502 27240 25558 27720 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 26146 27240 26202 27720 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 26882 27240 26938 27720 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 27526 27240 27582 27720 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 15290 27240 15346 27720 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 15934 27240 15990 27720 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 16578 27240 16634 27720 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 17314 27240 17370 27720 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 17958 27240 18014 27720 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 18694 27240 18750 27720 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 19338 27240 19394 27720 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 20074 27240 20130 27720 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 20718 27240 20774 27720 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 4352 480 4472 6 prog_clk
port 82 nsew default input
rlabel metal3 s 27520 0 28000 120 6 right_bottom_grid_pin_1_
port 83 nsew default input
rlabel metal3 s 27520 23392 28000 23512 6 right_top_grid_pin_42_
port 84 nsew default input
rlabel metal3 s 27520 23936 28000 24056 6 right_top_grid_pin_43_
port 85 nsew default input
rlabel metal3 s 27520 24480 28000 24600 6 right_top_grid_pin_44_
port 86 nsew default input
rlabel metal3 s 27520 25024 28000 25144 6 right_top_grid_pin_45_
port 87 nsew default input
rlabel metal3 s 27520 25704 28000 25824 6 right_top_grid_pin_46_
port 88 nsew default input
rlabel metal3 s 27520 26248 28000 26368 6 right_top_grid_pin_47_
port 89 nsew default input
rlabel metal3 s 27520 26792 28000 26912 6 right_top_grid_pin_48_
port 90 nsew default input
rlabel metal3 s 27520 27336 28000 27456 6 right_top_grid_pin_49_
port 91 nsew default input
rlabel metal2 s 294 27240 350 27720 6 top_left_grid_pin_1_
port 92 nsew default input
rlabel metal4 s 5611 1848 5931 25336 6 vpwr
port 93 nsew default input
rlabel metal4 s 10277 1848 10597 25336 6 vgnd
port 94 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 27720
<< end >>
