magic
tech sky130A
magscale 1 2
timestamp 1608762278
<< checkpaint >>
rect -1260 -1260 24060 24060
<< locali >>
rect 16405 19703 16439 19873
rect 10149 19159 10183 19261
rect 12449 19159 12483 19329
rect 19349 19159 19383 19261
rect 8125 18751 8159 18921
rect 6929 17731 6963 17833
rect 3893 17595 3927 17697
rect 4169 16575 4203 16745
rect 11529 16643 11563 16745
rect 12173 15487 12207 15589
rect 5549 15351 5583 15453
rect 13737 15419 13771 15589
rect 7297 14331 7331 14569
rect 17877 13787 17911 13957
rect 15025 13311 15059 13413
rect 17785 12835 17819 12937
rect 12173 12631 12207 12733
rect 9505 12223 9539 12393
rect 12725 12087 12759 12257
rect 18981 11747 19015 11849
rect 3893 10999 3927 11237
rect 15393 10999 15427 11101
rect 6837 10455 6871 10625
rect 5457 10217 5549 10251
rect 5457 9979 5491 10217
rect 16129 8891 16163 8993
rect 5457 7871 5491 8041
<< viali >>
rect 2053 20009 2087 20043
rect 9045 20009 9079 20043
rect 9781 20009 9815 20043
rect 10241 20009 10275 20043
rect 14473 20009 14507 20043
rect 15025 20009 15059 20043
rect 15669 20009 15703 20043
rect 16773 20009 16807 20043
rect 18521 20009 18555 20043
rect 19073 20009 19107 20043
rect 19625 20009 19659 20043
rect 7481 19941 7515 19975
rect 1869 19873 1903 19907
rect 2421 19873 2455 19907
rect 8125 19873 8159 19907
rect 10149 19873 10183 19907
rect 11989 19873 12023 19907
rect 13001 19873 13035 19907
rect 13737 19873 13771 19907
rect 14289 19873 14323 19907
rect 14841 19873 14875 19907
rect 15485 19873 15519 19907
rect 16037 19873 16071 19907
rect 16405 19873 16439 19907
rect 16589 19873 16623 19907
rect 17325 19873 17359 19907
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 19441 19873 19475 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 7573 19805 7607 19839
rect 7665 19805 7699 19839
rect 9137 19805 9171 19839
rect 9321 19805 9355 19839
rect 10333 19805 10367 19839
rect 13093 19805 13127 19839
rect 13185 19805 13219 19839
rect 8309 19737 8343 19771
rect 16221 19737 16255 19771
rect 17509 19737 17543 19771
rect 20177 19737 20211 19771
rect 2605 19669 2639 19703
rect 7113 19669 7147 19703
rect 8677 19669 8711 19703
rect 12173 19669 12207 19703
rect 12633 19669 12667 19703
rect 13921 19669 13955 19703
rect 16405 19669 16439 19703
rect 20729 19669 20763 19703
rect 3525 19465 3559 19499
rect 5733 19465 5767 19499
rect 12541 19465 12575 19499
rect 19625 19465 19659 19499
rect 7297 19329 7331 19363
rect 12449 19329 12483 19363
rect 13185 19329 13219 19363
rect 17509 19329 17543 19363
rect 18889 19329 18923 19363
rect 1869 19261 1903 19295
rect 2421 19261 2455 19295
rect 3341 19261 3375 19295
rect 3985 19261 4019 19295
rect 5549 19261 5583 19295
rect 7021 19261 7055 19295
rect 7757 19261 7791 19295
rect 9597 19261 9631 19295
rect 10149 19261 10183 19295
rect 10333 19261 10367 19295
rect 10589 19261 10623 19295
rect 4721 19193 4755 19227
rect 8002 19193 8036 19227
rect 9873 19193 9907 19227
rect 14013 19261 14047 19295
rect 14749 19261 14783 19295
rect 15301 19261 15335 19295
rect 16037 19261 16071 19295
rect 18153 19261 18187 19295
rect 18705 19261 18739 19295
rect 19349 19261 19383 19295
rect 19441 19261 19475 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 13001 19193 13035 19227
rect 14289 19193 14323 19227
rect 15577 19193 15611 19227
rect 17325 19193 17359 19227
rect 2053 19125 2087 19159
rect 2605 19125 2639 19159
rect 9137 19125 9171 19159
rect 10149 19125 10183 19159
rect 11713 19125 11747 19159
rect 12449 19125 12483 19159
rect 12909 19125 12943 19159
rect 13553 19125 13587 19159
rect 14933 19125 14967 19159
rect 16221 19125 16255 19159
rect 16865 19125 16899 19159
rect 17233 19125 17267 19159
rect 18337 19125 18371 19159
rect 19349 19125 19383 19159
rect 20177 19125 20211 19159
rect 20729 19125 20763 19159
rect 2053 18921 2087 18955
rect 2605 18921 2639 18955
rect 3157 18921 3191 18955
rect 8125 18921 8159 18955
rect 11069 18921 11103 18955
rect 13093 18921 13127 18955
rect 15761 18921 15795 18955
rect 17785 18921 17819 18955
rect 18797 18921 18831 18955
rect 20269 18921 20303 18955
rect 6828 18853 6862 18887
rect 1869 18785 1903 18819
rect 2421 18785 2455 18819
rect 2973 18785 3007 18819
rect 4077 18785 4111 18819
rect 9956 18853 9990 18887
rect 11980 18853 12014 18887
rect 13614 18853 13648 18887
rect 18337 18853 18371 18887
rect 19257 18853 19291 18887
rect 8585 18785 8619 18819
rect 9689 18785 9723 18819
rect 15669 18785 15703 18819
rect 16405 18785 16439 18819
rect 16672 18785 16706 18819
rect 18061 18785 18095 18819
rect 19165 18785 19199 18819
rect 20177 18785 20211 18819
rect 6561 18717 6595 18751
rect 8125 18717 8159 18751
rect 8677 18717 8711 18751
rect 8769 18717 8803 18751
rect 11713 18717 11747 18751
rect 13369 18717 13403 18751
rect 15853 18717 15887 18751
rect 19349 18717 19383 18751
rect 20361 18717 20395 18751
rect 20913 18717 20947 18751
rect 4261 18649 4295 18683
rect 14749 18649 14783 18683
rect 19809 18649 19843 18683
rect 7941 18581 7975 18615
rect 8217 18581 8251 18615
rect 15301 18581 15335 18615
rect 1961 18377 1995 18411
rect 2513 18377 2547 18411
rect 9505 18377 9539 18411
rect 12541 18377 12575 18411
rect 13737 18377 13771 18411
rect 17141 18377 17175 18411
rect 17601 18377 17635 18411
rect 19717 18377 19751 18411
rect 3065 18309 3099 18343
rect 11069 18309 11103 18343
rect 6101 18241 6135 18275
rect 6837 18241 6871 18275
rect 8493 18241 8527 18275
rect 10057 18241 10091 18275
rect 10517 18241 10551 18275
rect 11621 18241 11655 18275
rect 13185 18241 13219 18275
rect 14105 18241 14139 18275
rect 20269 18241 20303 18275
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 2881 18173 2915 18207
rect 3433 18173 3467 18207
rect 5917 18173 5951 18207
rect 7104 18173 7138 18207
rect 13553 18173 13587 18207
rect 14372 18173 14406 18207
rect 15761 18173 15795 18207
rect 17417 18173 17451 18207
rect 18061 18173 18095 18207
rect 20177 18173 20211 18207
rect 20729 18173 20763 18207
rect 11529 18105 11563 18139
rect 12909 18105 12943 18139
rect 16006 18105 16040 18139
rect 18306 18105 18340 18139
rect 20085 18105 20119 18139
rect 3617 18037 3651 18071
rect 8217 18037 8251 18071
rect 9873 18037 9907 18071
rect 9965 18037 9999 18071
rect 11437 18037 11471 18071
rect 13001 18037 13035 18071
rect 15485 18037 15519 18071
rect 19441 18037 19475 18071
rect 20913 18037 20947 18071
rect 6929 17833 6963 17867
rect 7113 17833 7147 17867
rect 7481 17833 7515 17867
rect 7573 17833 7607 17867
rect 8585 17833 8619 17867
rect 9873 17833 9907 17867
rect 12081 17833 12115 17867
rect 12541 17833 12575 17867
rect 15301 17833 15335 17867
rect 15669 17833 15703 17867
rect 16497 17833 16531 17867
rect 16865 17833 16899 17867
rect 17509 17833 17543 17867
rect 17877 17833 17911 17867
rect 20913 17833 20947 17867
rect 2513 17765 2547 17799
rect 18880 17765 18914 17799
rect 1685 17697 1719 17731
rect 2237 17697 2271 17731
rect 3893 17697 3927 17731
rect 5089 17697 5123 17731
rect 5365 17697 5399 17731
rect 5825 17697 5859 17731
rect 6929 17697 6963 17731
rect 8493 17697 8527 17731
rect 9689 17697 9723 17731
rect 10425 17697 10459 17731
rect 10692 17697 10726 17731
rect 12449 17697 12483 17731
rect 13093 17697 13127 17731
rect 14565 17697 14599 17731
rect 15761 17697 15795 17731
rect 17969 17697 18003 17731
rect 20269 17697 20303 17731
rect 7757 17629 7791 17663
rect 8769 17629 8803 17663
rect 12633 17629 12667 17663
rect 13277 17629 13311 17663
rect 14657 17629 14691 17663
rect 14841 17629 14875 17663
rect 15853 17629 15887 17663
rect 16957 17629 16991 17663
rect 17049 17629 17083 17663
rect 18061 17629 18095 17663
rect 18613 17629 18647 17663
rect 1869 17561 1903 17595
rect 3893 17561 3927 17595
rect 6009 17561 6043 17595
rect 11805 17561 11839 17595
rect 14197 17561 14231 17595
rect 8125 17493 8159 17527
rect 19993 17493 20027 17527
rect 20453 17493 20487 17527
rect 2513 17289 2547 17323
rect 3065 17289 3099 17323
rect 3617 17289 3651 17323
rect 5457 17289 5491 17323
rect 10885 17289 10919 17323
rect 14381 17221 14415 17255
rect 4997 17153 5031 17187
rect 6009 17153 6043 17187
rect 7481 17153 7515 17187
rect 8309 17153 8343 17187
rect 8493 17153 8527 17187
rect 9137 17153 9171 17187
rect 11529 17153 11563 17187
rect 11897 17153 11931 17187
rect 12633 17153 12667 17187
rect 13553 17153 13587 17187
rect 13737 17153 13771 17187
rect 15025 17153 15059 17187
rect 16589 17153 16623 17187
rect 18613 17153 18647 17187
rect 19625 17153 19659 17187
rect 1777 17085 1811 17119
rect 2329 17085 2363 17119
rect 2881 17085 2915 17119
rect 3433 17085 3467 17119
rect 7205 17085 7239 17119
rect 8217 17085 8251 17119
rect 8861 17085 8895 17119
rect 13461 17085 13495 17119
rect 15393 17085 15427 17119
rect 16313 17085 16347 17119
rect 17141 17085 17175 17119
rect 20545 17085 20579 17119
rect 5917 17017 5951 17051
rect 11345 17017 11379 17051
rect 14841 17017 14875 17051
rect 15669 17017 15703 17051
rect 17417 17017 17451 17051
rect 18429 17017 18463 17051
rect 1961 16949 1995 16983
rect 4445 16949 4479 16983
rect 4813 16949 4847 16983
rect 4905 16949 4939 16983
rect 5825 16949 5859 16983
rect 6837 16949 6871 16983
rect 7297 16949 7331 16983
rect 7849 16949 7883 16983
rect 11253 16949 11287 16983
rect 13093 16949 13127 16983
rect 14749 16949 14783 16983
rect 18061 16949 18095 16983
rect 18521 16949 18555 16983
rect 19073 16949 19107 16983
rect 19441 16949 19475 16983
rect 19533 16949 19567 16983
rect 20085 16949 20119 16983
rect 20729 16949 20763 16983
rect 2605 16745 2639 16779
rect 4169 16745 4203 16779
rect 5641 16745 5675 16779
rect 10701 16745 10735 16779
rect 11529 16745 11563 16779
rect 13001 16745 13035 16779
rect 14473 16745 14507 16779
rect 15301 16745 15335 16779
rect 15761 16745 15795 16779
rect 17877 16745 17911 16779
rect 18613 16745 18647 16779
rect 20361 16745 20395 16779
rect 1777 16609 1811 16643
rect 2973 16609 3007 16643
rect 3065 16609 3099 16643
rect 4528 16677 4562 16711
rect 6162 16677 6196 16711
rect 7818 16677 7852 16711
rect 10149 16677 10183 16711
rect 13369 16677 13403 16711
rect 13461 16677 13495 16711
rect 16764 16677 16798 16711
rect 7573 16609 7607 16643
rect 10057 16609 10091 16643
rect 11069 16609 11103 16643
rect 11529 16609 11563 16643
rect 12081 16609 12115 16643
rect 14381 16609 14415 16643
rect 15669 16609 15703 16643
rect 16497 16609 16531 16643
rect 18429 16609 18463 16643
rect 19248 16609 19282 16643
rect 3249 16541 3283 16575
rect 4169 16541 4203 16575
rect 4261 16541 4295 16575
rect 5917 16541 5951 16575
rect 10241 16541 10275 16575
rect 11161 16541 11195 16575
rect 11345 16541 11379 16575
rect 12173 16541 12207 16575
rect 12265 16541 12299 16575
rect 13645 16541 13679 16575
rect 14565 16541 14599 16575
rect 15853 16541 15887 16575
rect 18981 16541 19015 16575
rect 1961 16473 1995 16507
rect 8953 16473 8987 16507
rect 9689 16473 9723 16507
rect 11713 16473 11747 16507
rect 14013 16473 14047 16507
rect 7297 16405 7331 16439
rect 4997 16201 5031 16235
rect 6009 16201 6043 16235
rect 8217 16201 8251 16235
rect 10517 16201 10551 16235
rect 16037 16201 16071 16235
rect 16497 16201 16531 16235
rect 16865 16201 16899 16235
rect 20269 16201 20303 16235
rect 4445 16133 4479 16167
rect 10149 16133 10183 16167
rect 12633 16133 12667 16167
rect 5549 16065 5583 16099
rect 8769 16065 8803 16099
rect 11161 16065 11195 16099
rect 11897 16065 11931 16099
rect 13001 16065 13035 16099
rect 17509 16065 17543 16099
rect 1777 15997 1811 16031
rect 2329 15997 2363 16031
rect 3065 15997 3099 16031
rect 5457 15997 5491 16031
rect 6193 15997 6227 16031
rect 6837 15997 6871 16031
rect 8677 15997 8711 16031
rect 9036 15997 9070 16031
rect 10977 15997 11011 16031
rect 11621 15997 11655 16031
rect 12817 15997 12851 16031
rect 13268 15997 13302 16031
rect 14657 15997 14691 16031
rect 16313 15997 16347 16031
rect 18337 15997 18371 16031
rect 18889 15997 18923 16031
rect 20545 15997 20579 16031
rect 3332 15929 3366 15963
rect 7104 15929 7138 15963
rect 10885 15929 10919 15963
rect 14902 15929 14936 15963
rect 19156 15929 19190 15963
rect 1961 15861 1995 15895
rect 2513 15861 2547 15895
rect 5365 15861 5399 15895
rect 8493 15861 8527 15895
rect 14381 15861 14415 15895
rect 17233 15861 17267 15895
rect 17325 15861 17359 15895
rect 18521 15861 18555 15895
rect 20729 15861 20763 15895
rect 3249 15657 3283 15691
rect 4629 15657 4663 15691
rect 5089 15657 5123 15691
rect 5641 15657 5675 15691
rect 7389 15657 7423 15691
rect 8033 15657 8067 15691
rect 8493 15657 8527 15691
rect 11989 15657 12023 15691
rect 13921 15657 13955 15691
rect 14381 15657 14415 15691
rect 18061 15657 18095 15691
rect 19073 15657 19107 15691
rect 3157 15589 3191 15623
rect 6009 15589 6043 15623
rect 12173 15589 12207 15623
rect 12532 15589 12566 15623
rect 13737 15589 13771 15623
rect 15660 15589 15694 15623
rect 17509 15589 17543 15623
rect 18429 15589 18463 15623
rect 20361 15589 20395 15623
rect 1777 15521 1811 15555
rect 4997 15521 5031 15555
rect 7481 15521 7515 15555
rect 8401 15521 8435 15555
rect 9045 15521 9079 15555
rect 10609 15521 10643 15555
rect 10876 15521 10910 15555
rect 3433 15453 3467 15487
rect 5273 15453 5307 15487
rect 5549 15453 5583 15487
rect 6101 15453 6135 15487
rect 6193 15453 6227 15487
rect 7573 15453 7607 15487
rect 8677 15453 8711 15487
rect 12173 15453 12207 15487
rect 12265 15453 12299 15487
rect 2789 15385 2823 15419
rect 14289 15521 14323 15555
rect 15393 15521 15427 15555
rect 17417 15521 17451 15555
rect 18521 15521 18555 15555
rect 19441 15521 19475 15555
rect 20085 15521 20119 15555
rect 14473 15453 14507 15487
rect 17601 15453 17635 15487
rect 18705 15453 18739 15487
rect 19533 15453 19567 15487
rect 19625 15453 19659 15487
rect 7021 15385 7055 15419
rect 13737 15385 13771 15419
rect 16773 15385 16807 15419
rect 1961 15317 1995 15351
rect 5549 15317 5583 15351
rect 13645 15317 13679 15351
rect 17049 15317 17083 15351
rect 4169 15113 4203 15147
rect 7389 15113 7423 15147
rect 8401 15113 8435 15147
rect 11069 15113 11103 15147
rect 13277 15113 13311 15147
rect 19441 15113 19475 15147
rect 3709 15045 3743 15079
rect 11345 15045 11379 15079
rect 14105 15045 14139 15079
rect 17693 15045 17727 15079
rect 1869 14977 1903 15011
rect 4813 14977 4847 15011
rect 5181 14977 5215 15011
rect 6193 14977 6227 15011
rect 6377 14977 6411 15011
rect 8033 14977 8067 15011
rect 8953 14977 8987 15011
rect 11989 14977 12023 15011
rect 13001 14977 13035 15011
rect 13829 14977 13863 15011
rect 14657 14977 14691 15011
rect 15577 14977 15611 15011
rect 19993 14977 20027 15011
rect 1593 14909 1627 14943
rect 2329 14909 2363 14943
rect 6101 14909 6135 14943
rect 9689 14909 9723 14943
rect 9956 14909 9990 14943
rect 13645 14909 13679 14943
rect 14473 14909 14507 14943
rect 15301 14909 15335 14943
rect 16129 14909 16163 14943
rect 16313 14909 16347 14943
rect 16580 14909 16614 14943
rect 18061 14909 18095 14943
rect 19809 14909 19843 14943
rect 20545 14909 20579 14943
rect 2596 14841 2630 14875
rect 4537 14841 4571 14875
rect 8769 14841 8803 14875
rect 8861 14841 8895 14875
rect 11713 14841 11747 14875
rect 12909 14841 12943 14875
rect 13737 14841 13771 14875
rect 18306 14841 18340 14875
rect 20821 14841 20855 14875
rect 4629 14773 4663 14807
rect 5733 14773 5767 14807
rect 7757 14773 7791 14807
rect 7849 14773 7883 14807
rect 11805 14773 11839 14807
rect 12449 14773 12483 14807
rect 12817 14773 12851 14807
rect 14565 14773 14599 14807
rect 14933 14773 14967 14807
rect 15393 14773 15427 14807
rect 15945 14773 15979 14807
rect 2789 14569 2823 14603
rect 4353 14569 4387 14603
rect 4721 14569 4755 14603
rect 7021 14569 7055 14603
rect 7297 14569 7331 14603
rect 10333 14569 10367 14603
rect 11345 14569 11379 14603
rect 12173 14569 12207 14603
rect 13369 14569 13403 14603
rect 13921 14569 13955 14603
rect 14749 14569 14783 14603
rect 15301 14569 15335 14603
rect 18429 14569 18463 14603
rect 18889 14569 18923 14603
rect 19257 14569 19291 14603
rect 4813 14501 4847 14535
rect 2145 14433 2179 14467
rect 3157 14433 3191 14467
rect 5365 14433 5399 14467
rect 5621 14433 5655 14467
rect 7205 14433 7239 14467
rect 2237 14365 2271 14399
rect 2421 14365 2455 14399
rect 3249 14365 3283 14399
rect 3433 14365 3467 14399
rect 4905 14365 4939 14399
rect 19625 14501 19659 14535
rect 7656 14433 7690 14467
rect 11713 14433 11747 14467
rect 13277 14433 13311 14467
rect 14105 14433 14139 14467
rect 15669 14433 15703 14467
rect 16497 14433 16531 14467
rect 17316 14433 17350 14467
rect 18705 14433 18739 14467
rect 20269 14433 20303 14467
rect 7389 14365 7423 14399
rect 10425 14365 10459 14399
rect 10609 14365 10643 14399
rect 11805 14365 11839 14399
rect 11989 14365 12023 14399
rect 13461 14365 13495 14399
rect 15761 14365 15795 14399
rect 15853 14365 15887 14399
rect 17049 14365 17083 14399
rect 19717 14365 19751 14399
rect 19809 14365 19843 14399
rect 20913 14365 20947 14399
rect 1777 14297 1811 14331
rect 7297 14297 7331 14331
rect 6745 14229 6779 14263
rect 8769 14229 8803 14263
rect 9965 14229 9999 14263
rect 12909 14229 12943 14263
rect 16681 14229 16715 14263
rect 20453 14229 20487 14263
rect 1685 14025 1719 14059
rect 2881 14025 2915 14059
rect 6285 14025 6319 14059
rect 8401 14025 8435 14059
rect 10885 14025 10919 14059
rect 16957 14025 16991 14059
rect 18061 14025 18095 14059
rect 19349 14025 19383 14059
rect 20361 14025 20395 14059
rect 4629 13957 4663 13991
rect 13829 13957 13863 13991
rect 17877 13957 17911 13991
rect 2329 13889 2363 13923
rect 9505 13889 9539 13923
rect 9689 13889 9723 13923
rect 10517 13889 10551 13923
rect 10609 13889 10643 13923
rect 11437 13889 11471 13923
rect 16313 13889 16347 13923
rect 17417 13889 17451 13923
rect 17601 13889 17635 13923
rect 2145 13821 2179 13855
rect 2697 13821 2731 13855
rect 3249 13821 3283 13855
rect 4905 13821 4939 13855
rect 5161 13821 5195 13855
rect 7021 13821 7055 13855
rect 7288 13821 7322 13855
rect 11345 13821 11379 13855
rect 12449 13821 12483 13855
rect 12716 13821 12750 13855
rect 14105 13821 14139 13855
rect 18521 13889 18555 13923
rect 18613 13889 18647 13923
rect 19993 13889 20027 13923
rect 20913 13889 20947 13923
rect 19809 13821 19843 13855
rect 3516 13753 3550 13787
rect 9413 13753 9447 13787
rect 11253 13753 11287 13787
rect 14372 13753 14406 13787
rect 16221 13753 16255 13787
rect 17877 13753 17911 13787
rect 18429 13753 18463 13787
rect 20821 13753 20855 13787
rect 2053 13685 2087 13719
rect 9045 13685 9079 13719
rect 10057 13685 10091 13719
rect 10425 13685 10459 13719
rect 15485 13685 15519 13719
rect 15761 13685 15795 13719
rect 16129 13685 16163 13719
rect 17325 13685 17359 13719
rect 19717 13685 19751 13719
rect 20729 13685 20763 13719
rect 2237 13481 2271 13515
rect 6101 13481 6135 13515
rect 8309 13481 8343 13515
rect 8769 13481 8803 13515
rect 11345 13481 11379 13515
rect 12817 13481 12851 13515
rect 13369 13481 13403 13515
rect 14657 13481 14691 13515
rect 15485 13481 15519 13515
rect 15853 13481 15887 13515
rect 19993 13481 20027 13515
rect 20453 13481 20487 13515
rect 1777 13413 1811 13447
rect 3525 13413 3559 13447
rect 6561 13413 6595 13447
rect 8677 13413 8711 13447
rect 10232 13413 10266 13447
rect 13461 13413 13495 13447
rect 14565 13413 14599 13447
rect 15025 13413 15059 13447
rect 16856 13413 16890 13447
rect 18880 13413 18914 13447
rect 1501 13345 1535 13379
rect 2605 13345 2639 13379
rect 3249 13345 3283 13379
rect 4721 13345 4755 13379
rect 4813 13345 4847 13379
rect 6469 13345 6503 13379
rect 7481 13345 7515 13379
rect 9965 13345 9999 13379
rect 11704 13345 11738 13379
rect 15945 13345 15979 13379
rect 18613 13345 18647 13379
rect 20269 13345 20303 13379
rect 2697 13277 2731 13311
rect 2789 13277 2823 13311
rect 4905 13277 4939 13311
rect 6653 13277 6687 13311
rect 7573 13277 7607 13311
rect 7665 13277 7699 13311
rect 8861 13277 8895 13311
rect 11437 13277 11471 13311
rect 13645 13277 13679 13311
rect 14749 13277 14783 13311
rect 15025 13277 15059 13311
rect 16129 13277 16163 13311
rect 16589 13277 16623 13311
rect 13001 13209 13035 13243
rect 14197 13209 14231 13243
rect 4353 13141 4387 13175
rect 7113 13141 7147 13175
rect 17969 13141 18003 13175
rect 1869 12937 1903 12971
rect 3617 12937 3651 12971
rect 7941 12937 7975 12971
rect 8953 12937 8987 12971
rect 12633 12937 12667 12971
rect 15761 12937 15795 12971
rect 17785 12937 17819 12971
rect 19441 12937 19475 12971
rect 19993 12937 20027 12971
rect 6929 12869 6963 12903
rect 13001 12869 13035 12903
rect 16957 12869 16991 12903
rect 2237 12801 2271 12835
rect 4169 12801 4203 12835
rect 5181 12801 5215 12835
rect 7389 12801 7423 12835
rect 7573 12801 7607 12835
rect 8493 12801 8527 12835
rect 9505 12801 9539 12835
rect 13645 12801 13679 12835
rect 16037 12801 16071 12835
rect 17509 12801 17543 12835
rect 17785 12801 17819 12835
rect 20453 12801 20487 12835
rect 20545 12801 20579 12835
rect 1685 12733 1719 12767
rect 2504 12733 2538 12767
rect 7297 12733 7331 12767
rect 8309 12733 8343 12767
rect 9321 12733 9355 12767
rect 12173 12733 12207 12767
rect 12817 12733 12851 12767
rect 14381 12733 14415 12767
rect 14648 12733 14682 12767
rect 18061 12733 18095 12767
rect 18317 12733 18351 12767
rect 4997 12665 5031 12699
rect 8401 12665 8435 12699
rect 10333 12665 10367 12699
rect 13461 12665 13495 12699
rect 17325 12665 17359 12699
rect 20361 12665 20395 12699
rect 4629 12597 4663 12631
rect 5089 12597 5123 12631
rect 9413 12597 9447 12631
rect 11621 12597 11655 12631
rect 12173 12597 12207 12631
rect 13369 12597 13403 12631
rect 17417 12597 17451 12631
rect 2881 12393 2915 12427
rect 4261 12393 4295 12427
rect 4629 12393 4663 12427
rect 9505 12393 9539 12427
rect 9689 12393 9723 12427
rect 10057 12393 10091 12427
rect 12817 12393 12851 12427
rect 14657 12393 14691 12427
rect 17693 12393 17727 12427
rect 19809 12393 19843 12427
rect 20177 12393 20211 12427
rect 20913 12393 20947 12427
rect 1768 12325 1802 12359
rect 1501 12257 1535 12291
rect 4721 12257 4755 12291
rect 5897 12257 5931 12291
rect 7297 12257 7331 12291
rect 7564 12257 7598 12291
rect 18429 12325 18463 12359
rect 19349 12325 19383 12359
rect 11152 12257 11186 12291
rect 12725 12257 12759 12291
rect 13185 12257 13219 12291
rect 14013 12257 14047 12291
rect 14565 12257 14599 12291
rect 15301 12257 15335 12291
rect 16580 12257 16614 12291
rect 18337 12257 18371 12291
rect 19073 12257 19107 12291
rect 4813 12189 4847 12223
rect 5641 12189 5675 12223
rect 9505 12189 9539 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 10885 12189 10919 12223
rect 7021 12121 7055 12155
rect 8677 12121 8711 12155
rect 12265 12121 12299 12155
rect 13277 12189 13311 12223
rect 13461 12189 13495 12223
rect 14749 12189 14783 12223
rect 16313 12189 16347 12223
rect 18613 12189 18647 12223
rect 20269 12189 20303 12223
rect 20453 12189 20487 12223
rect 12725 12053 12759 12087
rect 13829 12053 13863 12087
rect 14197 12053 14231 12087
rect 17969 12053 18003 12087
rect 2329 11849 2363 11883
rect 5733 11849 5767 11883
rect 7849 11849 7883 11883
rect 10149 11849 10183 11883
rect 13829 11849 13863 11883
rect 14105 11849 14139 11883
rect 18981 11849 19015 11883
rect 19165 11849 19199 11883
rect 20177 11849 20211 11883
rect 16129 11781 16163 11815
rect 2973 11713 3007 11747
rect 3985 11713 4019 11747
rect 4353 11713 4387 11747
rect 7021 11713 7055 11747
rect 10609 11713 10643 11747
rect 10793 11713 10827 11747
rect 11897 11713 11931 11747
rect 14657 11713 14691 11747
rect 15669 11713 15703 11747
rect 16681 11713 16715 11747
rect 17417 11713 17451 11747
rect 18705 11713 18739 11747
rect 18981 11713 19015 11747
rect 19717 11713 19751 11747
rect 20729 11713 20763 11747
rect 8033 11645 8067 11679
rect 8217 11645 8251 11679
rect 8484 11645 8518 11679
rect 10517 11645 10551 11679
rect 12449 11645 12483 11679
rect 14473 11645 14507 11679
rect 17233 11645 17267 11679
rect 18521 11645 18555 11679
rect 19533 11645 19567 11679
rect 2697 11577 2731 11611
rect 4620 11577 4654 11611
rect 11713 11577 11747 11611
rect 12716 11577 12750 11611
rect 14565 11577 14599 11611
rect 16589 11577 16623 11611
rect 19625 11577 19659 11611
rect 20637 11577 20671 11611
rect 1501 11509 1535 11543
rect 2789 11509 2823 11543
rect 3341 11509 3375 11543
rect 3709 11509 3743 11543
rect 3801 11509 3835 11543
rect 9597 11509 9631 11543
rect 11345 11509 11379 11543
rect 11805 11509 11839 11543
rect 15117 11509 15151 11543
rect 15485 11509 15519 11543
rect 15577 11509 15611 11543
rect 16497 11509 16531 11543
rect 18153 11509 18187 11543
rect 18613 11509 18647 11543
rect 20545 11509 20579 11543
rect 1961 11305 1995 11339
rect 2973 11305 3007 11339
rect 4077 11305 4111 11339
rect 5549 11305 5583 11339
rect 6653 11305 6687 11339
rect 8217 11305 8251 11339
rect 10057 11305 10091 11339
rect 11161 11305 11195 11339
rect 11713 11305 11747 11339
rect 17141 11305 17175 11339
rect 17693 11305 17727 11339
rect 18705 11305 18739 11339
rect 19165 11305 19199 11339
rect 19717 11305 19751 11339
rect 20177 11305 20211 11339
rect 2329 11237 2363 11271
rect 2421 11237 2455 11271
rect 3341 11237 3375 11271
rect 3893 11237 3927 11271
rect 12992 11237 13026 11271
rect 18153 11237 18187 11271
rect 20085 11237 20119 11271
rect 1869 11169 1903 11203
rect 2513 11101 2547 11135
rect 3433 11101 3467 11135
rect 3617 11101 3651 11135
rect 4445 11169 4479 11203
rect 4537 11169 4571 11203
rect 5457 11169 5491 11203
rect 6561 11169 6595 11203
rect 7573 11169 7607 11203
rect 7665 11169 7699 11203
rect 8585 11169 8619 11203
rect 10149 11169 10183 11203
rect 11069 11169 11103 11203
rect 12081 11169 12115 11203
rect 15669 11169 15703 11203
rect 15761 11169 15795 11203
rect 16028 11169 16062 11203
rect 18061 11169 18095 11203
rect 19073 11169 19107 11203
rect 4629 11101 4663 11135
rect 5733 11101 5767 11135
rect 6745 11101 6779 11135
rect 7757 11101 7791 11135
rect 8677 11101 8711 11135
rect 8769 11101 8803 11135
rect 10241 11101 10275 11135
rect 11345 11101 11379 11135
rect 12173 11101 12207 11135
rect 12357 11101 12391 11135
rect 12725 11101 12759 11135
rect 15393 11101 15427 11135
rect 18245 11101 18279 11135
rect 19257 11101 19291 11135
rect 20269 11101 20303 11135
rect 6193 11033 6227 11067
rect 7205 11033 7239 11067
rect 10701 11033 10735 11067
rect 14105 11033 14139 11067
rect 3893 10965 3927 10999
rect 5089 10965 5123 10999
rect 9689 10965 9723 10999
rect 15393 10965 15427 10999
rect 15485 10965 15519 10999
rect 2881 10761 2915 10795
rect 4813 10761 4847 10795
rect 5733 10761 5767 10795
rect 7573 10761 7607 10795
rect 12633 10761 12667 10795
rect 13645 10761 13679 10795
rect 16037 10761 16071 10795
rect 16313 10761 16347 10795
rect 18613 10761 18647 10795
rect 19625 10761 19659 10795
rect 5089 10693 5123 10727
rect 7021 10693 7055 10727
rect 6285 10625 6319 10659
rect 6837 10625 6871 10659
rect 8217 10625 8251 10659
rect 10057 10625 10091 10659
rect 13277 10625 13311 10659
rect 14197 10625 14231 10659
rect 16865 10625 16899 10659
rect 18061 10625 18095 10659
rect 19165 10625 19199 10659
rect 20177 10625 20211 10659
rect 20821 10625 20855 10659
rect 1501 10557 1535 10591
rect 1768 10557 1802 10591
rect 3433 10557 3467 10591
rect 3700 10557 3734 10591
rect 5273 10557 5307 10591
rect 6101 10557 6135 10591
rect 7205 10557 7239 10591
rect 7941 10557 7975 10591
rect 9873 10557 9907 10591
rect 10517 10557 10551 10591
rect 13093 10557 13127 10591
rect 14013 10557 14047 10591
rect 14657 10557 14691 10591
rect 16773 10557 16807 10591
rect 18981 10557 19015 10591
rect 20637 10557 20671 10591
rect 10784 10489 10818 10523
rect 14924 10489 14958 10523
rect 19993 10489 20027 10523
rect 6193 10421 6227 10455
rect 6837 10421 6871 10455
rect 8033 10421 8067 10455
rect 9505 10421 9539 10455
rect 9965 10421 9999 10455
rect 11897 10421 11931 10455
rect 13001 10421 13035 10455
rect 14105 10421 14139 10455
rect 16681 10421 16715 10455
rect 19073 10421 19107 10455
rect 20085 10421 20119 10455
rect 1961 10217 1995 10251
rect 2973 10217 3007 10251
rect 4629 10217 4663 10251
rect 5549 10217 5583 10251
rect 7021 10217 7055 10251
rect 9321 10217 9355 10251
rect 10057 10217 10091 10251
rect 10149 10217 10183 10251
rect 17509 10217 17543 10251
rect 17877 10217 17911 10251
rect 18061 10217 18095 10251
rect 19257 10217 19291 10251
rect 2421 10149 2455 10183
rect 1409 10081 1443 10115
rect 2329 10081 2363 10115
rect 3341 10081 3375 10115
rect 4169 10081 4203 10115
rect 4997 10081 5031 10115
rect 2513 10013 2547 10047
rect 3433 10013 3467 10047
rect 3617 10013 3651 10047
rect 5089 10013 5123 10047
rect 5273 10013 5307 10047
rect 8208 10149 8242 10183
rect 11152 10149 11186 10183
rect 13737 10149 13771 10183
rect 13829 10149 13863 10183
rect 16396 10149 16430 10183
rect 19717 10149 19751 10183
rect 5908 10081 5942 10115
rect 7849 10081 7883 10115
rect 18429 10081 18463 10115
rect 19625 10081 19659 10115
rect 5641 10013 5675 10047
rect 7941 10013 7975 10047
rect 10241 10013 10275 10047
rect 10885 10013 10919 10047
rect 12725 10013 12759 10047
rect 13921 10013 13955 10047
rect 16129 10013 16163 10047
rect 18521 10013 18555 10047
rect 18613 10013 18647 10047
rect 19809 10013 19843 10047
rect 1593 9945 1627 9979
rect 5457 9945 5491 9979
rect 9689 9945 9723 9979
rect 7665 9877 7699 9911
rect 12265 9877 12299 9911
rect 13369 9877 13403 9911
rect 7021 9673 7055 9707
rect 1777 9605 1811 9639
rect 4169 9605 4203 9639
rect 4537 9605 4571 9639
rect 5641 9605 5675 9639
rect 12081 9605 12115 9639
rect 12449 9605 12483 9639
rect 16589 9605 16623 9639
rect 18889 9605 18923 9639
rect 2421 9537 2455 9571
rect 5181 9537 5215 9571
rect 6285 9537 6319 9571
rect 7665 9537 7699 9571
rect 10333 9537 10367 9571
rect 10517 9537 10551 9571
rect 13001 9537 13035 9571
rect 13553 9537 13587 9571
rect 17417 9537 17451 9571
rect 19533 9537 19567 9571
rect 20545 9537 20579 9571
rect 2145 9469 2179 9503
rect 2789 9469 2823 9503
rect 6101 9469 6135 9503
rect 8033 9469 8067 9503
rect 8289 9469 8323 9503
rect 10241 9469 10275 9503
rect 12265 9469 12299 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 15209 9469 15243 9503
rect 18153 9469 18187 9503
rect 19349 9469 19383 9503
rect 3034 9401 3068 9435
rect 4997 9401 5031 9435
rect 7481 9401 7515 9435
rect 13820 9401 13854 9435
rect 15476 9401 15510 9435
rect 17325 9401 17359 9435
rect 18429 9401 18463 9435
rect 20269 9401 20303 9435
rect 2237 9333 2271 9367
rect 4905 9333 4939 9367
rect 6009 9333 6043 9367
rect 7389 9333 7423 9367
rect 9413 9333 9447 9367
rect 9873 9333 9907 9367
rect 14933 9333 14967 9367
rect 16865 9333 16899 9367
rect 17233 9333 17267 9367
rect 19257 9333 19291 9367
rect 19901 9333 19935 9367
rect 20361 9333 20395 9367
rect 4261 9129 4295 9163
rect 4629 9129 4663 9163
rect 8493 9129 8527 9163
rect 14197 9129 14231 9163
rect 16773 9129 16807 9163
rect 1777 9061 1811 9095
rect 3525 9061 3559 9095
rect 7849 9061 7883 9095
rect 10324 9061 10358 9095
rect 1501 8993 1535 9027
rect 2605 8993 2639 9027
rect 3249 8993 3283 9027
rect 5641 8993 5675 9027
rect 7941 8993 7975 9027
rect 12081 8993 12115 9027
rect 12348 8993 12382 9027
rect 14565 8993 14599 9027
rect 15669 8993 15703 9027
rect 15761 8993 15795 9027
rect 16129 8993 16163 9027
rect 16681 8993 16715 9027
rect 17325 8993 17359 9027
rect 18788 8993 18822 9027
rect 2697 8925 2731 8959
rect 2881 8925 2915 8959
rect 4721 8925 4755 8959
rect 4905 8925 4939 8959
rect 5733 8925 5767 8959
rect 5917 8925 5951 8959
rect 8033 8925 8067 8959
rect 10057 8925 10091 8959
rect 14657 8925 14691 8959
rect 14841 8925 14875 8959
rect 15945 8925 15979 8959
rect 16865 8925 16899 8959
rect 18521 8925 18555 8959
rect 2237 8857 2271 8891
rect 13461 8857 13495 8891
rect 16129 8857 16163 8891
rect 19901 8857 19935 8891
rect 5273 8789 5307 8823
rect 7481 8789 7515 8823
rect 11437 8789 11471 8823
rect 15301 8789 15335 8823
rect 16313 8789 16347 8823
rect 3065 8585 3099 8619
rect 4629 8585 4663 8619
rect 5733 8585 5767 8619
rect 14105 8585 14139 8619
rect 19441 8585 19475 8619
rect 3617 8517 3651 8551
rect 16589 8517 16623 8551
rect 4169 8449 4203 8483
rect 5273 8449 5307 8483
rect 6285 8449 6319 8483
rect 7665 8449 7699 8483
rect 10701 8449 10735 8483
rect 10793 8449 10827 8483
rect 11805 8449 11839 8483
rect 14749 8449 14783 8483
rect 15853 8449 15887 8483
rect 17049 8449 17083 8483
rect 17233 8449 17267 8483
rect 20453 8449 20487 8483
rect 1685 8381 1719 8415
rect 5089 8381 5123 8415
rect 6193 8381 6227 8415
rect 8585 8381 8619 8415
rect 8841 8381 8875 8415
rect 11713 8381 11747 8415
rect 12449 8381 12483 8415
rect 14565 8381 14599 8415
rect 16957 8381 16991 8415
rect 18061 8381 18095 8415
rect 1952 8313 1986 8347
rect 3985 8313 4019 8347
rect 6101 8313 6135 8347
rect 10609 8313 10643 8347
rect 11621 8313 11655 8347
rect 12716 8313 12750 8347
rect 14473 8313 14507 8347
rect 18328 8313 18362 8347
rect 20177 8313 20211 8347
rect 20821 8313 20855 8347
rect 4077 8245 4111 8279
rect 4997 8245 5031 8279
rect 7021 8245 7055 8279
rect 7389 8245 7423 8279
rect 7481 8245 7515 8279
rect 9965 8245 9999 8279
rect 10241 8245 10275 8279
rect 11253 8245 11287 8279
rect 13829 8245 13863 8279
rect 15301 8245 15335 8279
rect 15669 8245 15703 8279
rect 15761 8245 15795 8279
rect 19809 8245 19843 8279
rect 20269 8245 20303 8279
rect 1777 8041 1811 8075
rect 2237 8041 2271 8075
rect 2789 8041 2823 8075
rect 5457 8041 5491 8075
rect 7757 8041 7791 8075
rect 8309 8041 8343 8075
rect 8769 8041 8803 8075
rect 10149 8041 10183 8075
rect 10701 8041 10735 8075
rect 15669 8041 15703 8075
rect 19165 8041 19199 8075
rect 20177 8041 20211 8075
rect 4997 7973 5031 8007
rect 2145 7905 2179 7939
rect 3157 7905 3191 7939
rect 3249 7905 3283 7939
rect 10057 7973 10091 8007
rect 11069 7973 11103 8007
rect 15761 7973 15795 8007
rect 17294 7973 17328 8007
rect 20269 7973 20303 8007
rect 5897 7905 5931 7939
rect 7665 7905 7699 7939
rect 8677 7905 8711 7939
rect 13001 7905 13035 7939
rect 19073 7905 19107 7939
rect 2329 7837 2363 7871
rect 3433 7837 3467 7871
rect 5089 7837 5123 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 5641 7837 5675 7871
rect 7941 7837 7975 7871
rect 8861 7837 8895 7871
rect 10241 7837 10275 7871
rect 11161 7837 11195 7871
rect 11345 7837 11379 7871
rect 13093 7837 13127 7871
rect 13277 7837 13311 7871
rect 15853 7837 15887 7871
rect 17049 7837 17083 7871
rect 19349 7837 19383 7871
rect 20453 7837 20487 7871
rect 7021 7769 7055 7803
rect 7297 7769 7331 7803
rect 9689 7769 9723 7803
rect 15301 7769 15335 7803
rect 4629 7701 4663 7735
rect 12633 7701 12667 7735
rect 18429 7701 18463 7735
rect 18705 7701 18739 7735
rect 19809 7701 19843 7735
rect 18061 7497 18095 7531
rect 19257 7497 19291 7531
rect 20269 7497 20303 7531
rect 3709 7429 3743 7463
rect 3985 7429 4019 7463
rect 9873 7429 9907 7463
rect 4537 7361 4571 7395
rect 4997 7361 5031 7395
rect 18613 7361 18647 7395
rect 19717 7361 19751 7395
rect 19809 7361 19843 7395
rect 20729 7361 20763 7395
rect 20821 7361 20855 7395
rect 2329 7293 2363 7327
rect 2596 7293 2630 7327
rect 4353 7293 4387 7327
rect 6837 7293 6871 7327
rect 7093 7293 7127 7327
rect 8493 7293 8527 7327
rect 18429 7293 18463 7327
rect 19625 7293 19659 7327
rect 20637 7293 20671 7327
rect 5264 7225 5298 7259
rect 8760 7225 8794 7259
rect 4445 7157 4479 7191
rect 6377 7157 6411 7191
rect 8217 7157 8251 7191
rect 18521 7157 18555 7191
rect 2789 6953 2823 6987
rect 17969 6953 18003 6987
rect 3157 6817 3191 6851
rect 5365 6817 5399 6851
rect 6009 6817 6043 6851
rect 16589 6817 16623 6851
rect 16856 6817 16890 6851
rect 19064 6817 19098 6851
rect 3249 6749 3283 6783
rect 3341 6749 3375 6783
rect 5457 6749 5491 6783
rect 5549 6749 5583 6783
rect 18797 6749 18831 6783
rect 4997 6613 5031 6647
rect 20177 6613 20211 6647
rect 2973 6409 3007 6443
rect 5089 6409 5123 6443
rect 20453 6409 20487 6443
rect 1593 6273 1627 6307
rect 3249 6273 3283 6307
rect 5549 6273 5583 6307
rect 5733 6273 5767 6307
rect 18521 6273 18555 6307
rect 19073 6273 19107 6307
rect 5457 6205 5491 6239
rect 18337 6205 18371 6239
rect 1860 6137 1894 6171
rect 19340 6137 19374 6171
rect 20729 6069 20763 6103
rect 20177 5729 20211 5763
rect 20269 5661 20303 5695
rect 20361 5661 20395 5695
rect 19625 5593 19659 5627
rect 19809 5525 19843 5559
rect 19809 5321 19843 5355
rect 20269 5185 20303 5219
rect 20453 5185 20487 5219
rect 20177 5117 20211 5151
rect 4905 3009 4939 3043
rect 4629 2941 4663 2975
rect 5549 2941 5583 2975
rect 15209 2941 15243 2975
rect 5825 2873 5859 2907
rect 15485 2873 15519 2907
<< metal1 >>
rect 4062 20952 4068 21004
rect 4120 20992 4126 21004
rect 5718 20992 5724 21004
rect 4120 20964 5724 20992
rect 4120 20952 4126 20964
rect 5718 20952 5724 20964
rect 5776 20952 5782 21004
rect 9766 20680 9772 20732
rect 9824 20720 9830 20732
rect 10318 20720 10324 20732
rect 9824 20692 10324 20720
rect 9824 20680 9830 20692
rect 10318 20680 10324 20692
rect 10376 20680 10382 20732
rect 14366 20612 14372 20664
rect 14424 20652 14430 20664
rect 19610 20652 19616 20664
rect 14424 20624 19616 20652
rect 14424 20612 14430 20624
rect 19610 20612 19616 20624
rect 19668 20612 19674 20664
rect 12250 20544 12256 20596
rect 12308 20584 12314 20596
rect 16666 20584 16672 20596
rect 12308 20556 16672 20584
rect 12308 20544 12314 20556
rect 16666 20544 16672 20556
rect 16724 20544 16730 20596
rect 15654 20408 15660 20460
rect 15712 20448 15718 20460
rect 17862 20448 17868 20460
rect 15712 20420 17868 20448
rect 15712 20408 15718 20420
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 10226 20340 10232 20392
rect 10284 20380 10290 20392
rect 17678 20380 17684 20392
rect 10284 20352 17684 20380
rect 10284 20340 10290 20352
rect 17678 20340 17684 20352
rect 17736 20340 17742 20392
rect 14550 20272 14556 20324
rect 14608 20312 14614 20324
rect 17034 20312 17040 20324
rect 14608 20284 17040 20312
rect 14608 20272 14614 20284
rect 17034 20272 17040 20284
rect 17092 20272 17098 20324
rect 15102 20204 15108 20256
rect 15160 20244 15166 20256
rect 19150 20244 19156 20256
rect 15160 20216 19156 20244
rect 15160 20204 15166 20216
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 2041 20043 2099 20049
rect 2041 20009 2053 20043
rect 2087 20040 2099 20043
rect 2774 20040 2780 20052
rect 2087 20012 2780 20040
rect 2087 20009 2099 20012
rect 2041 20003 2099 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 9033 20043 9091 20049
rect 9033 20009 9045 20043
rect 9079 20040 9091 20043
rect 9769 20043 9827 20049
rect 9769 20040 9781 20043
rect 9079 20012 9781 20040
rect 9079 20009 9091 20012
rect 9033 20003 9091 20009
rect 9769 20009 9781 20012
rect 9815 20009 9827 20043
rect 10226 20040 10232 20052
rect 10187 20012 10232 20040
rect 9769 20003 9827 20009
rect 10226 20000 10232 20012
rect 10284 20000 10290 20052
rect 14366 20000 14372 20052
rect 14424 20040 14430 20052
rect 14461 20043 14519 20049
rect 14461 20040 14473 20043
rect 14424 20012 14473 20040
rect 14424 20000 14430 20012
rect 14461 20009 14473 20012
rect 14507 20009 14519 20043
rect 14461 20003 14519 20009
rect 15013 20043 15071 20049
rect 15013 20009 15025 20043
rect 15059 20040 15071 20043
rect 15102 20040 15108 20052
rect 15059 20012 15108 20040
rect 15059 20009 15071 20012
rect 15013 20003 15071 20009
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15654 20040 15660 20052
rect 15615 20012 15660 20040
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 16761 20043 16819 20049
rect 16761 20009 16773 20043
rect 16807 20040 16819 20043
rect 17494 20040 17500 20052
rect 16807 20012 17500 20040
rect 16807 20009 16819 20012
rect 16761 20003 16819 20009
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 18506 20040 18512 20052
rect 18467 20012 18512 20040
rect 18506 20000 18512 20012
rect 18564 20000 18570 20052
rect 19058 20040 19064 20052
rect 19019 20012 19064 20040
rect 19058 20000 19064 20012
rect 19116 20000 19122 20052
rect 19242 20000 19248 20052
rect 19300 20040 19306 20052
rect 19613 20043 19671 20049
rect 19613 20040 19625 20043
rect 19300 20012 19625 20040
rect 19300 20000 19306 20012
rect 19613 20009 19625 20012
rect 19659 20009 19671 20043
rect 19613 20003 19671 20009
rect 7469 19975 7527 19981
rect 7469 19941 7481 19975
rect 7515 19972 7527 19975
rect 8478 19972 8484 19984
rect 7515 19944 8484 19972
rect 7515 19941 7527 19944
rect 7469 19935 7527 19941
rect 8478 19932 8484 19944
rect 8536 19932 8542 19984
rect 15562 19932 15568 19984
rect 15620 19972 15626 19984
rect 15620 19944 16620 19972
rect 15620 19932 15626 19944
rect 1857 19907 1915 19913
rect 1857 19873 1869 19907
rect 1903 19873 1915 19907
rect 1857 19867 1915 19873
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19904 2467 19907
rect 3694 19904 3700 19916
rect 2455 19876 3700 19904
rect 2455 19873 2467 19876
rect 2409 19867 2467 19873
rect 1872 19836 1900 19867
rect 3694 19864 3700 19876
rect 3752 19864 3758 19916
rect 7742 19864 7748 19916
rect 7800 19904 7806 19916
rect 8113 19907 8171 19913
rect 8113 19904 8125 19907
rect 7800 19876 8125 19904
rect 7800 19864 7806 19876
rect 8113 19873 8125 19876
rect 8159 19873 8171 19907
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 8113 19867 8171 19873
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 11977 19907 12035 19913
rect 11977 19873 11989 19907
rect 12023 19904 12035 19907
rect 12158 19904 12164 19916
rect 12023 19876 12164 19904
rect 12023 19873 12035 19876
rect 11977 19867 12035 19873
rect 12158 19864 12164 19876
rect 12216 19864 12222 19916
rect 12986 19904 12992 19916
rect 12947 19876 12992 19904
rect 12986 19864 12992 19876
rect 13044 19864 13050 19916
rect 13538 19864 13544 19916
rect 13596 19904 13602 19916
rect 13725 19907 13783 19913
rect 13725 19904 13737 19907
rect 13596 19876 13737 19904
rect 13596 19864 13602 19876
rect 13725 19873 13737 19876
rect 13771 19873 13783 19907
rect 13725 19867 13783 19873
rect 13998 19864 14004 19916
rect 14056 19904 14062 19916
rect 14277 19907 14335 19913
rect 14277 19904 14289 19907
rect 14056 19876 14289 19904
rect 14056 19864 14062 19876
rect 14277 19873 14289 19876
rect 14323 19873 14335 19907
rect 14826 19904 14832 19916
rect 14787 19876 14832 19904
rect 14277 19867 14335 19873
rect 14826 19864 14832 19876
rect 14884 19864 14890 19916
rect 15470 19904 15476 19916
rect 15431 19876 15476 19904
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 16592 19913 16620 19944
rect 16850 19932 16856 19984
rect 16908 19972 16914 19984
rect 16908 19944 18920 19972
rect 16908 19932 16914 19944
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 16393 19907 16451 19913
rect 16393 19904 16405 19907
rect 16071 19876 16405 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 16393 19873 16405 19876
rect 16439 19873 16451 19907
rect 16393 19867 16451 19873
rect 16577 19907 16635 19913
rect 16577 19873 16589 19907
rect 16623 19873 16635 19907
rect 16577 19867 16635 19873
rect 16666 19864 16672 19916
rect 16724 19904 16730 19916
rect 17313 19907 17371 19913
rect 17313 19904 17325 19907
rect 16724 19876 17325 19904
rect 16724 19864 16730 19876
rect 17313 19873 17325 19876
rect 17359 19873 17371 19907
rect 17313 19867 17371 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18506 19904 18512 19916
rect 18371 19876 18512 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18506 19864 18512 19876
rect 18564 19864 18570 19916
rect 18892 19913 18920 19944
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19873 18935 19907
rect 18877 19867 18935 19873
rect 19429 19907 19487 19913
rect 19429 19873 19441 19907
rect 19475 19904 19487 19907
rect 19518 19904 19524 19916
rect 19475 19876 19524 19904
rect 19475 19873 19487 19876
rect 19429 19867 19487 19873
rect 19518 19864 19524 19876
rect 19576 19864 19582 19916
rect 19981 19907 20039 19913
rect 19981 19873 19993 19907
rect 20027 19904 20039 19907
rect 20254 19904 20260 19916
rect 20027 19876 20260 19904
rect 20027 19873 20039 19876
rect 19981 19867 20039 19873
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 20533 19907 20591 19913
rect 20533 19873 20545 19907
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 4982 19836 4988 19848
rect 1872 19808 4988 19836
rect 4982 19796 4988 19808
rect 5040 19796 5046 19848
rect 7558 19836 7564 19848
rect 7519 19808 7564 19836
rect 7558 19796 7564 19808
rect 7616 19796 7622 19848
rect 7653 19839 7711 19845
rect 7653 19805 7665 19839
rect 7699 19805 7711 19839
rect 9122 19836 9128 19848
rect 9083 19808 9128 19836
rect 7653 19799 7711 19805
rect 6914 19728 6920 19780
rect 6972 19768 6978 19780
rect 7668 19768 7696 19799
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 10226 19836 10232 19848
rect 9355 19808 10232 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 10318 19796 10324 19848
rect 10376 19836 10382 19848
rect 13078 19836 13084 19848
rect 10376 19808 10421 19836
rect 13039 19808 13084 19836
rect 10376 19796 10382 19808
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 18782 19836 18788 19848
rect 13228 19808 13273 19836
rect 17420 19808 18788 19836
rect 13228 19796 13234 19808
rect 6972 19740 7696 19768
rect 8297 19771 8355 19777
rect 6972 19728 6978 19740
rect 8297 19737 8309 19771
rect 8343 19768 8355 19771
rect 14550 19768 14556 19780
rect 8343 19740 14556 19768
rect 8343 19737 8355 19740
rect 8297 19731 8355 19737
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 16209 19771 16267 19777
rect 16209 19737 16221 19771
rect 16255 19768 16267 19771
rect 17420 19768 17448 19808
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 20548 19836 20576 19867
rect 19444 19808 20576 19836
rect 19444 19780 19472 19808
rect 16255 19740 17448 19768
rect 17497 19771 17555 19777
rect 16255 19737 16267 19740
rect 16209 19731 16267 19737
rect 17497 19737 17509 19771
rect 17543 19768 17555 19771
rect 18322 19768 18328 19780
rect 17543 19740 18328 19768
rect 17543 19737 17555 19740
rect 17497 19731 17555 19737
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 19426 19728 19432 19780
rect 19484 19728 19490 19780
rect 20162 19768 20168 19780
rect 20123 19740 20168 19768
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 2590 19700 2596 19712
rect 2551 19672 2596 19700
rect 2590 19660 2596 19672
rect 2648 19660 2654 19712
rect 7101 19703 7159 19709
rect 7101 19669 7113 19703
rect 7147 19700 7159 19703
rect 7466 19700 7472 19712
rect 7147 19672 7472 19700
rect 7147 19669 7159 19672
rect 7101 19663 7159 19669
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 8665 19703 8723 19709
rect 8665 19669 8677 19703
rect 8711 19700 8723 19703
rect 9582 19700 9588 19712
rect 8711 19672 9588 19700
rect 8711 19669 8723 19672
rect 8665 19663 8723 19669
rect 9582 19660 9588 19672
rect 9640 19660 9646 19712
rect 12161 19703 12219 19709
rect 12161 19669 12173 19703
rect 12207 19700 12219 19703
rect 12250 19700 12256 19712
rect 12207 19672 12256 19700
rect 12207 19669 12219 19672
rect 12161 19663 12219 19669
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12621 19703 12679 19709
rect 12621 19669 12633 19703
rect 12667 19700 12679 19703
rect 13814 19700 13820 19712
rect 12667 19672 13820 19700
rect 12667 19669 12679 19672
rect 12621 19663 12679 19669
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 13906 19660 13912 19712
rect 13964 19700 13970 19712
rect 16393 19703 16451 19709
rect 13964 19672 14009 19700
rect 13964 19660 13970 19672
rect 16393 19669 16405 19703
rect 16439 19700 16451 19703
rect 17954 19700 17960 19712
rect 16439 19672 17960 19700
rect 16439 19669 16451 19672
rect 16393 19663 16451 19669
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 20717 19703 20775 19709
rect 20717 19700 20729 19703
rect 20680 19672 20729 19700
rect 20680 19660 20686 19672
rect 20717 19669 20729 19672
rect 20763 19669 20775 19703
rect 20717 19663 20775 19669
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 3510 19496 3516 19508
rect 3471 19468 3516 19496
rect 3510 19456 3516 19468
rect 3568 19456 3574 19508
rect 5718 19496 5724 19508
rect 5679 19468 5724 19496
rect 5718 19456 5724 19468
rect 5776 19456 5782 19508
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 7926 19496 7932 19508
rect 7616 19468 7932 19496
rect 7616 19456 7622 19468
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 12529 19499 12587 19505
rect 12529 19465 12541 19499
rect 12575 19496 12587 19499
rect 13078 19496 13084 19508
rect 12575 19468 13084 19496
rect 12575 19465 12587 19468
rect 12529 19459 12587 19465
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 13906 19456 13912 19508
rect 13964 19496 13970 19508
rect 19610 19496 19616 19508
rect 13964 19468 19012 19496
rect 19571 19468 19616 19496
rect 13964 19456 13970 19468
rect 7742 19428 7748 19440
rect 7300 19400 7748 19428
rect 7300 19369 7328 19400
rect 7742 19388 7748 19400
rect 7800 19388 7806 19440
rect 14826 19388 14832 19440
rect 14884 19428 14890 19440
rect 14884 19400 18920 19428
rect 14884 19388 14890 19400
rect 7285 19363 7343 19369
rect 3252 19332 3464 19360
rect 198 19252 204 19304
rect 256 19292 262 19304
rect 1857 19295 1915 19301
rect 1857 19292 1869 19295
rect 256 19264 1869 19292
rect 256 19252 262 19264
rect 1857 19261 1869 19264
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 2409 19295 2467 19301
rect 2409 19261 2421 19295
rect 2455 19292 2467 19295
rect 3252 19292 3280 19332
rect 2455 19264 3280 19292
rect 3329 19295 3387 19301
rect 2455 19261 2467 19264
rect 2409 19255 2467 19261
rect 3329 19261 3341 19295
rect 3375 19261 3387 19295
rect 3329 19255 3387 19261
rect 2866 19224 2872 19236
rect 2608 19196 2872 19224
rect 2038 19156 2044 19168
rect 1999 19128 2044 19156
rect 2038 19116 2044 19128
rect 2096 19116 2102 19168
rect 2608 19165 2636 19196
rect 2866 19184 2872 19196
rect 2924 19184 2930 19236
rect 2593 19159 2651 19165
rect 2593 19125 2605 19159
rect 2639 19125 2651 19159
rect 3344 19156 3372 19255
rect 3436 19224 3464 19332
rect 7285 19329 7297 19363
rect 7331 19329 7343 19363
rect 7285 19323 7343 19329
rect 10226 19320 10232 19372
rect 10284 19360 10290 19372
rect 12437 19363 12495 19369
rect 10284 19332 10456 19360
rect 10284 19320 10290 19332
rect 3970 19292 3976 19304
rect 3931 19264 3976 19292
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 5166 19292 5172 19304
rect 4080 19264 5172 19292
rect 4080 19224 4108 19264
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5537 19295 5595 19301
rect 5537 19261 5549 19295
rect 5583 19292 5595 19295
rect 6086 19292 6092 19304
rect 5583 19264 6092 19292
rect 5583 19261 5595 19264
rect 5537 19255 5595 19261
rect 6086 19252 6092 19264
rect 6144 19252 6150 19304
rect 6178 19252 6184 19304
rect 6236 19292 6242 19304
rect 6822 19292 6828 19304
rect 6236 19264 6828 19292
rect 6236 19252 6242 19264
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 7006 19292 7012 19304
rect 6967 19264 7012 19292
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 7745 19295 7803 19301
rect 7745 19292 7757 19295
rect 7668 19264 7757 19292
rect 3436 19196 4108 19224
rect 4709 19227 4767 19233
rect 4709 19193 4721 19227
rect 4755 19224 4767 19227
rect 7558 19224 7564 19236
rect 4755 19196 7564 19224
rect 4755 19193 4767 19196
rect 4709 19187 4767 19193
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 6362 19156 6368 19168
rect 3344 19128 6368 19156
rect 2593 19119 2651 19125
rect 6362 19116 6368 19128
rect 6420 19116 6426 19168
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 7668 19156 7696 19264
rect 7745 19261 7757 19264
rect 7791 19292 7803 19295
rect 9582 19292 9588 19304
rect 7791 19264 9444 19292
rect 9543 19264 9588 19292
rect 7791 19261 7803 19264
rect 7745 19255 7803 19261
rect 7990 19227 8048 19233
rect 7990 19224 8002 19227
rect 7760 19196 8002 19224
rect 7760 19168 7788 19196
rect 7990 19193 8002 19196
rect 8036 19193 8048 19227
rect 7990 19187 8048 19193
rect 8110 19184 8116 19236
rect 8168 19224 8174 19236
rect 9306 19224 9312 19236
rect 8168 19196 9312 19224
rect 8168 19184 8174 19196
rect 9306 19184 9312 19196
rect 9364 19184 9370 19236
rect 9416 19224 9444 19264
rect 9582 19252 9588 19264
rect 9640 19252 9646 19304
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 9950 19292 9956 19304
rect 9824 19264 9956 19292
rect 9824 19252 9830 19264
rect 9950 19252 9956 19264
rect 10008 19252 10014 19304
rect 10137 19295 10195 19301
rect 10137 19261 10149 19295
rect 10183 19292 10195 19295
rect 10321 19295 10379 19301
rect 10321 19292 10333 19295
rect 10183 19264 10333 19292
rect 10183 19261 10195 19264
rect 10137 19255 10195 19261
rect 10321 19261 10333 19264
rect 10367 19261 10379 19295
rect 10428 19292 10456 19332
rect 12437 19329 12449 19363
rect 12483 19360 12495 19363
rect 13173 19363 13231 19369
rect 13173 19360 13185 19363
rect 12483 19332 13185 19360
rect 12483 19329 12495 19332
rect 12437 19323 12495 19329
rect 13173 19329 13185 19332
rect 13219 19360 13231 19363
rect 13262 19360 13268 19372
rect 13219 19332 13268 19360
rect 13219 19329 13231 19332
rect 13173 19323 13231 19329
rect 13262 19320 13268 19332
rect 13320 19320 13326 19372
rect 17494 19360 17500 19372
rect 17455 19332 17500 19360
rect 17494 19320 17500 19332
rect 17552 19320 17558 19372
rect 18892 19369 18920 19400
rect 18877 19363 18935 19369
rect 18877 19329 18889 19363
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 10577 19295 10635 19301
rect 10577 19292 10589 19295
rect 10428 19264 10589 19292
rect 10321 19255 10379 19261
rect 10577 19261 10589 19264
rect 10623 19292 10635 19295
rect 10962 19292 10968 19304
rect 10623 19264 10968 19292
rect 10623 19261 10635 19264
rect 10577 19255 10635 19261
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11974 19292 11980 19304
rect 11112 19264 11980 19292
rect 11112 19252 11118 19264
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 12250 19252 12256 19304
rect 12308 19292 12314 19304
rect 12308 19264 13308 19292
rect 12308 19252 12314 19264
rect 9674 19224 9680 19236
rect 9416 19196 9680 19224
rect 9674 19184 9680 19196
rect 9732 19184 9738 19236
rect 9861 19227 9919 19233
rect 9861 19193 9873 19227
rect 9907 19224 9919 19227
rect 10410 19224 10416 19236
rect 9907 19196 10416 19224
rect 9907 19193 9919 19196
rect 9861 19187 9919 19193
rect 10410 19184 10416 19196
rect 10468 19184 10474 19236
rect 10778 19184 10784 19236
rect 10836 19224 10842 19236
rect 12802 19224 12808 19236
rect 10836 19196 12808 19224
rect 10836 19184 10842 19196
rect 12802 19184 12808 19196
rect 12860 19224 12866 19236
rect 12989 19227 13047 19233
rect 12989 19224 13001 19227
rect 12860 19196 13001 19224
rect 12860 19184 12866 19196
rect 12989 19193 13001 19196
rect 13035 19193 13047 19227
rect 13280 19224 13308 19264
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 14001 19295 14059 19301
rect 14001 19292 14013 19295
rect 13872 19264 14013 19292
rect 13872 19252 13878 19264
rect 14001 19261 14013 19264
rect 14047 19261 14059 19295
rect 14001 19255 14059 19261
rect 14737 19295 14795 19301
rect 14737 19261 14749 19295
rect 14783 19292 14795 19295
rect 15102 19292 15108 19304
rect 14783 19264 15108 19292
rect 14783 19261 14795 19264
rect 14737 19255 14795 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15286 19292 15292 19304
rect 15247 19264 15292 19292
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 16025 19295 16083 19301
rect 16025 19261 16037 19295
rect 16071 19292 16083 19295
rect 16574 19292 16580 19304
rect 16071 19264 16580 19292
rect 16071 19261 16083 19264
rect 16025 19255 16083 19261
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 17402 19252 17408 19304
rect 17460 19292 17466 19304
rect 18141 19295 18199 19301
rect 18141 19292 18153 19295
rect 17460 19264 18153 19292
rect 17460 19252 17466 19264
rect 18141 19261 18153 19264
rect 18187 19261 18199 19295
rect 18141 19255 18199 19261
rect 18693 19295 18751 19301
rect 18693 19261 18705 19295
rect 18739 19292 18751 19295
rect 18782 19292 18788 19304
rect 18739 19264 18788 19292
rect 18739 19261 18751 19264
rect 18693 19255 18751 19261
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 14090 19224 14096 19236
rect 13280 19196 14096 19224
rect 12989 19187 13047 19193
rect 14090 19184 14096 19196
rect 14148 19184 14154 19236
rect 14277 19227 14335 19233
rect 14277 19193 14289 19227
rect 14323 19224 14335 19227
rect 15470 19224 15476 19236
rect 14323 19196 15476 19224
rect 14323 19193 14335 19196
rect 14277 19187 14335 19193
rect 15470 19184 15476 19196
rect 15528 19184 15534 19236
rect 15565 19227 15623 19233
rect 15565 19193 15577 19227
rect 15611 19224 15623 19227
rect 16666 19224 16672 19236
rect 15611 19196 16672 19224
rect 15611 19193 15623 19196
rect 15565 19187 15623 19193
rect 16666 19184 16672 19196
rect 16724 19184 16730 19236
rect 16758 19184 16764 19236
rect 16816 19224 16822 19236
rect 17313 19227 17371 19233
rect 17313 19224 17325 19227
rect 16816 19196 17325 19224
rect 16816 19184 16822 19196
rect 17313 19193 17325 19196
rect 17359 19193 17371 19227
rect 17313 19187 17371 19193
rect 17678 19184 17684 19236
rect 17736 19224 17742 19236
rect 18984 19224 19012 19468
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 19337 19295 19395 19301
rect 19337 19261 19349 19295
rect 19383 19292 19395 19295
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 19383 19264 19441 19292
rect 19383 19261 19395 19264
rect 19337 19255 19395 19261
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19429 19255 19487 19261
rect 19610 19252 19616 19304
rect 19668 19292 19674 19304
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19668 19264 19993 19292
rect 19668 19252 19674 19264
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 19981 19255 20039 19261
rect 20070 19252 20076 19304
rect 20128 19292 20134 19304
rect 20533 19295 20591 19301
rect 20533 19292 20545 19295
rect 20128 19264 20545 19292
rect 20128 19252 20134 19264
rect 20533 19261 20545 19264
rect 20579 19261 20591 19295
rect 20533 19255 20591 19261
rect 22094 19224 22100 19236
rect 17736 19196 18920 19224
rect 18984 19196 22100 19224
rect 17736 19184 17742 19196
rect 7340 19128 7696 19156
rect 7340 19116 7346 19128
rect 7742 19116 7748 19168
rect 7800 19116 7806 19168
rect 9125 19159 9183 19165
rect 9125 19125 9137 19159
rect 9171 19156 9183 19159
rect 10042 19156 10048 19168
rect 9171 19128 10048 19156
rect 9171 19125 9183 19128
rect 9125 19119 9183 19125
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 10137 19159 10195 19165
rect 10137 19125 10149 19159
rect 10183 19156 10195 19159
rect 10226 19156 10232 19168
rect 10183 19128 10232 19156
rect 10183 19125 10195 19128
rect 10137 19119 10195 19125
rect 10226 19116 10232 19128
rect 10284 19156 10290 19168
rect 11514 19156 11520 19168
rect 10284 19128 11520 19156
rect 10284 19116 10290 19128
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 11701 19159 11759 19165
rect 11701 19125 11713 19159
rect 11747 19156 11759 19159
rect 11974 19156 11980 19168
rect 11747 19128 11980 19156
rect 11747 19125 11759 19128
rect 11701 19119 11759 19125
rect 11974 19116 11980 19128
rect 12032 19156 12038 19168
rect 12437 19159 12495 19165
rect 12437 19156 12449 19159
rect 12032 19128 12449 19156
rect 12032 19116 12038 19128
rect 12437 19125 12449 19128
rect 12483 19125 12495 19159
rect 12894 19156 12900 19168
rect 12855 19128 12900 19156
rect 12437 19119 12495 19125
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 13541 19159 13599 19165
rect 13541 19156 13553 19159
rect 13136 19128 13553 19156
rect 13136 19116 13142 19128
rect 13541 19125 13553 19128
rect 13587 19125 13599 19159
rect 13541 19119 13599 19125
rect 14921 19159 14979 19165
rect 14921 19125 14933 19159
rect 14967 19156 14979 19159
rect 15378 19156 15384 19168
rect 14967 19128 15384 19156
rect 14967 19125 14979 19128
rect 14921 19119 14979 19125
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 16209 19159 16267 19165
rect 16209 19156 16221 19159
rect 15804 19128 16221 19156
rect 15804 19116 15810 19128
rect 16209 19125 16221 19128
rect 16255 19125 16267 19159
rect 16209 19119 16267 19125
rect 16853 19159 16911 19165
rect 16853 19125 16865 19159
rect 16899 19156 16911 19159
rect 16942 19156 16948 19168
rect 16899 19128 16948 19156
rect 16899 19125 16911 19128
rect 16853 19119 16911 19125
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 17218 19156 17224 19168
rect 17179 19128 17224 19156
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 18325 19159 18383 19165
rect 18325 19125 18337 19159
rect 18371 19156 18383 19159
rect 18598 19156 18604 19168
rect 18371 19128 18604 19156
rect 18371 19125 18383 19128
rect 18325 19119 18383 19125
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 18892 19156 18920 19196
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 19337 19159 19395 19165
rect 19337 19156 19349 19159
rect 18892 19128 19349 19156
rect 19337 19125 19349 19128
rect 19383 19125 19395 19159
rect 20162 19156 20168 19168
rect 20123 19128 20168 19156
rect 19337 19119 19395 19125
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 20530 19116 20536 19168
rect 20588 19156 20594 19168
rect 20717 19159 20775 19165
rect 20717 19156 20729 19159
rect 20588 19128 20729 19156
rect 20588 19116 20594 19128
rect 20717 19125 20729 19128
rect 20763 19125 20775 19159
rect 20717 19119 20775 19125
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2041 18955 2099 18961
rect 2041 18952 2053 18955
rect 2004 18924 2053 18952
rect 2004 18912 2010 18924
rect 2041 18921 2053 18924
rect 2087 18921 2099 18955
rect 2041 18915 2099 18921
rect 2593 18955 2651 18961
rect 2593 18921 2605 18955
rect 2639 18952 2651 18955
rect 2958 18952 2964 18964
rect 2639 18924 2964 18952
rect 2639 18921 2651 18924
rect 2593 18915 2651 18921
rect 2958 18912 2964 18924
rect 3016 18912 3022 18964
rect 3050 18912 3056 18964
rect 3108 18952 3114 18964
rect 3145 18955 3203 18961
rect 3145 18952 3157 18955
rect 3108 18924 3157 18952
rect 3108 18912 3114 18924
rect 3145 18921 3157 18924
rect 3191 18921 3203 18955
rect 3145 18915 3203 18921
rect 3602 18912 3608 18964
rect 3660 18952 3666 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 3660 18924 8125 18952
rect 3660 18912 3666 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 9030 18952 9036 18964
rect 8260 18924 9036 18952
rect 8260 18912 8266 18924
rect 9030 18912 9036 18924
rect 9088 18912 9094 18964
rect 10778 18952 10784 18964
rect 9600 18924 10784 18952
rect 1026 18844 1032 18896
rect 1084 18884 1090 18896
rect 1084 18856 2636 18884
rect 1084 18844 1090 18856
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18785 1915 18819
rect 1857 18779 1915 18785
rect 1872 18748 1900 18779
rect 2038 18776 2044 18828
rect 2096 18816 2102 18828
rect 2409 18819 2467 18825
rect 2409 18816 2421 18819
rect 2096 18788 2421 18816
rect 2096 18776 2102 18788
rect 2409 18785 2421 18788
rect 2455 18785 2467 18819
rect 2409 18779 2467 18785
rect 2130 18748 2136 18760
rect 1872 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 2608 18748 2636 18856
rect 2682 18844 2688 18896
rect 2740 18884 2746 18896
rect 6816 18887 6874 18893
rect 2740 18856 6776 18884
rect 2740 18844 2746 18856
rect 2961 18819 3019 18825
rect 2961 18785 2973 18819
rect 3007 18816 3019 18819
rect 3234 18816 3240 18828
rect 3007 18788 3240 18816
rect 3007 18785 3019 18788
rect 2961 18779 3019 18785
rect 3234 18776 3240 18788
rect 3292 18776 3298 18828
rect 3786 18776 3792 18828
rect 3844 18816 3850 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 3844 18788 4077 18816
rect 3844 18776 3850 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 6748 18816 6776 18856
rect 6816 18853 6828 18887
rect 6862 18884 6874 18887
rect 6914 18884 6920 18896
rect 6862 18856 6920 18884
rect 6862 18853 6874 18856
rect 6816 18847 6874 18853
rect 6914 18844 6920 18856
rect 6972 18884 6978 18896
rect 6972 18856 8984 18884
rect 6972 18844 6978 18856
rect 8386 18816 8392 18828
rect 4065 18779 4123 18785
rect 4172 18788 4384 18816
rect 6748 18788 8392 18816
rect 4172 18748 4200 18788
rect 2608 18720 4200 18748
rect 4356 18748 4384 18788
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18816 8631 18819
rect 8846 18816 8852 18828
rect 8619 18788 8852 18816
rect 8619 18785 8631 18788
rect 8573 18779 8631 18785
rect 8846 18776 8852 18788
rect 8904 18776 8910 18828
rect 4356 18720 6500 18748
rect 4249 18683 4307 18689
rect 4249 18649 4261 18683
rect 4295 18680 4307 18683
rect 5350 18680 5356 18692
rect 4295 18652 5356 18680
rect 4295 18649 4307 18652
rect 4249 18643 4307 18649
rect 5350 18640 5356 18652
rect 5408 18640 5414 18692
rect 3142 18572 3148 18624
rect 3200 18612 3206 18624
rect 5442 18612 5448 18624
rect 3200 18584 5448 18612
rect 3200 18572 3206 18584
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 6472 18612 6500 18720
rect 6546 18708 6552 18760
rect 6604 18748 6610 18760
rect 6604 18720 6649 18748
rect 6604 18708 6610 18720
rect 7558 18708 7564 18760
rect 7616 18708 7622 18760
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18748 8171 18751
rect 8294 18748 8300 18760
rect 8159 18720 8300 18748
rect 8159 18717 8171 18720
rect 8113 18711 8171 18717
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 8662 18748 8668 18760
rect 8623 18720 8668 18748
rect 8662 18708 8668 18720
rect 8720 18708 8726 18760
rect 8757 18751 8815 18757
rect 8757 18717 8769 18751
rect 8803 18748 8815 18751
rect 8956 18748 8984 18856
rect 8803 18720 8984 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 7576 18680 7604 18708
rect 7576 18652 8340 18680
rect 7558 18612 7564 18624
rect 6472 18584 7564 18612
rect 7558 18572 7564 18584
rect 7616 18572 7622 18624
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 7929 18615 7987 18621
rect 7929 18612 7941 18615
rect 7800 18584 7941 18612
rect 7800 18572 7806 18584
rect 7929 18581 7941 18584
rect 7975 18581 7987 18615
rect 8202 18612 8208 18624
rect 8163 18584 8208 18612
rect 7929 18575 7987 18581
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 8312 18612 8340 18652
rect 8386 18640 8392 18692
rect 8444 18680 8450 18692
rect 9600 18680 9628 18924
rect 10778 18912 10784 18924
rect 10836 18912 10842 18964
rect 10962 18912 10968 18964
rect 11020 18952 11026 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 11020 18924 11069 18952
rect 11020 18912 11026 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 11057 18915 11115 18921
rect 11514 18912 11520 18964
rect 11572 18952 11578 18964
rect 12710 18952 12716 18964
rect 11572 18924 12716 18952
rect 11572 18912 11578 18924
rect 12710 18912 12716 18924
rect 12768 18912 12774 18964
rect 13081 18955 13139 18961
rect 13081 18921 13093 18955
rect 13127 18952 13139 18955
rect 13170 18952 13176 18964
rect 13127 18924 13176 18952
rect 13127 18921 13139 18924
rect 13081 18915 13139 18921
rect 13170 18912 13176 18924
rect 13228 18912 13234 18964
rect 15749 18955 15807 18961
rect 15749 18921 15761 18955
rect 15795 18952 15807 18955
rect 17402 18952 17408 18964
rect 15795 18924 17408 18952
rect 15795 18921 15807 18924
rect 15749 18915 15807 18921
rect 17402 18912 17408 18924
rect 17460 18912 17466 18964
rect 17494 18912 17500 18964
rect 17552 18952 17558 18964
rect 17773 18955 17831 18961
rect 17773 18952 17785 18955
rect 17552 18924 17785 18952
rect 17552 18912 17558 18924
rect 17773 18921 17785 18924
rect 17819 18921 17831 18955
rect 17773 18915 17831 18921
rect 18785 18955 18843 18961
rect 18785 18921 18797 18955
rect 18831 18952 18843 18955
rect 20257 18955 20315 18961
rect 20257 18952 20269 18955
rect 18831 18924 20269 18952
rect 18831 18921 18843 18924
rect 18785 18915 18843 18921
rect 20257 18921 20269 18924
rect 20303 18921 20315 18955
rect 20257 18915 20315 18921
rect 9944 18887 10002 18893
rect 9944 18853 9956 18887
rect 9990 18884 10002 18887
rect 10042 18884 10048 18896
rect 9990 18856 10048 18884
rect 9990 18853 10002 18856
rect 9944 18847 10002 18853
rect 10042 18844 10048 18856
rect 10100 18884 10106 18896
rect 10318 18884 10324 18896
rect 10100 18856 10324 18884
rect 10100 18844 10106 18856
rect 10318 18844 10324 18856
rect 10376 18844 10382 18896
rect 11974 18893 11980 18896
rect 11968 18884 11980 18893
rect 11935 18856 11980 18884
rect 11968 18847 11980 18856
rect 11974 18844 11980 18847
rect 12032 18844 12038 18896
rect 13188 18884 13216 18912
rect 13602 18887 13660 18893
rect 13602 18884 13614 18887
rect 13188 18856 13614 18884
rect 13602 18853 13614 18856
rect 13648 18853 13660 18887
rect 15562 18884 15568 18896
rect 13602 18847 13660 18853
rect 13740 18856 15568 18884
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 9732 18788 9777 18816
rect 9732 18776 9738 18788
rect 10410 18776 10416 18828
rect 10468 18816 10474 18828
rect 13740 18816 13768 18856
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 16942 18844 16948 18896
rect 17000 18884 17006 18896
rect 17000 18856 17540 18884
rect 17000 18844 17006 18856
rect 10468 18788 13768 18816
rect 10468 18776 10474 18788
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 15657 18819 15715 18825
rect 15657 18816 15669 18819
rect 14240 18788 15669 18816
rect 14240 18776 14246 18788
rect 15657 18785 15669 18788
rect 15703 18785 15715 18819
rect 15657 18779 15715 18785
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 16393 18819 16451 18825
rect 16393 18816 16405 18819
rect 15804 18788 16405 18816
rect 15804 18776 15810 18788
rect 16393 18785 16405 18788
rect 16439 18785 16451 18819
rect 16393 18779 16451 18785
rect 16660 18819 16718 18825
rect 16660 18785 16672 18819
rect 16706 18816 16718 18819
rect 17034 18816 17040 18828
rect 16706 18788 17040 18816
rect 16706 18785 16718 18788
rect 16660 18779 16718 18785
rect 17034 18776 17040 18788
rect 17092 18776 17098 18828
rect 17512 18816 17540 18856
rect 17954 18844 17960 18896
rect 18012 18884 18018 18896
rect 18325 18887 18383 18893
rect 18325 18884 18337 18887
rect 18012 18856 18337 18884
rect 18012 18844 18018 18856
rect 18325 18853 18337 18856
rect 18371 18853 18383 18887
rect 18325 18847 18383 18853
rect 18690 18844 18696 18896
rect 18748 18884 18754 18896
rect 19245 18887 19303 18893
rect 19245 18884 19257 18887
rect 18748 18856 19257 18884
rect 18748 18844 18754 18856
rect 19245 18853 19257 18856
rect 19291 18853 19303 18887
rect 19245 18847 19303 18853
rect 18049 18819 18107 18825
rect 18049 18816 18061 18819
rect 17512 18788 18061 18816
rect 18049 18785 18061 18788
rect 18095 18785 18107 18819
rect 18049 18779 18107 18785
rect 18966 18776 18972 18828
rect 19024 18816 19030 18828
rect 19153 18819 19211 18825
rect 19153 18816 19165 18819
rect 19024 18788 19165 18816
rect 19024 18776 19030 18788
rect 19153 18785 19165 18788
rect 19199 18785 19211 18819
rect 19153 18779 19211 18785
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20165 18819 20223 18825
rect 20165 18816 20177 18819
rect 19760 18788 20177 18816
rect 19760 18776 19766 18788
rect 20165 18785 20177 18788
rect 20211 18785 20223 18819
rect 20165 18779 20223 18785
rect 11514 18708 11520 18760
rect 11572 18748 11578 18760
rect 11701 18751 11759 18757
rect 11701 18748 11713 18751
rect 11572 18720 11713 18748
rect 11572 18708 11578 18720
rect 11701 18717 11713 18720
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 12710 18708 12716 18760
rect 12768 18748 12774 18760
rect 13170 18748 13176 18760
rect 12768 18720 13176 18748
rect 12768 18708 12774 18720
rect 13170 18708 13176 18720
rect 13228 18748 13234 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 13228 18720 13369 18748
rect 13228 18708 13234 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18717 15899 18751
rect 19334 18748 19340 18760
rect 19295 18720 19340 18748
rect 15841 18711 15899 18717
rect 14734 18680 14740 18692
rect 8444 18652 9628 18680
rect 14647 18652 14740 18680
rect 8444 18640 8450 18652
rect 14734 18640 14740 18652
rect 14792 18680 14798 18692
rect 15856 18680 15884 18711
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 20349 18751 20407 18757
rect 20349 18748 20361 18751
rect 20036 18720 20361 18748
rect 20036 18708 20042 18720
rect 20349 18717 20361 18720
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20772 18720 20913 18748
rect 20772 18708 20778 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 14792 18652 15884 18680
rect 14792 18640 14798 18652
rect 18782 18640 18788 18692
rect 18840 18680 18846 18692
rect 19797 18683 19855 18689
rect 19797 18680 19809 18683
rect 18840 18652 19809 18680
rect 18840 18640 18846 18652
rect 19797 18649 19809 18652
rect 19843 18649 19855 18683
rect 19797 18643 19855 18649
rect 9582 18612 9588 18624
rect 8312 18584 9588 18612
rect 9582 18572 9588 18584
rect 9640 18572 9646 18624
rect 9858 18572 9864 18624
rect 9916 18612 9922 18624
rect 14458 18612 14464 18624
rect 9916 18584 14464 18612
rect 9916 18572 9922 18584
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 15289 18615 15347 18621
rect 15289 18581 15301 18615
rect 15335 18612 15347 18615
rect 15654 18612 15660 18624
rect 15335 18584 15660 18612
rect 15335 18581 15347 18584
rect 15289 18575 15347 18581
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 2774 18408 2780 18420
rect 2547 18380 2780 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 3510 18408 3516 18420
rect 2976 18380 3516 18408
rect 2222 18300 2228 18352
rect 2280 18340 2286 18352
rect 2976 18340 3004 18380
rect 3510 18368 3516 18380
rect 3568 18368 3574 18420
rect 8662 18408 8668 18420
rect 5920 18380 8668 18408
rect 2280 18312 3004 18340
rect 3053 18343 3111 18349
rect 2280 18300 2286 18312
rect 3053 18309 3065 18343
rect 3099 18340 3111 18343
rect 3970 18340 3976 18352
rect 3099 18312 3976 18340
rect 3099 18309 3111 18312
rect 3053 18303 3111 18309
rect 3970 18300 3976 18312
rect 4028 18300 4034 18352
rect 1854 18232 1860 18284
rect 1912 18272 1918 18284
rect 5920 18272 5948 18380
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 9122 18368 9128 18420
rect 9180 18408 9186 18420
rect 9493 18411 9551 18417
rect 9493 18408 9505 18411
rect 9180 18380 9505 18408
rect 9180 18368 9186 18380
rect 9493 18377 9505 18380
rect 9539 18377 9551 18411
rect 9493 18371 9551 18377
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 10410 18408 10416 18420
rect 9640 18380 10416 18408
rect 9640 18368 9646 18380
rect 10410 18368 10416 18380
rect 10468 18368 10474 18420
rect 11146 18368 11152 18420
rect 11204 18408 11210 18420
rect 11698 18408 11704 18420
rect 11204 18380 11704 18408
rect 11204 18368 11210 18380
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 12529 18411 12587 18417
rect 12529 18377 12541 18411
rect 12575 18408 12587 18411
rect 12986 18408 12992 18420
rect 12575 18380 12992 18408
rect 12575 18377 12587 18380
rect 12529 18371 12587 18377
rect 12986 18368 12992 18380
rect 13044 18368 13050 18420
rect 13170 18368 13176 18420
rect 13228 18368 13234 18420
rect 13725 18411 13783 18417
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 15010 18408 15016 18420
rect 13771 18380 15016 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 15010 18368 15016 18380
rect 15068 18368 15074 18420
rect 15396 18380 16988 18408
rect 8570 18300 8576 18352
rect 8628 18340 8634 18352
rect 10870 18340 10876 18352
rect 8628 18312 10876 18340
rect 8628 18300 8634 18312
rect 10870 18300 10876 18312
rect 10928 18300 10934 18352
rect 11057 18343 11115 18349
rect 11057 18309 11069 18343
rect 11103 18340 11115 18343
rect 12710 18340 12716 18352
rect 11103 18312 12716 18340
rect 11103 18309 11115 18312
rect 11057 18303 11115 18309
rect 12710 18300 12716 18312
rect 12768 18300 12774 18352
rect 12894 18300 12900 18352
rect 12952 18340 12958 18352
rect 13188 18340 13216 18368
rect 12952 18312 14136 18340
rect 12952 18300 12958 18312
rect 6086 18272 6092 18284
rect 1912 18244 5948 18272
rect 6047 18244 6092 18272
rect 1912 18232 1918 18244
rect 6086 18232 6092 18244
rect 6144 18232 6150 18284
rect 6546 18232 6552 18284
rect 6604 18272 6610 18284
rect 6825 18275 6883 18281
rect 6825 18272 6837 18275
rect 6604 18244 6837 18272
rect 6604 18232 6610 18244
rect 6825 18241 6837 18244
rect 6871 18241 6883 18275
rect 8478 18272 8484 18284
rect 8439 18244 8484 18272
rect 6825 18235 6883 18241
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2314 18204 2320 18216
rect 2275 18176 2320 18204
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 2958 18204 2964 18216
rect 2915 18176 2964 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 2958 18164 2964 18176
rect 3016 18164 3022 18216
rect 3421 18207 3479 18213
rect 3421 18173 3433 18207
rect 3467 18204 3479 18207
rect 3878 18204 3884 18216
rect 3467 18176 3884 18204
rect 3467 18173 3479 18176
rect 3421 18167 3479 18173
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 5905 18207 5963 18213
rect 5905 18173 5917 18207
rect 5951 18204 5963 18207
rect 6730 18204 6736 18216
rect 5951 18176 6736 18204
rect 5951 18173 5963 18176
rect 5905 18167 5963 18173
rect 6730 18164 6736 18176
rect 6788 18164 6794 18216
rect 4798 18096 4804 18148
rect 4856 18136 4862 18148
rect 5350 18136 5356 18148
rect 4856 18108 5356 18136
rect 4856 18096 4862 18108
rect 5350 18096 5356 18108
rect 5408 18096 5414 18148
rect 1394 18028 1400 18080
rect 1452 18068 1458 18080
rect 2866 18068 2872 18080
rect 1452 18040 2872 18068
rect 1452 18028 1458 18040
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 3602 18068 3608 18080
rect 3563 18040 3608 18068
rect 3602 18028 3608 18040
rect 3660 18028 3666 18080
rect 5902 18028 5908 18080
rect 5960 18068 5966 18080
rect 6840 18068 6868 18235
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 10042 18272 10048 18284
rect 10003 18244 10048 18272
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 10134 18232 10140 18284
rect 10192 18272 10198 18284
rect 10505 18275 10563 18281
rect 10505 18272 10517 18275
rect 10192 18244 10517 18272
rect 10192 18232 10198 18244
rect 10505 18241 10517 18244
rect 10551 18241 10563 18275
rect 10505 18235 10563 18241
rect 11609 18275 11667 18281
rect 11609 18241 11621 18275
rect 11655 18241 11667 18275
rect 11609 18235 11667 18241
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 13262 18272 13268 18284
rect 13219 18244 13268 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 7092 18207 7150 18213
rect 7092 18173 7104 18207
rect 7138 18204 7150 18207
rect 11624 18204 11652 18235
rect 13262 18232 13268 18244
rect 13320 18232 13326 18284
rect 14108 18281 14136 18312
rect 14093 18275 14151 18281
rect 14093 18241 14105 18275
rect 14139 18241 14151 18275
rect 14093 18235 14151 18241
rect 11790 18204 11796 18216
rect 7138 18176 11796 18204
rect 7138 18173 7150 18176
rect 7092 18167 7150 18173
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 11974 18164 11980 18216
rect 12032 18204 12038 18216
rect 13541 18207 13599 18213
rect 13541 18204 13553 18207
rect 12032 18176 13553 18204
rect 12032 18164 12038 18176
rect 13541 18173 13553 18176
rect 13587 18173 13599 18207
rect 13541 18167 13599 18173
rect 14360 18207 14418 18213
rect 14360 18173 14372 18207
rect 14406 18204 14418 18207
rect 14734 18204 14740 18216
rect 14406 18176 14740 18204
rect 14406 18173 14418 18176
rect 14360 18167 14418 18173
rect 14734 18164 14740 18176
rect 14792 18204 14798 18216
rect 14792 18176 15056 18204
rect 14792 18164 14798 18176
rect 15028 18148 15056 18176
rect 9214 18096 9220 18148
rect 9272 18136 9278 18148
rect 10594 18136 10600 18148
rect 9272 18108 10600 18136
rect 9272 18096 9278 18108
rect 10594 18096 10600 18108
rect 10652 18096 10658 18148
rect 11146 18096 11152 18148
rect 11204 18136 11210 18148
rect 11517 18139 11575 18145
rect 11517 18136 11529 18139
rect 11204 18108 11529 18136
rect 11204 18096 11210 18108
rect 11517 18105 11529 18108
rect 11563 18105 11575 18139
rect 11517 18099 11575 18105
rect 12897 18139 12955 18145
rect 12897 18105 12909 18139
rect 12943 18136 12955 18139
rect 13078 18136 13084 18148
rect 12943 18108 13084 18136
rect 12943 18105 12955 18108
rect 12897 18099 12955 18105
rect 13078 18096 13084 18108
rect 13136 18096 13142 18148
rect 13170 18096 13176 18148
rect 13228 18136 13234 18148
rect 13630 18136 13636 18148
rect 13228 18108 13636 18136
rect 13228 18096 13234 18108
rect 13630 18096 13636 18108
rect 13688 18096 13694 18148
rect 15010 18096 15016 18148
rect 15068 18096 15074 18148
rect 5960 18040 6868 18068
rect 5960 18028 5966 18040
rect 6914 18028 6920 18080
rect 6972 18068 6978 18080
rect 8205 18071 8263 18077
rect 8205 18068 8217 18071
rect 6972 18040 8217 18068
rect 6972 18028 6978 18040
rect 8205 18037 8217 18040
rect 8251 18037 8263 18071
rect 8205 18031 8263 18037
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 9306 18068 9312 18080
rect 8352 18040 9312 18068
rect 8352 18028 8358 18040
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 9861 18071 9919 18077
rect 9861 18068 9873 18071
rect 9824 18040 9873 18068
rect 9824 18028 9830 18040
rect 9861 18037 9873 18040
rect 9907 18037 9919 18071
rect 9861 18031 9919 18037
rect 9953 18071 10011 18077
rect 9953 18037 9965 18071
rect 9999 18068 10011 18071
rect 10042 18068 10048 18080
rect 9999 18040 10048 18068
rect 9999 18037 10011 18040
rect 9953 18031 10011 18037
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 11422 18068 11428 18080
rect 11383 18040 11428 18068
rect 11422 18028 11428 18040
rect 11480 18028 11486 18080
rect 12986 18068 12992 18080
rect 12947 18040 12992 18068
rect 12986 18028 12992 18040
rect 13044 18068 13050 18080
rect 15396 18068 15424 18380
rect 16960 18340 16988 18380
rect 17034 18368 17040 18420
rect 17092 18408 17098 18420
rect 17129 18411 17187 18417
rect 17129 18408 17141 18411
rect 17092 18380 17141 18408
rect 17092 18368 17098 18380
rect 17129 18377 17141 18380
rect 17175 18377 17187 18411
rect 17129 18371 17187 18377
rect 17589 18411 17647 18417
rect 17589 18377 17601 18411
rect 17635 18408 17647 18411
rect 17770 18408 17776 18420
rect 17635 18380 17776 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 19518 18408 19524 18420
rect 17880 18380 19524 18408
rect 17880 18340 17908 18380
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 19702 18408 19708 18420
rect 19663 18380 19708 18408
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 16960 18312 17908 18340
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 20257 18275 20315 18281
rect 20257 18272 20269 18275
rect 19300 18244 20269 18272
rect 19300 18232 19306 18244
rect 20257 18241 20269 18244
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 15746 18204 15752 18216
rect 15707 18176 15752 18204
rect 15746 18164 15752 18176
rect 15804 18164 15810 18216
rect 16298 18164 16304 18216
rect 16356 18204 16362 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 16356 18176 17417 18204
rect 16356 18164 16362 18176
rect 17405 18173 17417 18176
rect 17451 18204 17463 18207
rect 17954 18204 17960 18216
rect 17451 18176 17960 18204
rect 17451 18173 17463 18176
rect 17405 18167 17463 18173
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 18598 18204 18604 18216
rect 18095 18176 18604 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 18782 18164 18788 18216
rect 18840 18204 18846 18216
rect 20165 18207 20223 18213
rect 20165 18204 20177 18207
rect 18840 18176 20177 18204
rect 18840 18164 18846 18176
rect 20165 18173 20177 18176
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 20717 18207 20775 18213
rect 20717 18173 20729 18207
rect 20763 18204 20775 18207
rect 20990 18204 20996 18216
rect 20763 18176 20996 18204
rect 20763 18173 20775 18176
rect 20717 18167 20775 18173
rect 20990 18164 20996 18176
rect 21048 18164 21054 18216
rect 15838 18136 15844 18148
rect 15488 18108 15844 18136
rect 15488 18077 15516 18108
rect 15838 18096 15844 18108
rect 15896 18136 15902 18148
rect 15994 18139 16052 18145
rect 15994 18136 16006 18139
rect 15896 18108 16006 18136
rect 15896 18096 15902 18108
rect 15994 18105 16006 18108
rect 16040 18105 16052 18139
rect 15994 18099 16052 18105
rect 17494 18096 17500 18148
rect 17552 18136 17558 18148
rect 18294 18139 18352 18145
rect 18294 18136 18306 18139
rect 17552 18108 18306 18136
rect 17552 18096 17558 18108
rect 18294 18105 18306 18108
rect 18340 18105 18352 18139
rect 18294 18099 18352 18105
rect 20073 18139 20131 18145
rect 20073 18105 20085 18139
rect 20119 18136 20131 18139
rect 20806 18136 20812 18148
rect 20119 18108 20812 18136
rect 20119 18105 20131 18108
rect 20073 18099 20131 18105
rect 20806 18096 20812 18108
rect 20864 18096 20870 18148
rect 13044 18040 15424 18068
rect 15473 18071 15531 18077
rect 13044 18028 13050 18040
rect 15473 18037 15485 18071
rect 15519 18037 15531 18071
rect 15473 18031 15531 18037
rect 19242 18028 19248 18080
rect 19300 18068 19306 18080
rect 19429 18071 19487 18077
rect 19429 18068 19441 18071
rect 19300 18040 19441 18068
rect 19300 18028 19306 18040
rect 19429 18037 19441 18040
rect 19475 18037 19487 18071
rect 19429 18031 19487 18037
rect 20622 18028 20628 18080
rect 20680 18068 20686 18080
rect 20901 18071 20959 18077
rect 20901 18068 20913 18071
rect 20680 18040 20913 18068
rect 20680 18028 20686 18040
rect 20901 18037 20913 18040
rect 20947 18037 20959 18071
rect 20901 18031 20959 18037
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 6917 17867 6975 17873
rect 6917 17864 6929 17867
rect 3568 17836 6929 17864
rect 3568 17824 3574 17836
rect 6917 17833 6929 17836
rect 6963 17833 6975 17867
rect 6917 17827 6975 17833
rect 7006 17824 7012 17876
rect 7064 17864 7070 17876
rect 7101 17867 7159 17873
rect 7101 17864 7113 17867
rect 7064 17836 7113 17864
rect 7064 17824 7070 17836
rect 7101 17833 7113 17836
rect 7147 17833 7159 17867
rect 7466 17864 7472 17876
rect 7427 17836 7472 17864
rect 7101 17827 7159 17833
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 7561 17867 7619 17873
rect 7561 17833 7573 17867
rect 7607 17864 7619 17867
rect 8202 17864 8208 17876
rect 7607 17836 8208 17864
rect 7607 17833 7619 17836
rect 7561 17827 7619 17833
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 8573 17867 8631 17873
rect 8573 17864 8585 17867
rect 8444 17836 8585 17864
rect 8444 17824 8450 17836
rect 8573 17833 8585 17836
rect 8619 17833 8631 17867
rect 9858 17864 9864 17876
rect 9819 17836 9864 17864
rect 8573 17827 8631 17833
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 11422 17824 11428 17876
rect 11480 17864 11486 17876
rect 12069 17867 12127 17873
rect 12069 17864 12081 17867
rect 11480 17836 12081 17864
rect 11480 17824 11486 17836
rect 12069 17833 12081 17836
rect 12115 17833 12127 17867
rect 12069 17827 12127 17833
rect 12529 17867 12587 17873
rect 12529 17833 12541 17867
rect 12575 17864 12587 17867
rect 13262 17864 13268 17876
rect 12575 17836 13268 17864
rect 12575 17833 12587 17836
rect 12529 17827 12587 17833
rect 13262 17824 13268 17836
rect 13320 17864 13326 17876
rect 14550 17864 14556 17876
rect 13320 17836 14556 17864
rect 13320 17824 13326 17836
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15654 17864 15660 17876
rect 15615 17836 15660 17864
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 16485 17867 16543 17873
rect 16485 17833 16497 17867
rect 16531 17864 16543 17867
rect 16758 17864 16764 17876
rect 16531 17836 16764 17864
rect 16531 17833 16543 17836
rect 16485 17827 16543 17833
rect 16758 17824 16764 17836
rect 16816 17824 16822 17876
rect 16853 17867 16911 17873
rect 16853 17833 16865 17867
rect 16899 17864 16911 17867
rect 16942 17864 16948 17876
rect 16899 17836 16948 17864
rect 16899 17833 16911 17836
rect 16853 17827 16911 17833
rect 16942 17824 16948 17836
rect 17000 17824 17006 17876
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 17497 17867 17555 17873
rect 17497 17864 17509 17867
rect 17276 17836 17509 17864
rect 17276 17824 17282 17836
rect 17497 17833 17509 17836
rect 17543 17833 17555 17867
rect 17497 17827 17555 17833
rect 17865 17867 17923 17873
rect 17865 17833 17877 17867
rect 17911 17864 17923 17867
rect 20714 17864 20720 17876
rect 17911 17836 20720 17864
rect 17911 17833 17923 17836
rect 17865 17827 17923 17833
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 20806 17824 20812 17876
rect 20864 17864 20870 17876
rect 20901 17867 20959 17873
rect 20901 17864 20913 17867
rect 20864 17836 20913 17864
rect 20864 17824 20870 17836
rect 20901 17833 20913 17836
rect 20947 17833 20959 17867
rect 20901 17827 20959 17833
rect 2314 17756 2320 17808
rect 2372 17796 2378 17808
rect 2501 17799 2559 17805
rect 2501 17796 2513 17799
rect 2372 17768 2513 17796
rect 2372 17756 2378 17768
rect 2501 17765 2513 17768
rect 2547 17765 2559 17799
rect 2501 17759 2559 17765
rect 9582 17756 9588 17808
rect 9640 17796 9646 17808
rect 18868 17799 18926 17805
rect 9640 17768 18644 17796
rect 9640 17756 9646 17768
rect 1670 17728 1676 17740
rect 1631 17700 1676 17728
rect 1670 17688 1676 17700
rect 1728 17688 1734 17740
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17697 2283 17731
rect 2225 17691 2283 17697
rect 2130 17660 2136 17672
rect 1872 17632 2136 17660
rect 1872 17601 1900 17632
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 2240 17660 2268 17691
rect 3326 17688 3332 17740
rect 3384 17728 3390 17740
rect 3881 17731 3939 17737
rect 3881 17728 3893 17731
rect 3384 17700 3893 17728
rect 3384 17688 3390 17700
rect 3881 17697 3893 17700
rect 3927 17697 3939 17731
rect 5074 17728 5080 17740
rect 5035 17700 5080 17728
rect 3881 17691 3939 17697
rect 5074 17688 5080 17700
rect 5132 17688 5138 17740
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17728 5411 17731
rect 5813 17731 5871 17737
rect 5813 17728 5825 17731
rect 5399 17700 5825 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 5813 17697 5825 17700
rect 5859 17697 5871 17731
rect 5813 17691 5871 17697
rect 6917 17731 6975 17737
rect 6917 17697 6929 17731
rect 6963 17728 6975 17731
rect 6963 17700 8432 17728
rect 6963 17697 6975 17700
rect 6917 17691 6975 17697
rect 7006 17660 7012 17672
rect 2240 17632 7012 17660
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 7742 17660 7748 17672
rect 7703 17632 7748 17660
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 8404 17660 8432 17700
rect 8478 17688 8484 17740
rect 8536 17728 8542 17740
rect 8536 17700 8581 17728
rect 8680 17700 9076 17728
rect 8536 17688 8542 17700
rect 8680 17660 8708 17700
rect 8404 17632 8708 17660
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17660 8815 17663
rect 8938 17660 8944 17672
rect 8803 17632 8944 17660
rect 8803 17629 8815 17632
rect 8757 17623 8815 17629
rect 8938 17620 8944 17632
rect 8996 17620 9002 17672
rect 9048 17660 9076 17700
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9180 17700 9689 17728
rect 9180 17688 9186 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 10226 17688 10232 17740
rect 10284 17728 10290 17740
rect 10413 17731 10471 17737
rect 10413 17728 10425 17731
rect 10284 17700 10425 17728
rect 10284 17688 10290 17700
rect 10413 17697 10425 17700
rect 10459 17697 10471 17731
rect 10413 17691 10471 17697
rect 10680 17731 10738 17737
rect 10680 17697 10692 17731
rect 10726 17728 10738 17731
rect 10962 17728 10968 17740
rect 10726 17700 10968 17728
rect 10726 17697 10738 17700
rect 10680 17691 10738 17697
rect 10962 17688 10968 17700
rect 11020 17688 11026 17740
rect 11882 17688 11888 17740
rect 11940 17728 11946 17740
rect 12437 17731 12495 17737
rect 12437 17728 12449 17731
rect 11940 17700 12449 17728
rect 11940 17688 11946 17700
rect 12437 17697 12449 17700
rect 12483 17697 12495 17731
rect 12437 17691 12495 17697
rect 12710 17688 12716 17740
rect 12768 17728 12774 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 12768 17700 13093 17728
rect 12768 17688 12774 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 14553 17731 14611 17737
rect 14553 17697 14565 17731
rect 14599 17728 14611 17731
rect 14918 17728 14924 17740
rect 14599 17700 14924 17728
rect 14599 17697 14611 17700
rect 14553 17691 14611 17697
rect 14918 17688 14924 17700
rect 14976 17688 14982 17740
rect 15749 17731 15807 17737
rect 15749 17728 15761 17731
rect 15120 17700 15761 17728
rect 10042 17660 10048 17672
rect 9048 17632 10048 17660
rect 10042 17620 10048 17632
rect 10100 17660 10106 17672
rect 10318 17660 10324 17672
rect 10100 17632 10324 17660
rect 10100 17620 10106 17632
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 12618 17660 12624 17672
rect 12579 17632 12624 17660
rect 12618 17620 12624 17632
rect 12676 17620 12682 17672
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17629 13323 17663
rect 13265 17623 13323 17629
rect 1857 17595 1915 17601
rect 1857 17561 1869 17595
rect 1903 17561 1915 17595
rect 1857 17555 1915 17561
rect 3881 17595 3939 17601
rect 3881 17561 3893 17595
rect 3927 17592 3939 17595
rect 5810 17592 5816 17604
rect 3927 17564 5816 17592
rect 3927 17561 3939 17564
rect 3881 17555 3939 17561
rect 5810 17552 5816 17564
rect 5868 17552 5874 17604
rect 5997 17595 6055 17601
rect 5997 17561 6009 17595
rect 6043 17592 6055 17595
rect 6043 17564 9260 17592
rect 6043 17561 6055 17564
rect 5997 17555 6055 17561
rect 1762 17484 1768 17536
rect 1820 17524 1826 17536
rect 3326 17524 3332 17536
rect 1820 17496 3332 17524
rect 1820 17484 1826 17496
rect 3326 17484 3332 17496
rect 3384 17484 3390 17536
rect 3418 17484 3424 17536
rect 3476 17524 3482 17536
rect 6914 17524 6920 17536
rect 3476 17496 6920 17524
rect 3476 17484 3482 17496
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 7190 17484 7196 17536
rect 7248 17524 7254 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7248 17496 8125 17524
rect 7248 17484 7254 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 9232 17524 9260 17564
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 10226 17592 10232 17604
rect 9364 17564 10232 17592
rect 9364 17552 9370 17564
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 11790 17592 11796 17604
rect 11751 17564 11796 17592
rect 11790 17552 11796 17564
rect 11848 17552 11854 17604
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 13280 17592 13308 17623
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 13688 17632 14657 17660
rect 13688 17620 13694 17632
rect 14645 17629 14657 17632
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17660 14887 17663
rect 15010 17660 15016 17672
rect 14875 17632 15016 17660
rect 14875 17629 14887 17632
rect 14829 17623 14887 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 12216 17564 13308 17592
rect 14185 17595 14243 17601
rect 12216 17552 12222 17564
rect 14185 17561 14197 17595
rect 14231 17592 14243 17595
rect 15120 17592 15148 17700
rect 15749 17697 15761 17700
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 17184 17700 17969 17728
rect 17184 17688 17190 17700
rect 17957 17697 17969 17700
rect 18003 17728 18015 17731
rect 18506 17728 18512 17740
rect 18003 17700 18512 17728
rect 18003 17697 18015 17700
rect 17957 17691 18015 17697
rect 18506 17688 18512 17700
rect 18564 17688 18570 17740
rect 18616 17728 18644 17768
rect 18868 17765 18880 17799
rect 18914 17796 18926 17799
rect 19242 17796 19248 17808
rect 18914 17768 19248 17796
rect 18914 17765 18926 17768
rect 18868 17759 18926 17765
rect 19242 17756 19248 17768
rect 19300 17756 19306 17808
rect 21726 17796 21732 17808
rect 19352 17768 21732 17796
rect 19352 17728 19380 17768
rect 21726 17756 21732 17768
rect 21784 17756 21790 17808
rect 20254 17728 20260 17740
rect 18616 17700 19380 17728
rect 20215 17700 20260 17728
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 15838 17660 15844 17672
rect 15799 17632 15844 17660
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16945 17663 17003 17669
rect 16945 17629 16957 17663
rect 16991 17629 17003 17663
rect 16945 17623 17003 17629
rect 14231 17564 15148 17592
rect 14231 17561 14243 17564
rect 14185 17555 14243 17561
rect 12250 17524 12256 17536
rect 9232 17496 12256 17524
rect 8113 17487 8171 17493
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 13446 17484 13452 17536
rect 13504 17524 13510 17536
rect 16960 17524 16988 17623
rect 17034 17620 17040 17672
rect 17092 17660 17098 17672
rect 18049 17663 18107 17669
rect 17092 17632 17137 17660
rect 17092 17620 17098 17632
rect 18049 17629 18061 17663
rect 18095 17629 18107 17663
rect 18598 17660 18604 17672
rect 18511 17632 18604 17660
rect 18049 17623 18107 17629
rect 17052 17592 17080 17620
rect 18064 17592 18092 17623
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 17052 17564 18092 17592
rect 13504 17496 16988 17524
rect 18616 17524 18644 17620
rect 18782 17524 18788 17536
rect 18616 17496 18788 17524
rect 13504 17484 13510 17496
rect 18782 17484 18788 17496
rect 18840 17484 18846 17536
rect 19794 17484 19800 17536
rect 19852 17524 19858 17536
rect 19978 17524 19984 17536
rect 19852 17496 19984 17524
rect 19852 17484 19858 17496
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 20438 17524 20444 17536
rect 20399 17496 20444 17524
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2774 17320 2780 17332
rect 2547 17292 2780 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3050 17320 3056 17332
rect 3011 17292 3056 17320
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 3142 17280 3148 17332
rect 3200 17320 3206 17332
rect 3605 17323 3663 17329
rect 3605 17320 3617 17323
rect 3200 17292 3617 17320
rect 3200 17280 3206 17292
rect 3605 17289 3617 17292
rect 3651 17289 3663 17323
rect 3605 17283 3663 17289
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 5132 17292 5457 17320
rect 5132 17280 5138 17292
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 5445 17283 5503 17289
rect 5810 17280 5816 17332
rect 5868 17320 5874 17332
rect 8018 17320 8024 17332
rect 5868 17292 8024 17320
rect 5868 17280 5874 17292
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 10778 17320 10784 17332
rect 8128 17292 10784 17320
rect 2866 17212 2872 17264
rect 2924 17252 2930 17264
rect 8128 17252 8156 17292
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 10873 17323 10931 17329
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 11146 17320 11152 17332
rect 10919 17292 11152 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 12618 17320 12624 17332
rect 11532 17292 12624 17320
rect 2924 17224 8156 17252
rect 8312 17224 9812 17252
rect 2924 17212 2930 17224
rect 4706 17144 4712 17196
rect 4764 17184 4770 17196
rect 4985 17187 5043 17193
rect 4985 17184 4997 17187
rect 4764 17156 4997 17184
rect 4764 17144 4770 17156
rect 4985 17153 4997 17156
rect 5031 17153 5043 17187
rect 5994 17184 6000 17196
rect 5955 17156 6000 17184
rect 4985 17147 5043 17153
rect 5994 17144 6000 17156
rect 6052 17144 6058 17196
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7466 17184 7472 17196
rect 6972 17156 7328 17184
rect 7427 17156 7472 17184
rect 6972 17144 6978 17156
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 1780 17048 1808 17079
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 1912 17088 2329 17116
rect 1912 17076 1918 17088
rect 2317 17085 2329 17088
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17085 2927 17119
rect 3418 17116 3424 17128
rect 3379 17088 3424 17116
rect 2869 17079 2927 17085
rect 2406 17048 2412 17060
rect 1780 17020 2412 17048
rect 2406 17008 2412 17020
rect 2464 17008 2470 17060
rect 2884 17048 2912 17079
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 6270 17116 6276 17128
rect 3528 17088 6276 17116
rect 3528 17048 3556 17088
rect 6270 17076 6276 17088
rect 6328 17076 6334 17128
rect 7190 17116 7196 17128
rect 7151 17088 7196 17116
rect 7190 17076 7196 17088
rect 7248 17076 7254 17128
rect 7300 17116 7328 17156
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 7558 17144 7564 17196
rect 7616 17184 7622 17196
rect 8312 17193 8340 17224
rect 8297 17187 8355 17193
rect 8297 17184 8309 17187
rect 7616 17156 8309 17184
rect 7616 17144 7622 17156
rect 8297 17153 8309 17156
rect 8343 17153 8355 17187
rect 8297 17147 8355 17153
rect 8481 17187 8539 17193
rect 8481 17153 8493 17187
rect 8527 17184 8539 17187
rect 8938 17184 8944 17196
rect 8527 17156 8944 17184
rect 8527 17153 8539 17156
rect 8481 17147 8539 17153
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 9122 17184 9128 17196
rect 9083 17156 9128 17184
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 8205 17119 8263 17125
rect 7300 17088 8156 17116
rect 5905 17051 5963 17057
rect 5905 17048 5917 17051
rect 2884 17020 3556 17048
rect 4448 17020 5917 17048
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 4448 16989 4476 17020
rect 5905 17017 5917 17020
rect 5951 17017 5963 17051
rect 5905 17011 5963 17017
rect 4433 16983 4491 16989
rect 4433 16949 4445 16983
rect 4479 16949 4491 16983
rect 4798 16980 4804 16992
rect 4759 16952 4804 16980
rect 4433 16943 4491 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 5810 16980 5816 16992
rect 4948 16952 4993 16980
rect 5771 16952 5816 16980
rect 4948 16940 4954 16952
rect 5810 16940 5816 16952
rect 5868 16940 5874 16992
rect 6822 16980 6828 16992
rect 6783 16952 6828 16980
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 7285 16983 7343 16989
rect 7285 16949 7297 16983
rect 7331 16980 7343 16983
rect 7837 16983 7895 16989
rect 7837 16980 7849 16983
rect 7331 16952 7849 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 7837 16949 7849 16952
rect 7883 16949 7895 16983
rect 8128 16980 8156 17088
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 8662 17116 8668 17128
rect 8251 17088 8668 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17116 8907 17119
rect 9674 17116 9680 17128
rect 8895 17088 9680 17116
rect 8895 17085 8907 17088
rect 8849 17079 8907 17085
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 9784 17116 9812 17224
rect 10962 17212 10968 17264
rect 11020 17252 11026 17264
rect 11532 17252 11560 17292
rect 12618 17280 12624 17292
rect 12676 17320 12682 17332
rect 17862 17320 17868 17332
rect 12676 17292 17868 17320
rect 12676 17280 12682 17292
rect 17862 17280 17868 17292
rect 17920 17280 17926 17332
rect 14182 17252 14188 17264
rect 11020 17224 11560 17252
rect 11020 17212 11026 17224
rect 9858 17144 9864 17196
rect 9916 17184 9922 17196
rect 11054 17184 11060 17196
rect 9916 17156 11060 17184
rect 9916 17144 9922 17156
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 11532 17193 11560 17224
rect 12636 17224 14188 17252
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17153 11575 17187
rect 11882 17184 11888 17196
rect 11843 17156 11888 17184
rect 11517 17147 11575 17153
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 12636 17193 12664 17224
rect 14182 17212 14188 17224
rect 14240 17212 14246 17264
rect 14369 17255 14427 17261
rect 14369 17221 14381 17255
rect 14415 17221 14427 17255
rect 14369 17215 14427 17221
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 12860 17156 13553 17184
rect 12860 17144 12866 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13722 17184 13728 17196
rect 13683 17156 13728 17184
rect 13541 17147 13599 17153
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 13446 17116 13452 17128
rect 9784 17088 13308 17116
rect 13407 17088 13452 17116
rect 8294 17008 8300 17060
rect 8352 17048 8358 17060
rect 10962 17048 10968 17060
rect 8352 17020 10968 17048
rect 8352 17008 8358 17020
rect 10962 17008 10968 17020
rect 11020 17008 11026 17060
rect 11333 17051 11391 17057
rect 11333 17048 11345 17051
rect 11072 17020 11345 17048
rect 8570 16980 8576 16992
rect 8128 16952 8576 16980
rect 7837 16943 7895 16949
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 8662 16940 8668 16992
rect 8720 16980 8726 16992
rect 10226 16980 10232 16992
rect 8720 16952 10232 16980
rect 8720 16940 8726 16952
rect 10226 16940 10232 16952
rect 10284 16940 10290 16992
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 11072 16980 11100 17020
rect 11333 17017 11345 17020
rect 11379 17017 11391 17051
rect 11333 17011 11391 17017
rect 11422 17008 11428 17060
rect 11480 17048 11486 17060
rect 13280 17048 13308 17088
rect 13446 17076 13452 17088
rect 13504 17076 13510 17128
rect 14384 17116 14412 17215
rect 14550 17212 14556 17264
rect 14608 17252 14614 17264
rect 14608 17224 16160 17252
rect 14608 17212 14614 17224
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17184 15071 17187
rect 16022 17184 16028 17196
rect 15059 17156 16028 17184
rect 15059 17153 15071 17156
rect 15013 17147 15071 17153
rect 16022 17144 16028 17156
rect 16080 17144 16086 17196
rect 15381 17119 15439 17125
rect 15381 17116 15393 17119
rect 14384 17088 15393 17116
rect 15381 17085 15393 17088
rect 15427 17085 15439 17119
rect 15381 17079 15439 17085
rect 13906 17048 13912 17060
rect 11480 17020 13216 17048
rect 13280 17020 13912 17048
rect 11480 17008 11486 17020
rect 11238 16980 11244 16992
rect 10836 16952 11100 16980
rect 11151 16952 11244 16980
rect 10836 16940 10842 16952
rect 11238 16940 11244 16952
rect 11296 16980 11302 16992
rect 11882 16980 11888 16992
rect 11296 16952 11888 16980
rect 11296 16940 11302 16952
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 13078 16980 13084 16992
rect 13039 16952 13084 16980
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 13188 16980 13216 17020
rect 13906 17008 13912 17020
rect 13964 17008 13970 17060
rect 13998 17008 14004 17060
rect 14056 17048 14062 17060
rect 14829 17051 14887 17057
rect 14829 17048 14841 17051
rect 14056 17020 14841 17048
rect 14056 17008 14062 17020
rect 14829 17017 14841 17020
rect 14875 17017 14887 17051
rect 14829 17011 14887 17017
rect 14918 17008 14924 17060
rect 14976 17008 14982 17060
rect 15194 17008 15200 17060
rect 15252 17048 15258 17060
rect 15657 17051 15715 17057
rect 15657 17048 15669 17051
rect 15252 17020 15669 17048
rect 15252 17008 15258 17020
rect 15657 17017 15669 17020
rect 15703 17017 15715 17051
rect 16132 17048 16160 17224
rect 17494 17212 17500 17264
rect 17552 17252 17558 17264
rect 19150 17252 19156 17264
rect 17552 17224 19156 17252
rect 17552 17212 17558 17224
rect 19150 17212 19156 17224
rect 19208 17252 19214 17264
rect 20990 17252 20996 17264
rect 19208 17224 20996 17252
rect 19208 17212 19214 17224
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 16574 17184 16580 17196
rect 16535 17156 16580 17184
rect 16574 17144 16580 17156
rect 16632 17144 16638 17196
rect 16960 17156 17264 17184
rect 16301 17119 16359 17125
rect 16301 17085 16313 17119
rect 16347 17116 16359 17119
rect 16850 17116 16856 17128
rect 16347 17088 16856 17116
rect 16347 17085 16359 17088
rect 16301 17079 16359 17085
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 16960 17048 16988 17156
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17085 17187 17119
rect 17236 17116 17264 17156
rect 18322 17144 18328 17196
rect 18380 17184 18386 17196
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 18380 17156 18613 17184
rect 18380 17144 18386 17156
rect 18601 17153 18613 17156
rect 18647 17184 18659 17187
rect 18874 17184 18880 17196
rect 18647 17156 18880 17184
rect 18647 17153 18659 17156
rect 18601 17147 18659 17153
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 19242 17144 19248 17196
rect 19300 17184 19306 17196
rect 19613 17187 19671 17193
rect 19613 17184 19625 17187
rect 19300 17156 19625 17184
rect 19300 17144 19306 17156
rect 19613 17153 19625 17156
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 19518 17116 19524 17128
rect 17236 17088 19524 17116
rect 17129 17079 17187 17085
rect 16132 17020 16988 17048
rect 15657 17011 15715 17017
rect 13630 16980 13636 16992
rect 13188 16952 13636 16980
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 14090 16940 14096 16992
rect 14148 16980 14154 16992
rect 14737 16983 14795 16989
rect 14737 16980 14749 16983
rect 14148 16952 14749 16980
rect 14148 16940 14154 16952
rect 14737 16949 14749 16952
rect 14783 16949 14795 16983
rect 14936 16980 14964 17008
rect 15562 16980 15568 16992
rect 14936 16952 15568 16980
rect 14737 16943 14795 16949
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 17144 16980 17172 17079
rect 19518 17076 19524 17088
rect 19576 17076 19582 17128
rect 20530 17116 20536 17128
rect 20491 17088 20536 17116
rect 20530 17076 20536 17088
rect 20588 17076 20594 17128
rect 17218 17008 17224 17060
rect 17276 17048 17282 17060
rect 17405 17051 17463 17057
rect 17405 17048 17417 17051
rect 17276 17020 17417 17048
rect 17276 17008 17282 17020
rect 17405 17017 17417 17020
rect 17451 17017 17463 17051
rect 17405 17011 17463 17017
rect 17954 17008 17960 17060
rect 18012 17048 18018 17060
rect 18417 17051 18475 17057
rect 18417 17048 18429 17051
rect 18012 17020 18429 17048
rect 18012 17008 18018 17020
rect 18417 17017 18429 17020
rect 18463 17017 18475 17051
rect 18417 17011 18475 17017
rect 18049 16983 18107 16989
rect 18049 16980 18061 16983
rect 17144 16952 18061 16980
rect 18049 16949 18061 16952
rect 18095 16949 18107 16983
rect 18049 16943 18107 16949
rect 18509 16983 18567 16989
rect 18509 16949 18521 16983
rect 18555 16980 18567 16983
rect 19061 16983 19119 16989
rect 19061 16980 19073 16983
rect 18555 16952 19073 16980
rect 18555 16949 18567 16952
rect 18509 16943 18567 16949
rect 19061 16949 19073 16952
rect 19107 16949 19119 16983
rect 19061 16943 19119 16949
rect 19150 16940 19156 16992
rect 19208 16980 19214 16992
rect 19429 16983 19487 16989
rect 19429 16980 19441 16983
rect 19208 16952 19441 16980
rect 19208 16940 19214 16952
rect 19429 16949 19441 16952
rect 19475 16949 19487 16983
rect 19429 16943 19487 16949
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 19576 16952 19621 16980
rect 19576 16940 19582 16952
rect 19702 16940 19708 16992
rect 19760 16980 19766 16992
rect 20073 16983 20131 16989
rect 20073 16980 20085 16983
rect 19760 16952 20085 16980
rect 19760 16940 19766 16952
rect 20073 16949 20085 16952
rect 20119 16949 20131 16983
rect 20073 16943 20131 16949
rect 20346 16940 20352 16992
rect 20404 16980 20410 16992
rect 20717 16983 20775 16989
rect 20717 16980 20729 16983
rect 20404 16952 20729 16980
rect 20404 16940 20410 16952
rect 20717 16949 20729 16952
rect 20763 16949 20775 16983
rect 20717 16943 20775 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 2593 16779 2651 16785
rect 2593 16745 2605 16779
rect 2639 16776 2651 16779
rect 3234 16776 3240 16788
rect 2639 16748 3240 16776
rect 2639 16745 2651 16748
rect 2593 16739 2651 16745
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 4157 16779 4215 16785
rect 4157 16745 4169 16779
rect 4203 16776 4215 16779
rect 5534 16776 5540 16788
rect 4203 16748 5540 16776
rect 4203 16745 4215 16748
rect 4157 16739 4215 16745
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 5629 16779 5687 16785
rect 5629 16745 5641 16779
rect 5675 16745 5687 16779
rect 5629 16739 5687 16745
rect 566 16668 572 16720
rect 624 16708 630 16720
rect 4516 16711 4574 16717
rect 624 16680 3096 16708
rect 624 16668 630 16680
rect 1762 16640 1768 16652
rect 1723 16612 1768 16640
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 3068 16649 3096 16680
rect 4516 16677 4528 16711
rect 4562 16708 4574 16711
rect 4706 16708 4712 16720
rect 4562 16680 4712 16708
rect 4562 16677 4574 16680
rect 4516 16671 4574 16677
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 5644 16708 5672 16739
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 6880 16748 8524 16776
rect 6880 16736 6886 16748
rect 5994 16708 6000 16720
rect 5644 16680 6000 16708
rect 5994 16668 6000 16680
rect 6052 16708 6058 16720
rect 6150 16711 6208 16717
rect 6150 16708 6162 16711
rect 6052 16680 6162 16708
rect 6052 16668 6058 16680
rect 6150 16677 6162 16680
rect 6196 16677 6208 16711
rect 6150 16671 6208 16677
rect 7466 16668 7472 16720
rect 7524 16708 7530 16720
rect 7806 16711 7864 16717
rect 7806 16708 7818 16711
rect 7524 16680 7818 16708
rect 7524 16668 7530 16680
rect 7806 16677 7818 16680
rect 7852 16677 7864 16711
rect 8496 16708 8524 16748
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 10502 16776 10508 16788
rect 8628 16748 10508 16776
rect 8628 16736 8634 16748
rect 10502 16736 10508 16748
rect 10560 16736 10566 16788
rect 10689 16779 10747 16785
rect 10689 16745 10701 16779
rect 10735 16776 10747 16779
rect 11517 16779 11575 16785
rect 11517 16776 11529 16779
rect 10735 16748 11529 16776
rect 10735 16745 10747 16748
rect 10689 16739 10747 16745
rect 11517 16745 11529 16748
rect 11563 16745 11575 16779
rect 11517 16739 11575 16745
rect 12989 16779 13047 16785
rect 12989 16745 13001 16779
rect 13035 16776 13047 16779
rect 14461 16779 14519 16785
rect 14461 16776 14473 16779
rect 13035 16748 14473 16776
rect 13035 16745 13047 16748
rect 12989 16739 13047 16745
rect 14461 16745 14473 16748
rect 14507 16745 14519 16779
rect 14461 16739 14519 16745
rect 15010 16736 15016 16788
rect 15068 16776 15074 16788
rect 15289 16779 15347 16785
rect 15289 16776 15301 16779
rect 15068 16748 15301 16776
rect 15068 16736 15074 16748
rect 15289 16745 15301 16748
rect 15335 16745 15347 16779
rect 15289 16739 15347 16745
rect 15749 16779 15807 16785
rect 15749 16745 15761 16779
rect 15795 16776 15807 16779
rect 17494 16776 17500 16788
rect 15795 16748 17500 16776
rect 15795 16745 15807 16748
rect 15749 16739 15807 16745
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 17862 16776 17868 16788
rect 17823 16748 17868 16776
rect 17862 16736 17868 16748
rect 17920 16736 17926 16788
rect 18598 16776 18604 16788
rect 18559 16748 18604 16776
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 18874 16736 18880 16788
rect 18932 16776 18938 16788
rect 20349 16779 20407 16785
rect 20349 16776 20361 16779
rect 18932 16748 20361 16776
rect 18932 16736 18938 16748
rect 20349 16745 20361 16748
rect 20395 16745 20407 16779
rect 20349 16739 20407 16745
rect 10137 16711 10195 16717
rect 10137 16708 10149 16711
rect 8496 16680 10149 16708
rect 7806 16671 7864 16677
rect 10137 16677 10149 16680
rect 10183 16677 10195 16711
rect 10137 16671 10195 16677
rect 10226 16668 10232 16720
rect 10284 16708 10290 16720
rect 13357 16711 13415 16717
rect 13357 16708 13369 16711
rect 10284 16680 13369 16708
rect 10284 16668 10290 16680
rect 13357 16677 13369 16680
rect 13403 16677 13415 16711
rect 13357 16671 13415 16677
rect 13449 16711 13507 16717
rect 13449 16677 13461 16711
rect 13495 16708 13507 16711
rect 13906 16708 13912 16720
rect 13495 16680 13912 16708
rect 13495 16677 13507 16680
rect 13449 16671 13507 16677
rect 13906 16668 13912 16680
rect 13964 16708 13970 16720
rect 14642 16708 14648 16720
rect 13964 16680 14648 16708
rect 13964 16668 13970 16680
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 16752 16711 16810 16717
rect 16752 16677 16764 16711
rect 16798 16708 16810 16711
rect 18322 16708 18328 16720
rect 16798 16680 18328 16708
rect 16798 16677 16810 16680
rect 16752 16671 16810 16677
rect 18322 16668 18328 16680
rect 18380 16668 18386 16720
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2924 16612 2973 16640
rect 2924 16600 2930 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 3053 16643 3111 16649
rect 3053 16609 3065 16643
rect 3099 16640 3111 16643
rect 3099 16612 7144 16640
rect 3099 16609 3111 16612
rect 3053 16603 3111 16609
rect 3237 16575 3295 16581
rect 3237 16541 3249 16575
rect 3283 16572 3295 16575
rect 3326 16572 3332 16584
rect 3283 16544 3332 16572
rect 3283 16541 3295 16544
rect 3237 16535 3295 16541
rect 3326 16532 3332 16544
rect 3384 16532 3390 16584
rect 3602 16532 3608 16584
rect 3660 16572 3666 16584
rect 4157 16575 4215 16581
rect 4157 16572 4169 16575
rect 3660 16544 4169 16572
rect 3660 16532 3666 16544
rect 4157 16541 4169 16544
rect 4203 16572 4215 16575
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 4203 16544 4261 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 5534 16532 5540 16584
rect 5592 16572 5598 16584
rect 5902 16572 5908 16584
rect 5592 16544 5908 16572
rect 5592 16532 5598 16544
rect 5902 16532 5908 16544
rect 5960 16532 5966 16584
rect 7116 16572 7144 16612
rect 7190 16600 7196 16652
rect 7248 16640 7254 16652
rect 7561 16643 7619 16649
rect 7561 16640 7573 16643
rect 7248 16612 7573 16640
rect 7248 16600 7254 16612
rect 7561 16609 7573 16612
rect 7607 16609 7619 16643
rect 8294 16640 8300 16652
rect 7561 16603 7619 16609
rect 7668 16612 8300 16640
rect 7668 16572 7696 16612
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 8444 16612 10057 16640
rect 8444 16600 8450 16612
rect 10045 16609 10057 16612
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 10318 16600 10324 16652
rect 10376 16640 10382 16652
rect 11057 16643 11115 16649
rect 10376 16612 10916 16640
rect 10376 16600 10382 16612
rect 9030 16572 9036 16584
rect 7116 16544 7696 16572
rect 8943 16544 9036 16572
rect 1946 16504 1952 16516
rect 1907 16476 1952 16504
rect 1946 16464 1952 16476
rect 2004 16464 2010 16516
rect 8956 16513 8984 16544
rect 9030 16532 9036 16544
rect 9088 16572 9094 16584
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 9088 16544 10241 16572
rect 9088 16532 9094 16544
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 10888 16572 10916 16612
rect 11057 16609 11069 16643
rect 11103 16640 11115 16643
rect 11238 16640 11244 16652
rect 11103 16612 11244 16640
rect 11103 16609 11115 16612
rect 11057 16603 11115 16609
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16640 11575 16643
rect 12069 16643 12127 16649
rect 12069 16640 12081 16643
rect 11563 16612 12081 16640
rect 11563 16609 11575 16612
rect 11517 16603 11575 16609
rect 12069 16609 12081 16612
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 13078 16600 13084 16652
rect 13136 16640 13142 16652
rect 14369 16643 14427 16649
rect 14369 16640 14381 16643
rect 13136 16612 14381 16640
rect 13136 16600 13142 16612
rect 14369 16609 14381 16612
rect 14415 16609 14427 16643
rect 14369 16603 14427 16609
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15160 16612 15669 16640
rect 15160 16600 15166 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 15930 16640 15936 16652
rect 15804 16612 15936 16640
rect 15804 16600 15810 16612
rect 15930 16600 15936 16612
rect 15988 16640 15994 16652
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 15988 16612 16497 16640
rect 15988 16600 15994 16612
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 16485 16603 16543 16609
rect 18417 16643 18475 16649
rect 18417 16609 18429 16643
rect 18463 16640 18475 16643
rect 19058 16640 19064 16652
rect 18463 16612 19064 16640
rect 18463 16609 18475 16612
rect 18417 16603 18475 16609
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 19242 16649 19248 16652
rect 19236 16640 19248 16649
rect 19203 16612 19248 16640
rect 19236 16603 19248 16612
rect 19242 16600 19248 16603
rect 19300 16600 19306 16652
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 10888 16544 11161 16572
rect 10229 16535 10287 16541
rect 11149 16541 11161 16544
rect 11195 16541 11207 16575
rect 11149 16535 11207 16541
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16541 11391 16575
rect 12158 16572 12164 16584
rect 12119 16544 12164 16572
rect 11333 16535 11391 16541
rect 8941 16507 8999 16513
rect 7208 16476 7512 16504
rect 2038 16396 2044 16448
rect 2096 16436 2102 16448
rect 7208 16436 7236 16476
rect 2096 16408 7236 16436
rect 2096 16396 2102 16408
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 7484 16436 7512 16476
rect 8941 16473 8953 16507
rect 8987 16473 8999 16507
rect 8941 16467 8999 16473
rect 9674 16464 9680 16516
rect 9732 16504 9738 16516
rect 9732 16476 9777 16504
rect 9732 16464 9738 16476
rect 11054 16464 11060 16516
rect 11112 16504 11118 16516
rect 11348 16504 11376 16535
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 13630 16572 13636 16584
rect 12308 16544 12353 16572
rect 13591 16544 13636 16572
rect 12308 16532 12314 16544
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 14550 16572 14556 16584
rect 14511 16544 14556 16572
rect 14550 16532 14556 16544
rect 14608 16532 14614 16584
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 18782 16532 18788 16584
rect 18840 16572 18846 16584
rect 18969 16575 19027 16581
rect 18969 16572 18981 16575
rect 18840 16544 18981 16572
rect 18840 16532 18846 16544
rect 18969 16541 18981 16544
rect 19015 16541 19027 16575
rect 18969 16535 19027 16541
rect 11112 16476 11376 16504
rect 11701 16507 11759 16513
rect 11112 16464 11118 16476
rect 11701 16473 11713 16507
rect 11747 16504 11759 16507
rect 13998 16504 14004 16516
rect 11747 16476 12664 16504
rect 13959 16476 14004 16504
rect 11747 16473 11759 16476
rect 11701 16467 11759 16473
rect 12342 16436 12348 16448
rect 7340 16408 7385 16436
rect 7484 16408 12348 16436
rect 7340 16396 7346 16408
rect 12342 16396 12348 16408
rect 12400 16396 12406 16448
rect 12636 16436 12664 16476
rect 13998 16464 14004 16476
rect 14056 16464 14062 16516
rect 14274 16436 14280 16448
rect 12636 16408 14280 16436
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 14642 16396 14648 16448
rect 14700 16436 14706 16448
rect 17770 16436 17776 16448
rect 14700 16408 17776 16436
rect 14700 16396 14706 16408
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 17862 16396 17868 16448
rect 17920 16436 17926 16448
rect 19978 16436 19984 16448
rect 17920 16408 19984 16436
rect 17920 16396 17926 16408
rect 19978 16396 19984 16408
rect 20036 16396 20042 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 4798 16192 4804 16244
rect 4856 16232 4862 16244
rect 4985 16235 5043 16241
rect 4985 16232 4997 16235
rect 4856 16204 4997 16232
rect 4856 16192 4862 16204
rect 4985 16201 4997 16204
rect 5031 16201 5043 16235
rect 4985 16195 5043 16201
rect 5258 16192 5264 16244
rect 5316 16232 5322 16244
rect 5718 16232 5724 16244
rect 5316 16204 5724 16232
rect 5316 16192 5322 16204
rect 5718 16192 5724 16204
rect 5776 16192 5782 16244
rect 5902 16192 5908 16244
rect 5960 16232 5966 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5960 16204 6009 16232
rect 5960 16192 5966 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 5997 16195 6055 16201
rect 7466 16192 7472 16244
rect 7524 16232 7530 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 7524 16204 8217 16232
rect 7524 16192 7530 16204
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 8205 16195 8263 16201
rect 9398 16192 9404 16244
rect 9456 16232 9462 16244
rect 10318 16232 10324 16244
rect 9456 16204 10324 16232
rect 9456 16192 9462 16204
rect 10318 16192 10324 16204
rect 10376 16192 10382 16244
rect 10505 16235 10563 16241
rect 10505 16201 10517 16235
rect 10551 16232 10563 16235
rect 12158 16232 12164 16244
rect 10551 16204 12164 16232
rect 10551 16201 10563 16204
rect 10505 16195 10563 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 12342 16192 12348 16244
rect 12400 16232 12406 16244
rect 15562 16232 15568 16244
rect 12400 16204 15568 16232
rect 12400 16192 12406 16204
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 16022 16232 16028 16244
rect 15983 16204 16028 16232
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 16206 16192 16212 16244
rect 16264 16232 16270 16244
rect 16485 16235 16543 16241
rect 16485 16232 16497 16235
rect 16264 16204 16497 16232
rect 16264 16192 16270 16204
rect 16485 16201 16497 16204
rect 16531 16201 16543 16235
rect 16850 16232 16856 16244
rect 16811 16204 16856 16232
rect 16485 16195 16543 16201
rect 16850 16192 16856 16204
rect 16908 16192 16914 16244
rect 17034 16192 17040 16244
rect 17092 16232 17098 16244
rect 17092 16204 18828 16232
rect 17092 16192 17098 16204
rect 4433 16167 4491 16173
rect 4433 16133 4445 16167
rect 4479 16164 4491 16167
rect 4706 16164 4712 16176
rect 4479 16136 4712 16164
rect 4479 16133 4491 16136
rect 4433 16127 4491 16133
rect 4706 16124 4712 16136
rect 4764 16164 4770 16176
rect 5166 16164 5172 16176
rect 4764 16136 5172 16164
rect 4764 16124 4770 16136
rect 5166 16124 5172 16136
rect 5224 16124 5230 16176
rect 10137 16167 10195 16173
rect 10137 16133 10149 16167
rect 10183 16133 10195 16167
rect 10137 16127 10195 16133
rect 5258 16056 5264 16108
rect 5316 16096 5322 16108
rect 5537 16099 5595 16105
rect 5537 16096 5549 16099
rect 5316 16068 5549 16096
rect 5316 16056 5322 16068
rect 5537 16065 5549 16068
rect 5583 16065 5595 16099
rect 5537 16059 5595 16065
rect 6196 16068 6960 16096
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 15997 1823 16031
rect 2314 16028 2320 16040
rect 2275 16000 2320 16028
rect 1765 15991 1823 15997
rect 1780 15960 1808 15991
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 3050 16028 3056 16040
rect 2963 16000 3056 16028
rect 3050 15988 3056 16000
rect 3108 16028 3114 16040
rect 3602 16028 3608 16040
rect 3108 16000 3608 16028
rect 3108 15988 3114 16000
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 5442 16028 5448 16040
rect 5403 16000 5448 16028
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 6196 16037 6224 16068
rect 6932 16040 6960 16068
rect 8478 16056 8484 16108
rect 8536 16096 8542 16108
rect 8757 16099 8815 16105
rect 8757 16096 8769 16099
rect 8536 16068 8769 16096
rect 8536 16056 8542 16068
rect 8757 16065 8769 16068
rect 8803 16065 8815 16099
rect 10152 16096 10180 16127
rect 11330 16124 11336 16176
rect 11388 16164 11394 16176
rect 12621 16167 12679 16173
rect 12621 16164 12633 16167
rect 11388 16136 12633 16164
rect 11388 16124 11394 16136
rect 12621 16133 12633 16136
rect 12667 16164 12679 16167
rect 12894 16164 12900 16176
rect 12667 16136 12900 16164
rect 12667 16133 12679 16136
rect 12621 16127 12679 16133
rect 12894 16124 12900 16136
rect 12952 16164 12958 16176
rect 12952 16136 13032 16164
rect 12952 16124 12958 16136
rect 11054 16096 11060 16108
rect 10152 16068 11060 16096
rect 8757 16059 8815 16065
rect 11054 16056 11060 16068
rect 11112 16096 11118 16108
rect 11149 16099 11207 16105
rect 11149 16096 11161 16099
rect 11112 16068 11161 16096
rect 11112 16056 11118 16068
rect 11149 16065 11161 16068
rect 11195 16096 11207 16099
rect 11698 16096 11704 16108
rect 11195 16068 11704 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16096 11943 16099
rect 11974 16096 11980 16108
rect 11931 16068 11980 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 11974 16056 11980 16068
rect 12032 16056 12038 16108
rect 13004 16105 13032 16136
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13998 16056 14004 16108
rect 14056 16096 14062 16108
rect 17497 16099 17555 16105
rect 14056 16068 14780 16096
rect 14056 16056 14062 16068
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 15997 6239 16031
rect 6181 15991 6239 15997
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 3142 15960 3148 15972
rect 1780 15932 3148 15960
rect 3142 15920 3148 15932
rect 3200 15920 3206 15972
rect 3320 15963 3378 15969
rect 3320 15929 3332 15963
rect 3366 15960 3378 15963
rect 3418 15960 3424 15972
rect 3366 15932 3424 15960
rect 3366 15929 3378 15932
rect 3320 15923 3378 15929
rect 3418 15920 3424 15932
rect 3476 15920 3482 15972
rect 3970 15920 3976 15972
rect 4028 15960 4034 15972
rect 6638 15960 6644 15972
rect 4028 15932 6644 15960
rect 4028 15920 4034 15932
rect 6638 15920 6644 15932
rect 6696 15920 6702 15972
rect 1946 15892 1952 15904
rect 1907 15864 1952 15892
rect 1946 15852 1952 15864
rect 2004 15852 2010 15904
rect 2498 15892 2504 15904
rect 2459 15864 2504 15892
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 5074 15852 5080 15904
rect 5132 15892 5138 15904
rect 5353 15895 5411 15901
rect 5353 15892 5365 15895
rect 5132 15864 5365 15892
rect 5132 15852 5138 15864
rect 5353 15861 5365 15864
rect 5399 15861 5411 15895
rect 6840 15892 6868 15991
rect 6914 15988 6920 16040
rect 6972 16028 6978 16040
rect 9030 16037 9036 16040
rect 8665 16031 8723 16037
rect 8665 16028 8677 16031
rect 6972 16000 8677 16028
rect 6972 15988 6978 16000
rect 8665 15997 8677 16000
rect 8711 15997 8723 16031
rect 9024 16028 9036 16037
rect 8991 16000 9036 16028
rect 8665 15991 8723 15997
rect 9024 15991 9036 16000
rect 9030 15988 9036 15991
rect 9088 15988 9094 16040
rect 10962 16028 10968 16040
rect 10923 16000 10968 16028
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 11609 16031 11667 16037
rect 11609 15997 11621 16031
rect 11655 16028 11667 16031
rect 12342 16028 12348 16040
rect 11655 16000 12348 16028
rect 11655 15997 11667 16000
rect 11609 15991 11667 15997
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 12805 16031 12863 16037
rect 12805 15997 12817 16031
rect 12851 15997 12863 16031
rect 12805 15991 12863 15997
rect 13256 16031 13314 16037
rect 13256 15997 13268 16031
rect 13302 16028 13314 16031
rect 13630 16028 13636 16040
rect 13302 16000 13636 16028
rect 13302 15997 13314 16000
rect 13256 15991 13314 15997
rect 7092 15963 7150 15969
rect 7092 15929 7104 15963
rect 7138 15960 7150 15963
rect 7282 15960 7288 15972
rect 7138 15932 7288 15960
rect 7138 15929 7150 15932
rect 7092 15923 7150 15929
rect 7282 15920 7288 15932
rect 7340 15960 7346 15972
rect 8938 15960 8944 15972
rect 7340 15932 8944 15960
rect 7340 15920 7346 15932
rect 8938 15920 8944 15932
rect 8996 15920 9002 15972
rect 9306 15920 9312 15972
rect 9364 15960 9370 15972
rect 10226 15960 10232 15972
rect 9364 15932 10232 15960
rect 9364 15920 9370 15932
rect 10226 15920 10232 15932
rect 10284 15920 10290 15972
rect 10778 15920 10784 15972
rect 10836 15960 10842 15972
rect 10873 15963 10931 15969
rect 10873 15960 10885 15963
rect 10836 15932 10885 15960
rect 10836 15920 10842 15932
rect 10873 15929 10885 15932
rect 10919 15929 10931 15963
rect 12820 15960 12848 15991
rect 13630 15988 13636 16000
rect 13688 15988 13694 16040
rect 14645 16031 14703 16037
rect 14645 16028 14657 16031
rect 14016 16000 14657 16028
rect 13906 15960 13912 15972
rect 12820 15932 13912 15960
rect 10873 15923 10931 15929
rect 13906 15920 13912 15932
rect 13964 15920 13970 15972
rect 7190 15892 7196 15904
rect 6840 15864 7196 15892
rect 5353 15855 5411 15861
rect 7190 15852 7196 15864
rect 7248 15892 7254 15904
rect 8478 15892 8484 15904
rect 7248 15864 8484 15892
rect 7248 15852 7254 15864
rect 8478 15852 8484 15864
rect 8536 15852 8542 15904
rect 12894 15852 12900 15904
rect 12952 15892 12958 15904
rect 14016 15892 14044 16000
rect 14645 15997 14657 16000
rect 14691 15997 14703 16031
rect 14752 16028 14780 16068
rect 15672 16068 17356 16096
rect 15672 16028 15700 16068
rect 14752 16000 15700 16028
rect 16301 16031 16359 16037
rect 14645 15991 14703 15997
rect 16301 15997 16313 16031
rect 16347 16028 16359 16031
rect 17218 16028 17224 16040
rect 16347 16000 17224 16028
rect 16347 15997 16359 16000
rect 16301 15991 16359 15997
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 17328 16028 17356 16068
rect 17497 16065 17509 16099
rect 17543 16096 17555 16099
rect 18046 16096 18052 16108
rect 17543 16068 18052 16096
rect 17543 16065 17555 16068
rect 17497 16059 17555 16065
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 18800 16096 18828 16204
rect 19242 16192 19248 16244
rect 19300 16232 19306 16244
rect 20257 16235 20315 16241
rect 20257 16232 20269 16235
rect 19300 16204 20269 16232
rect 19300 16192 19306 16204
rect 20257 16201 20269 16204
rect 20303 16201 20315 16235
rect 20257 16195 20315 16201
rect 18800 16068 19012 16096
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 17328 16000 18337 16028
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 18414 15988 18420 16040
rect 18472 16028 18478 16040
rect 18782 16028 18788 16040
rect 18472 16000 18788 16028
rect 18472 15988 18478 16000
rect 18782 15988 18788 16000
rect 18840 16028 18846 16040
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18840 16000 18889 16028
rect 18840 15988 18846 16000
rect 18877 15997 18889 16000
rect 18923 15997 18935 16031
rect 18984 16028 19012 16068
rect 18984 16000 19932 16028
rect 18877 15991 18935 15997
rect 14550 15960 14556 15972
rect 14384 15932 14556 15960
rect 14384 15904 14412 15932
rect 14550 15920 14556 15932
rect 14608 15960 14614 15972
rect 14890 15963 14948 15969
rect 14890 15960 14902 15963
rect 14608 15932 14902 15960
rect 14608 15920 14614 15932
rect 14890 15929 14902 15932
rect 14936 15929 14948 15963
rect 14890 15923 14948 15929
rect 15194 15920 15200 15972
rect 15252 15960 15258 15972
rect 17034 15960 17040 15972
rect 15252 15932 17040 15960
rect 15252 15920 15258 15932
rect 17034 15920 17040 15932
rect 17092 15920 17098 15972
rect 18598 15960 18604 15972
rect 17236 15932 18604 15960
rect 14366 15892 14372 15904
rect 12952 15864 14044 15892
rect 14327 15864 14372 15892
rect 12952 15852 12958 15864
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 17236 15901 17264 15932
rect 18598 15920 18604 15932
rect 18656 15920 18662 15972
rect 19144 15963 19202 15969
rect 19144 15929 19156 15963
rect 19190 15960 19202 15963
rect 19610 15960 19616 15972
rect 19190 15932 19616 15960
rect 19190 15929 19202 15932
rect 19144 15923 19202 15929
rect 19610 15920 19616 15932
rect 19668 15920 19674 15972
rect 19904 15960 19932 16000
rect 19978 15988 19984 16040
rect 20036 16028 20042 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20036 16000 20545 16028
rect 20036 15988 20042 16000
rect 20533 15997 20545 16000
rect 20579 16028 20591 16031
rect 21082 16028 21088 16040
rect 20579 16000 21088 16028
rect 20579 15997 20591 16000
rect 20533 15991 20591 15997
rect 21082 15988 21088 16000
rect 21140 15988 21146 16040
rect 20162 15960 20168 15972
rect 19904 15932 20168 15960
rect 20162 15920 20168 15932
rect 20220 15960 20226 15972
rect 20990 15960 20996 15972
rect 20220 15932 20996 15960
rect 20220 15920 20226 15932
rect 20990 15920 20996 15932
rect 21048 15920 21054 15972
rect 17221 15895 17279 15901
rect 17221 15861 17233 15895
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 18506 15892 18512 15904
rect 17368 15864 17413 15892
rect 18467 15864 18512 15892
rect 17368 15852 17374 15864
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 20717 15895 20775 15901
rect 20717 15892 20729 15895
rect 20680 15864 20729 15892
rect 20680 15852 20686 15864
rect 20717 15861 20729 15864
rect 20763 15861 20775 15895
rect 20717 15855 20775 15861
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 3234 15688 3240 15700
rect 3195 15660 3240 15688
rect 3234 15648 3240 15660
rect 3292 15648 3298 15700
rect 4617 15691 4675 15697
rect 4617 15657 4629 15691
rect 4663 15657 4675 15691
rect 4617 15651 4675 15657
rect 5077 15691 5135 15697
rect 5077 15657 5089 15691
rect 5123 15688 5135 15691
rect 5534 15688 5540 15700
rect 5123 15660 5540 15688
rect 5123 15657 5135 15660
rect 5077 15651 5135 15657
rect 3145 15623 3203 15629
rect 3145 15589 3157 15623
rect 3191 15620 3203 15623
rect 3510 15620 3516 15632
rect 3191 15592 3516 15620
rect 3191 15589 3203 15592
rect 3145 15583 3203 15589
rect 3510 15580 3516 15592
rect 3568 15580 3574 15632
rect 4632 15620 4660 15651
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 5629 15691 5687 15697
rect 5629 15657 5641 15691
rect 5675 15688 5687 15691
rect 5810 15688 5816 15700
rect 5675 15660 5816 15688
rect 5675 15657 5687 15660
rect 5629 15651 5687 15657
rect 5810 15648 5816 15660
rect 5868 15648 5874 15700
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 7423 15660 8033 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 8021 15657 8033 15660
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 11882 15688 11888 15700
rect 8527 15660 11888 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 11977 15691 12035 15697
rect 11977 15657 11989 15691
rect 12023 15688 12035 15691
rect 12023 15660 12296 15688
rect 12023 15657 12035 15660
rect 11977 15651 12035 15657
rect 5997 15623 6055 15629
rect 5997 15620 6009 15623
rect 4632 15592 6009 15620
rect 5997 15589 6009 15592
rect 6043 15589 6055 15623
rect 5997 15583 6055 15589
rect 6638 15580 6644 15632
rect 6696 15620 6702 15632
rect 8662 15620 8668 15632
rect 6696 15592 8668 15620
rect 6696 15580 6702 15592
rect 8662 15580 8668 15592
rect 8720 15580 8726 15632
rect 11330 15620 11336 15632
rect 10612 15592 11336 15620
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 3602 15552 3608 15564
rect 1811 15524 3608 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 3602 15512 3608 15524
rect 3660 15512 3666 15564
rect 4982 15552 4988 15564
rect 4943 15524 4988 15552
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 5166 15512 5172 15564
rect 5224 15552 5230 15564
rect 7469 15555 7527 15561
rect 5224 15524 6224 15552
rect 5224 15512 5230 15524
rect 3418 15484 3424 15496
rect 3331 15456 3424 15484
rect 3418 15444 3424 15456
rect 3476 15484 3482 15496
rect 5258 15484 5264 15496
rect 3476 15456 5028 15484
rect 5219 15456 5264 15484
rect 3476 15444 3482 15456
rect 2777 15419 2835 15425
rect 2777 15385 2789 15419
rect 2823 15416 2835 15419
rect 4890 15416 4896 15428
rect 2823 15388 4896 15416
rect 2823 15385 2835 15388
rect 2777 15379 2835 15385
rect 4890 15376 4896 15388
rect 4948 15376 4954 15428
rect 5000 15416 5028 15456
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 6196 15493 6224 15524
rect 7469 15521 7481 15555
rect 7515 15552 7527 15555
rect 8294 15552 8300 15564
rect 7515 15524 8300 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 10612 15561 10640 15592
rect 11330 15580 11336 15592
rect 11388 15620 11394 15632
rect 12161 15623 12219 15629
rect 12161 15620 12173 15623
rect 11388 15592 12173 15620
rect 11388 15580 11394 15592
rect 12161 15589 12173 15592
rect 12207 15589 12219 15623
rect 12268 15620 12296 15660
rect 12342 15648 12348 15700
rect 12400 15688 12406 15700
rect 13909 15691 13967 15697
rect 13909 15688 13921 15691
rect 12400 15660 13921 15688
rect 12400 15648 12406 15660
rect 13909 15657 13921 15660
rect 13955 15657 13967 15691
rect 13909 15651 13967 15657
rect 14274 15648 14280 15700
rect 14332 15688 14338 15700
rect 14369 15691 14427 15697
rect 14369 15688 14381 15691
rect 14332 15660 14381 15688
rect 14332 15648 14338 15660
rect 14369 15657 14381 15660
rect 14415 15657 14427 15691
rect 14369 15651 14427 15657
rect 14476 15660 17448 15688
rect 12520 15623 12578 15629
rect 12520 15620 12532 15623
rect 12268 15592 12532 15620
rect 12161 15583 12219 15589
rect 12520 15589 12532 15592
rect 12566 15620 12578 15623
rect 13725 15623 13783 15629
rect 13725 15620 13737 15623
rect 12566 15592 13737 15620
rect 12566 15589 12578 15592
rect 12520 15583 12578 15589
rect 13725 15589 13737 15592
rect 13771 15589 13783 15623
rect 14476 15620 14504 15660
rect 13725 15583 13783 15589
rect 13823 15592 14504 15620
rect 15648 15623 15706 15629
rect 10870 15561 10876 15564
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15552 8447 15555
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 8435 15524 9045 15552
rect 8435 15521 8447 15524
rect 8389 15515 8447 15521
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 9033 15515 9091 15521
rect 10597 15555 10655 15561
rect 10597 15521 10609 15555
rect 10643 15521 10655 15555
rect 10864 15552 10876 15561
rect 10831 15524 10876 15552
rect 10597 15515 10655 15521
rect 10864 15515 10876 15524
rect 10870 15512 10876 15515
rect 10928 15512 10934 15564
rect 13823 15552 13851 15592
rect 15648 15589 15660 15623
rect 15694 15620 15706 15623
rect 16022 15620 16028 15632
rect 15694 15592 16028 15620
rect 15694 15589 15706 15592
rect 15648 15583 15706 15589
rect 16022 15580 16028 15592
rect 16080 15580 16086 15632
rect 14274 15552 14280 15564
rect 12084 15524 13851 15552
rect 14235 15524 14280 15552
rect 5537 15487 5595 15493
rect 5537 15453 5549 15487
rect 5583 15484 5595 15487
rect 6089 15487 6147 15493
rect 6089 15484 6101 15487
rect 5583 15456 6101 15484
rect 5583 15453 5595 15456
rect 5537 15447 5595 15453
rect 6089 15453 6101 15456
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 6181 15487 6239 15493
rect 6181 15453 6193 15487
rect 6227 15453 6239 15487
rect 7558 15484 7564 15496
rect 7519 15456 7564 15484
rect 6181 15447 6239 15453
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 8665 15487 8723 15493
rect 8665 15453 8677 15487
rect 8711 15484 8723 15487
rect 8938 15484 8944 15496
rect 8711 15456 8944 15484
rect 8711 15453 8723 15456
rect 8665 15447 8723 15453
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 5276 15416 5304 15444
rect 5000 15388 5304 15416
rect 7009 15419 7067 15425
rect 7009 15385 7021 15419
rect 7055 15416 7067 15419
rect 8386 15416 8392 15428
rect 7055 15388 8392 15416
rect 7055 15385 7067 15388
rect 7009 15379 7067 15385
rect 8386 15376 8392 15388
rect 8444 15376 8450 15428
rect 1946 15348 1952 15360
rect 1907 15320 1952 15348
rect 1946 15308 1952 15320
rect 2004 15308 2010 15360
rect 2314 15308 2320 15360
rect 2372 15348 2378 15360
rect 3970 15348 3976 15360
rect 2372 15320 3976 15348
rect 2372 15308 2378 15320
rect 3970 15308 3976 15320
rect 4028 15308 4034 15360
rect 4154 15308 4160 15360
rect 4212 15348 4218 15360
rect 5537 15351 5595 15357
rect 5537 15348 5549 15351
rect 4212 15320 5549 15348
rect 4212 15308 4218 15320
rect 5537 15317 5549 15320
rect 5583 15317 5595 15351
rect 5537 15311 5595 15317
rect 6270 15308 6276 15360
rect 6328 15348 6334 15360
rect 12084 15348 12112 15524
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 15381 15555 15439 15561
rect 15381 15521 15393 15555
rect 15427 15552 15439 15555
rect 15930 15552 15936 15564
rect 15427 15524 15936 15552
rect 15427 15521 15439 15524
rect 15381 15515 15439 15521
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 17420 15561 17448 15660
rect 17954 15648 17960 15700
rect 18012 15688 18018 15700
rect 18049 15691 18107 15697
rect 18049 15688 18061 15691
rect 18012 15660 18061 15688
rect 18012 15648 18018 15660
rect 18049 15657 18061 15660
rect 18095 15657 18107 15691
rect 18690 15688 18696 15700
rect 18049 15651 18107 15657
rect 18156 15660 18696 15688
rect 17494 15580 17500 15632
rect 17552 15620 17558 15632
rect 18156 15620 18184 15660
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 19061 15691 19119 15697
rect 19061 15657 19073 15691
rect 19107 15688 19119 15691
rect 19518 15688 19524 15700
rect 19107 15660 19524 15688
rect 19107 15657 19119 15660
rect 19061 15651 19119 15657
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 17552 15592 18184 15620
rect 18417 15623 18475 15629
rect 17552 15580 17558 15592
rect 18417 15589 18429 15623
rect 18463 15620 18475 15623
rect 19702 15620 19708 15632
rect 18463 15592 19708 15620
rect 18463 15589 18475 15592
rect 18417 15583 18475 15589
rect 19702 15580 19708 15592
rect 19760 15580 19766 15632
rect 20349 15623 20407 15629
rect 20349 15589 20361 15623
rect 20395 15620 20407 15623
rect 20530 15620 20536 15632
rect 20395 15592 20536 15620
rect 20395 15589 20407 15592
rect 20349 15583 20407 15589
rect 20530 15580 20536 15592
rect 20588 15580 20594 15632
rect 17405 15555 17463 15561
rect 17405 15521 17417 15555
rect 17451 15552 17463 15555
rect 18509 15555 18567 15561
rect 17451 15524 17724 15552
rect 17451 15521 17463 15524
rect 17405 15515 17463 15521
rect 12161 15487 12219 15493
rect 12161 15453 12173 15487
rect 12207 15484 12219 15487
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 12207 15456 12265 15484
rect 12207 15453 12219 15456
rect 12161 15447 12219 15453
rect 12253 15453 12265 15456
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 17589 15487 17647 15493
rect 17589 15453 17601 15487
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 6328 15320 12112 15348
rect 12268 15348 12296 15447
rect 13725 15419 13783 15425
rect 13725 15385 13737 15419
rect 13771 15416 13783 15419
rect 14476 15416 14504 15447
rect 13771 15388 14504 15416
rect 13771 15385 13783 15388
rect 13725 15379 13783 15385
rect 16574 15376 16580 15428
rect 16632 15416 16638 15428
rect 16761 15419 16819 15425
rect 16761 15416 16773 15419
rect 16632 15388 16773 15416
rect 16632 15376 16638 15388
rect 16761 15385 16773 15388
rect 16807 15416 16819 15419
rect 17604 15416 17632 15447
rect 16807 15388 17632 15416
rect 16807 15385 16819 15388
rect 16761 15379 16819 15385
rect 12618 15348 12624 15360
rect 12268 15320 12624 15348
rect 6328 15308 6334 15320
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 13630 15348 13636 15360
rect 13543 15320 13636 15348
rect 13630 15308 13636 15320
rect 13688 15348 13694 15360
rect 15746 15348 15752 15360
rect 13688 15320 15752 15348
rect 13688 15308 13694 15320
rect 15746 15308 15752 15320
rect 15804 15308 15810 15360
rect 17034 15348 17040 15360
rect 16995 15320 17040 15348
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 17586 15348 17592 15360
rect 17276 15320 17592 15348
rect 17276 15308 17282 15320
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 17696 15348 17724 15524
rect 18509 15521 18521 15555
rect 18555 15552 18567 15555
rect 19334 15552 19340 15564
rect 18555 15524 19340 15552
rect 18555 15521 18567 15524
rect 18509 15515 18567 15521
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 19886 15552 19892 15564
rect 19475 15524 19892 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 19886 15512 19892 15524
rect 19944 15512 19950 15564
rect 20070 15552 20076 15564
rect 20031 15524 20076 15552
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 18693 15487 18751 15493
rect 18693 15453 18705 15487
rect 18739 15484 18751 15487
rect 19242 15484 19248 15496
rect 18739 15456 19248 15484
rect 18739 15453 18751 15456
rect 18693 15447 18751 15453
rect 19242 15444 19248 15456
rect 19300 15444 19306 15496
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 17770 15376 17776 15428
rect 17828 15416 17834 15428
rect 19536 15416 19564 15447
rect 19610 15444 19616 15496
rect 19668 15484 19674 15496
rect 19668 15456 19713 15484
rect 19668 15444 19674 15456
rect 17828 15388 19564 15416
rect 17828 15376 17834 15388
rect 18874 15348 18880 15360
rect 17696 15320 18880 15348
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 4157 15147 4215 15153
rect 4157 15144 4169 15147
rect 1596 15116 4169 15144
rect 1596 14949 1624 15116
rect 4157 15113 4169 15116
rect 4203 15113 4215 15147
rect 4157 15107 4215 15113
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 7377 15147 7435 15153
rect 7377 15144 7389 15147
rect 7064 15116 7389 15144
rect 7064 15104 7070 15116
rect 7377 15113 7389 15116
rect 7423 15113 7435 15147
rect 7377 15107 7435 15113
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8389 15147 8447 15153
rect 8389 15144 8401 15147
rect 8352 15116 8401 15144
rect 8352 15104 8358 15116
rect 8389 15113 8401 15116
rect 8435 15113 8447 15147
rect 8389 15107 8447 15113
rect 10870 15104 10876 15156
rect 10928 15144 10934 15156
rect 11057 15147 11115 15153
rect 11057 15144 11069 15147
rect 10928 15116 11069 15144
rect 10928 15104 10934 15116
rect 11057 15113 11069 15116
rect 11103 15144 11115 15147
rect 11882 15144 11888 15156
rect 11103 15116 11888 15144
rect 11103 15113 11115 15116
rect 11057 15107 11115 15113
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 13265 15147 13323 15153
rect 12360 15116 12572 15144
rect 3418 15036 3424 15088
rect 3476 15076 3482 15088
rect 3697 15079 3755 15085
rect 3697 15076 3709 15079
rect 3476 15048 3709 15076
rect 3476 15036 3482 15048
rect 3697 15045 3709 15048
rect 3743 15045 3755 15079
rect 3697 15039 3755 15045
rect 6196 15048 9076 15076
rect 1854 15008 1860 15020
rect 1815 14980 1860 15008
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 4801 15011 4859 15017
rect 4801 14977 4813 15011
rect 4847 14977 4859 15011
rect 4801 14971 4859 14977
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14909 1639 14943
rect 1581 14903 1639 14909
rect 2317 14943 2375 14949
rect 2317 14909 2329 14943
rect 2363 14940 2375 14943
rect 3050 14940 3056 14952
rect 2363 14912 3056 14940
rect 2363 14909 2375 14912
rect 2317 14903 2375 14909
rect 3050 14900 3056 14912
rect 3108 14940 3114 14952
rect 3970 14940 3976 14952
rect 3108 14912 3976 14940
rect 3108 14900 3114 14912
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 4816 14940 4844 14971
rect 4982 14968 4988 15020
rect 5040 15008 5046 15020
rect 6196 15017 6224 15048
rect 5169 15011 5227 15017
rect 5169 15008 5181 15011
rect 5040 14980 5181 15008
rect 5040 14968 5046 14980
rect 5169 14977 5181 14980
rect 5215 14977 5227 15011
rect 5169 14971 5227 14977
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 14977 6239 15011
rect 6181 14971 6239 14977
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 6638 15008 6644 15020
rect 6411 14980 6644 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 7190 15008 7196 15020
rect 7064 14980 7196 15008
rect 7064 14968 7070 14980
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 8754 15008 8760 15020
rect 8067 14980 8760 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 8754 14968 8760 14980
rect 8812 14968 8818 15020
rect 8938 15008 8944 15020
rect 8899 14980 8944 15008
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 9048 15008 9076 15048
rect 9674 15036 9680 15088
rect 9732 15036 9738 15088
rect 11333 15079 11391 15085
rect 11333 15045 11345 15079
rect 11379 15076 11391 15079
rect 12360 15076 12388 15116
rect 11379 15048 12388 15076
rect 12544 15076 12572 15116
rect 13265 15113 13277 15147
rect 13311 15144 13323 15147
rect 14274 15144 14280 15156
rect 13311 15116 14280 15144
rect 13311 15113 13323 15116
rect 13265 15107 13323 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 19429 15147 19487 15153
rect 16316 15116 18000 15144
rect 14090 15076 14096 15088
rect 12544 15048 13645 15076
rect 14051 15048 14096 15076
rect 11379 15045 11391 15048
rect 11333 15039 11391 15045
rect 9692 15008 9720 15036
rect 9048 14980 9720 15008
rect 11698 14968 11704 15020
rect 11756 15008 11762 15020
rect 11977 15011 12035 15017
rect 11977 15008 11989 15011
rect 11756 14980 11989 15008
rect 11756 14968 11762 14980
rect 11977 14977 11989 14980
rect 12023 15008 12035 15011
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12023 14980 13001 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 13617 15008 13645 15048
rect 14090 15036 14096 15048
rect 14148 15036 14154 15088
rect 16316 15076 16344 15116
rect 14292 15048 16344 15076
rect 13814 15008 13820 15020
rect 13617 14980 13676 15008
rect 13775 14980 13820 15008
rect 12989 14971 13047 14977
rect 5442 14940 5448 14952
rect 4816 14912 5448 14940
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14940 6147 14943
rect 6270 14940 6276 14952
rect 6135 14912 6276 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 7208 14940 7236 14968
rect 9674 14940 9680 14952
rect 7208 14912 9680 14940
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 9944 14943 10002 14949
rect 9944 14909 9956 14943
rect 9990 14940 10002 14943
rect 11716 14940 11744 14968
rect 13648 14949 13676 14980
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 13633 14943 13691 14949
rect 9990 14912 11744 14940
rect 12452 14912 13124 14940
rect 9990 14909 10002 14912
rect 9944 14903 10002 14909
rect 2584 14875 2642 14881
rect 2584 14841 2596 14875
rect 2630 14872 2642 14875
rect 3234 14872 3240 14884
rect 2630 14844 3240 14872
rect 2630 14841 2642 14844
rect 2584 14835 2642 14841
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 4246 14832 4252 14884
rect 4304 14872 4310 14884
rect 4525 14875 4583 14881
rect 4525 14872 4537 14875
rect 4304 14844 4537 14872
rect 4304 14832 4310 14844
rect 4525 14841 4537 14844
rect 4571 14841 4583 14875
rect 4525 14835 4583 14841
rect 8662 14832 8668 14884
rect 8720 14872 8726 14884
rect 8757 14875 8815 14881
rect 8757 14872 8769 14875
rect 8720 14844 8769 14872
rect 8720 14832 8726 14844
rect 8757 14841 8769 14844
rect 8803 14841 8815 14875
rect 8757 14835 8815 14841
rect 8849 14875 8907 14881
rect 8849 14841 8861 14875
rect 8895 14872 8907 14875
rect 8938 14872 8944 14884
rect 8895 14844 8944 14872
rect 8895 14841 8907 14844
rect 8849 14835 8907 14841
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 11698 14872 11704 14884
rect 11659 14844 11704 14872
rect 11698 14832 11704 14844
rect 11756 14832 11762 14884
rect 4614 14804 4620 14816
rect 4575 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 4706 14764 4712 14816
rect 4764 14804 4770 14816
rect 5721 14807 5779 14813
rect 5721 14804 5733 14807
rect 4764 14776 5733 14804
rect 4764 14764 4770 14776
rect 5721 14773 5733 14776
rect 5767 14773 5779 14807
rect 7742 14804 7748 14816
rect 7703 14776 7748 14804
rect 5721 14767 5779 14773
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 7837 14807 7895 14813
rect 7837 14773 7849 14807
rect 7883 14804 7895 14807
rect 8294 14804 8300 14816
rect 7883 14776 8300 14804
rect 7883 14773 7895 14776
rect 7837 14767 7895 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 11514 14804 11520 14816
rect 9088 14776 11520 14804
rect 9088 14764 9094 14776
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 11790 14804 11796 14816
rect 11751 14776 11796 14804
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 12452 14813 12480 14912
rect 12897 14875 12955 14881
rect 12897 14841 12909 14875
rect 12943 14872 12955 14875
rect 12986 14872 12992 14884
rect 12943 14844 12992 14872
rect 12943 14841 12955 14844
rect 12897 14835 12955 14841
rect 12986 14832 12992 14844
rect 13044 14832 13050 14884
rect 13096 14872 13124 14912
rect 13633 14909 13645 14943
rect 13679 14909 13691 14943
rect 14292 14940 14320 15048
rect 17586 15036 17592 15088
rect 17644 15076 17650 15088
rect 17681 15079 17739 15085
rect 17681 15076 17693 15079
rect 17644 15048 17693 15076
rect 17644 15036 17650 15048
rect 17681 15045 17693 15048
rect 17727 15045 17739 15079
rect 17681 15039 17739 15045
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 14424 14980 14657 15008
rect 14424 14968 14430 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 15008 15623 15011
rect 15838 15008 15844 15020
rect 15611 14980 15844 15008
rect 15611 14977 15623 14980
rect 15565 14971 15623 14977
rect 15838 14968 15844 14980
rect 15896 14968 15902 15020
rect 17972 15008 18000 15116
rect 18064 15116 19012 15144
rect 18064 15088 18092 15116
rect 18046 15036 18052 15088
rect 18104 15036 18110 15088
rect 18984 15076 19012 15116
rect 19429 15113 19441 15147
rect 19475 15144 19487 15147
rect 19610 15144 19616 15156
rect 19475 15116 19616 15144
rect 19475 15113 19487 15116
rect 19429 15107 19487 15113
rect 19610 15104 19616 15116
rect 19668 15104 19674 15156
rect 18984 15048 20576 15076
rect 16040 14980 16436 15008
rect 17972 14980 18184 15008
rect 13633 14903 13691 14909
rect 13832 14912 14320 14940
rect 14461 14943 14519 14949
rect 13725 14875 13783 14881
rect 13725 14872 13737 14875
rect 13096 14844 13737 14872
rect 13725 14841 13737 14844
rect 13771 14841 13783 14875
rect 13725 14835 13783 14841
rect 12437 14807 12495 14813
rect 12437 14773 12449 14807
rect 12483 14773 12495 14807
rect 12437 14767 12495 14773
rect 12805 14807 12863 14813
rect 12805 14773 12817 14807
rect 12851 14804 12863 14807
rect 13832 14804 13860 14912
rect 14461 14909 14473 14943
rect 14507 14940 14519 14943
rect 15010 14940 15016 14952
rect 14507 14912 15016 14940
rect 14507 14909 14519 14912
rect 14461 14903 14519 14909
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14940 15347 14943
rect 16040 14940 16068 14980
rect 15335 14912 16068 14940
rect 16117 14943 16175 14949
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 16117 14909 16129 14943
rect 16163 14909 16175 14943
rect 16117 14903 16175 14909
rect 16301 14943 16359 14949
rect 16301 14909 16313 14943
rect 16347 14909 16359 14943
rect 16301 14903 16359 14909
rect 13906 14832 13912 14884
rect 13964 14872 13970 14884
rect 16132 14872 16160 14903
rect 13964 14844 16160 14872
rect 13964 14832 13970 14844
rect 12851 14776 13860 14804
rect 14553 14807 14611 14813
rect 12851 14773 12863 14776
rect 12805 14767 12863 14773
rect 14553 14773 14565 14807
rect 14599 14804 14611 14807
rect 14921 14807 14979 14813
rect 14921 14804 14933 14807
rect 14599 14776 14933 14804
rect 14599 14773 14611 14776
rect 14553 14767 14611 14773
rect 14921 14773 14933 14776
rect 14967 14773 14979 14807
rect 14921 14767 14979 14773
rect 15381 14807 15439 14813
rect 15381 14773 15393 14807
rect 15427 14804 15439 14807
rect 15838 14804 15844 14816
rect 15427 14776 15844 14804
rect 15427 14773 15439 14776
rect 15381 14767 15439 14773
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 15933 14807 15991 14813
rect 15933 14773 15945 14807
rect 15979 14804 15991 14807
rect 16022 14804 16028 14816
rect 15979 14776 16028 14804
rect 15979 14773 15991 14776
rect 15933 14767 15991 14773
rect 16022 14764 16028 14776
rect 16080 14804 16086 14816
rect 16316 14804 16344 14903
rect 16408 14872 16436 14980
rect 16574 14949 16580 14952
rect 16568 14940 16580 14949
rect 16535 14912 16580 14940
rect 16568 14903 16580 14912
rect 16574 14900 16580 14903
rect 16632 14900 16638 14952
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17604 14912 18061 14940
rect 17494 14872 17500 14884
rect 16408 14844 17500 14872
rect 17494 14832 17500 14844
rect 17552 14832 17558 14884
rect 17604 14804 17632 14912
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18156 14940 18184 14980
rect 19058 14968 19064 15020
rect 19116 15008 19122 15020
rect 19981 15011 20039 15017
rect 19981 15008 19993 15011
rect 19116 14980 19993 15008
rect 19116 14968 19122 14980
rect 19981 14977 19993 14980
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 18782 14940 18788 14952
rect 18156 14912 18788 14940
rect 18049 14903 18107 14909
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 20548 14949 20576 15048
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14909 19855 14943
rect 19797 14903 19855 14909
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 17954 14832 17960 14884
rect 18012 14872 18018 14884
rect 18294 14875 18352 14881
rect 18294 14872 18306 14875
rect 18012 14844 18306 14872
rect 18012 14832 18018 14844
rect 18294 14841 18306 14844
rect 18340 14841 18352 14875
rect 19812 14872 19840 14903
rect 18294 14835 18352 14841
rect 18432 14844 19840 14872
rect 20809 14875 20867 14881
rect 16080 14776 17632 14804
rect 16080 14764 16086 14776
rect 17862 14764 17868 14816
rect 17920 14804 17926 14816
rect 18432 14804 18460 14844
rect 20809 14841 20821 14875
rect 20855 14841 20867 14875
rect 20809 14835 20867 14841
rect 17920 14776 18460 14804
rect 17920 14764 17926 14776
rect 18690 14764 18696 14816
rect 18748 14804 18754 14816
rect 20824 14804 20852 14835
rect 18748 14776 20852 14804
rect 18748 14764 18754 14776
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1670 14560 1676 14612
rect 1728 14560 1734 14612
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 4154 14600 4160 14612
rect 2823 14572 4160 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 4341 14603 4399 14609
rect 4341 14569 4353 14603
rect 4387 14600 4399 14603
rect 4614 14600 4620 14612
rect 4387 14572 4620 14600
rect 4387 14569 4399 14572
rect 4341 14563 4399 14569
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 4764 14572 4809 14600
rect 4764 14560 4770 14572
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 7009 14603 7067 14609
rect 7009 14600 7021 14603
rect 6972 14572 7021 14600
rect 6972 14560 6978 14572
rect 7009 14569 7021 14572
rect 7055 14569 7067 14603
rect 7009 14563 7067 14569
rect 7285 14603 7343 14609
rect 7285 14569 7297 14603
rect 7331 14600 7343 14603
rect 7331 14572 8524 14600
rect 7331 14569 7343 14572
rect 7285 14563 7343 14569
rect 1688 14532 1716 14560
rect 3326 14532 3332 14544
rect 1688 14504 3332 14532
rect 3326 14492 3332 14504
rect 3384 14492 3390 14544
rect 4801 14535 4859 14541
rect 4801 14501 4813 14535
rect 4847 14532 4859 14535
rect 6086 14532 6092 14544
rect 4847 14504 6092 14532
rect 4847 14501 4859 14504
rect 4801 14495 4859 14501
rect 6086 14492 6092 14504
rect 6144 14492 6150 14544
rect 7098 14492 7104 14544
rect 7156 14532 7162 14544
rect 7156 14504 8432 14532
rect 7156 14492 7162 14504
rect 1670 14424 1676 14476
rect 1728 14464 1734 14476
rect 2133 14467 2191 14473
rect 2133 14464 2145 14467
rect 1728 14436 2145 14464
rect 1728 14424 1734 14436
rect 2133 14433 2145 14436
rect 2179 14433 2191 14467
rect 2133 14427 2191 14433
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14464 3203 14467
rect 3602 14464 3608 14476
rect 3191 14436 3608 14464
rect 3191 14433 3203 14436
rect 3145 14427 3203 14433
rect 3602 14424 3608 14436
rect 3660 14424 3666 14476
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 4028 14436 5365 14464
rect 4028 14424 4034 14436
rect 5353 14433 5365 14436
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 5442 14424 5448 14476
rect 5500 14464 5506 14476
rect 5609 14467 5667 14473
rect 5609 14464 5621 14467
rect 5500 14436 5621 14464
rect 5500 14424 5506 14436
rect 5609 14433 5621 14436
rect 5655 14433 5667 14467
rect 7190 14464 7196 14476
rect 7151 14436 7196 14464
rect 5609 14427 5667 14433
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 7644 14467 7702 14473
rect 7644 14433 7656 14467
rect 7690 14464 7702 14467
rect 8110 14464 8116 14476
rect 7690 14436 8116 14464
rect 7690 14433 7702 14436
rect 7644 14427 7702 14433
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 2222 14396 2228 14408
rect 2183 14368 2228 14396
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 2409 14399 2467 14405
rect 2409 14365 2421 14399
rect 2455 14396 2467 14399
rect 2774 14396 2780 14408
rect 2455 14368 2780 14396
rect 2455 14365 2467 14368
rect 2409 14359 2467 14365
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14365 3295 14399
rect 3418 14396 3424 14408
rect 3379 14368 3424 14396
rect 3237 14359 3295 14365
rect 1765 14331 1823 14337
rect 1765 14297 1777 14331
rect 1811 14328 1823 14331
rect 2958 14328 2964 14340
rect 1811 14300 2964 14328
rect 1811 14297 1823 14300
rect 1765 14291 1823 14297
rect 2958 14288 2964 14300
rect 3016 14288 3022 14340
rect 3252 14328 3280 14359
rect 3418 14356 3424 14368
rect 3476 14356 3482 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 4893 14399 4951 14405
rect 4893 14396 4905 14399
rect 4856 14368 4905 14396
rect 4856 14356 4862 14368
rect 4893 14365 4905 14368
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 7006 14356 7012 14408
rect 7064 14396 7070 14408
rect 7377 14399 7435 14405
rect 7377 14396 7389 14399
rect 7064 14368 7389 14396
rect 7064 14356 7070 14368
rect 7377 14365 7389 14368
rect 7423 14365 7435 14399
rect 8404 14396 8432 14504
rect 8496 14464 8524 14572
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10321 14603 10379 14609
rect 10321 14600 10333 14603
rect 9824 14572 10333 14600
rect 9824 14560 9830 14572
rect 10321 14569 10333 14572
rect 10367 14569 10379 14603
rect 10321 14563 10379 14569
rect 11333 14603 11391 14609
rect 11333 14569 11345 14603
rect 11379 14569 11391 14603
rect 11333 14563 11391 14569
rect 10226 14492 10232 14544
rect 10284 14532 10290 14544
rect 11348 14532 11376 14563
rect 11698 14560 11704 14612
rect 11756 14600 11762 14612
rect 12161 14603 12219 14609
rect 12161 14600 12173 14603
rect 11756 14572 12173 14600
rect 11756 14560 11762 14572
rect 12161 14569 12173 14572
rect 12207 14569 12219 14603
rect 12161 14563 12219 14569
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 13357 14603 13415 14609
rect 13357 14600 13369 14603
rect 12584 14572 13369 14600
rect 12584 14560 12590 14572
rect 13357 14569 13369 14572
rect 13403 14569 13415 14603
rect 13906 14600 13912 14612
rect 13867 14572 13912 14600
rect 13357 14563 13415 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 14737 14603 14795 14609
rect 14737 14569 14749 14603
rect 14783 14600 14795 14603
rect 15102 14600 15108 14612
rect 14783 14572 15108 14600
rect 14783 14569 14795 14572
rect 14737 14563 14795 14569
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14600 15347 14603
rect 17862 14600 17868 14612
rect 15335 14572 17868 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 17954 14560 17960 14612
rect 18012 14600 18018 14612
rect 18417 14603 18475 14609
rect 18417 14600 18429 14603
rect 18012 14572 18429 14600
rect 18012 14560 18018 14572
rect 18417 14569 18429 14572
rect 18463 14569 18475 14603
rect 18874 14600 18880 14612
rect 18835 14572 18880 14600
rect 18417 14563 18475 14569
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 19245 14603 19303 14609
rect 19245 14569 19257 14603
rect 19291 14600 19303 14603
rect 20070 14600 20076 14612
rect 19291 14572 20076 14600
rect 19291 14569 19303 14572
rect 19245 14563 19303 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 16114 14532 16120 14544
rect 10284 14504 11183 14532
rect 11348 14504 16120 14532
rect 10284 14492 10290 14504
rect 11054 14464 11060 14476
rect 8496 14436 11060 14464
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 11155 14464 11183 14504
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 17770 14532 17776 14544
rect 16500 14504 17776 14532
rect 11701 14467 11759 14473
rect 11701 14464 11713 14467
rect 11155 14436 11713 14464
rect 11701 14433 11713 14436
rect 11747 14464 11759 14467
rect 12434 14464 12440 14476
rect 11747 14436 12440 14464
rect 11747 14433 11759 14436
rect 11701 14427 11759 14433
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 13265 14467 13323 14473
rect 13265 14464 13277 14467
rect 13044 14436 13277 14464
rect 13044 14424 13050 14436
rect 13265 14433 13277 14436
rect 13311 14433 13323 14467
rect 14090 14464 14096 14476
rect 14051 14436 14096 14464
rect 13265 14427 13323 14433
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 15654 14464 15660 14476
rect 15615 14436 15660 14464
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 16500 14473 16528 14504
rect 17770 14492 17776 14504
rect 17828 14492 17834 14544
rect 19613 14535 19671 14541
rect 19613 14501 19625 14535
rect 19659 14532 19671 14535
rect 20162 14532 20168 14544
rect 19659 14504 20168 14532
rect 19659 14501 19671 14504
rect 19613 14495 19671 14501
rect 20162 14492 20168 14504
rect 20220 14492 20226 14544
rect 16485 14467 16543 14473
rect 16485 14433 16497 14467
rect 16531 14433 16543 14467
rect 16485 14427 16543 14433
rect 17304 14467 17362 14473
rect 17304 14433 17316 14467
rect 17350 14464 17362 14467
rect 17586 14464 17592 14476
rect 17350 14436 17592 14464
rect 17350 14433 17362 14436
rect 17304 14427 17362 14433
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 18690 14464 18696 14476
rect 18651 14436 18696 14464
rect 18690 14424 18696 14436
rect 18748 14424 18754 14476
rect 20070 14424 20076 14476
rect 20128 14464 20134 14476
rect 20257 14467 20315 14473
rect 20257 14464 20269 14467
rect 20128 14436 20269 14464
rect 20128 14424 20134 14436
rect 20257 14433 20269 14436
rect 20303 14433 20315 14467
rect 20257 14427 20315 14433
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 8404 14368 10425 14396
rect 7377 14359 7435 14365
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 10778 14396 10784 14408
rect 10643 14368 10784 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 10870 14356 10876 14408
rect 10928 14396 10934 14408
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 10928 14368 11805 14396
rect 10928 14356 10934 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14396 12035 14399
rect 12023 14368 12664 14396
rect 12023 14365 12035 14368
rect 11977 14359 12035 14365
rect 7285 14331 7343 14337
rect 7285 14328 7297 14331
rect 3252 14300 3372 14328
rect 3344 14260 3372 14300
rect 6288 14300 7297 14328
rect 3510 14260 3516 14272
rect 3344 14232 3516 14260
rect 3510 14220 3516 14232
rect 3568 14260 3574 14272
rect 6288 14260 6316 14300
rect 7285 14297 7297 14300
rect 7331 14297 7343 14331
rect 7285 14291 7343 14297
rect 12636 14272 12664 14368
rect 12710 14356 12716 14408
rect 12768 14396 12774 14408
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 12768 14368 13461 14396
rect 12768 14356 12774 14368
rect 13449 14365 13461 14368
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 3568 14232 6316 14260
rect 6733 14263 6791 14269
rect 3568 14220 3574 14232
rect 6733 14229 6745 14263
rect 6779 14260 6791 14263
rect 7558 14260 7564 14272
rect 6779 14232 7564 14260
rect 6779 14229 6791 14232
rect 6733 14223 6791 14229
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 8754 14260 8760 14272
rect 8715 14232 8760 14260
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 9953 14263 10011 14269
rect 9953 14229 9965 14263
rect 9999 14260 10011 14263
rect 11974 14260 11980 14272
rect 9999 14232 11980 14260
rect 9999 14229 10011 14232
rect 9953 14223 10011 14229
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12618 14220 12624 14272
rect 12676 14220 12682 14272
rect 12894 14260 12900 14272
rect 12855 14232 12900 14260
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 13464 14260 13492 14359
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 13872 14368 15761 14396
rect 13872 14356 13878 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15470 14288 15476 14340
rect 15528 14328 15534 14340
rect 15856 14328 15884 14359
rect 16022 14356 16028 14408
rect 16080 14396 16086 14408
rect 17037 14399 17095 14405
rect 17037 14396 17049 14399
rect 16080 14368 17049 14396
rect 16080 14356 16086 14368
rect 17037 14365 17049 14368
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19705 14399 19763 14405
rect 19705 14396 19717 14399
rect 19392 14368 19717 14396
rect 19392 14356 19398 14368
rect 19705 14365 19717 14368
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 19794 14356 19800 14408
rect 19852 14396 19858 14408
rect 20901 14399 20959 14405
rect 19852 14368 19897 14396
rect 19852 14356 19858 14368
rect 20901 14365 20913 14399
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 15528 14300 15884 14328
rect 15528 14288 15534 14300
rect 18690 14288 18696 14340
rect 18748 14328 18754 14340
rect 20916 14328 20944 14359
rect 18748 14300 20944 14328
rect 18748 14288 18754 14300
rect 16298 14260 16304 14272
rect 13464 14232 16304 14260
rect 16298 14220 16304 14232
rect 16356 14220 16362 14272
rect 16669 14263 16727 14269
rect 16669 14229 16681 14263
rect 16715 14260 16727 14263
rect 17678 14260 17684 14272
rect 16715 14232 17684 14260
rect 16715 14229 16727 14232
rect 16669 14223 16727 14229
rect 17678 14220 17684 14232
rect 17736 14220 17742 14272
rect 20438 14260 20444 14272
rect 20399 14232 20444 14260
rect 20438 14220 20444 14232
rect 20496 14220 20502 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1670 14056 1676 14068
rect 1631 14028 1676 14056
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 2866 14056 2872 14068
rect 2827 14028 2872 14056
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 6273 14059 6331 14065
rect 6273 14056 6285 14059
rect 5592 14028 6285 14056
rect 5592 14016 5598 14028
rect 6273 14025 6285 14028
rect 6319 14025 6331 14059
rect 6273 14019 6331 14025
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8386 14056 8392 14068
rect 8168 14028 8392 14056
rect 8168 14016 8174 14028
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 9582 14056 9588 14068
rect 9508 14028 9588 14056
rect 4617 13991 4675 13997
rect 4617 13957 4629 13991
rect 4663 13988 4675 13991
rect 4798 13988 4804 14000
rect 4663 13960 4804 13988
rect 4663 13957 4675 13960
rect 4617 13951 4675 13957
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 2314 13920 2320 13932
rect 2275 13892 2320 13920
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 4816 13920 4844 13948
rect 9508 13929 9536 14028
rect 9582 14016 9588 14028
rect 9640 14056 9646 14068
rect 10870 14056 10876 14068
rect 9640 14028 10723 14056
rect 10831 14028 10876 14056
rect 9640 14016 9646 14028
rect 9493 13923 9551 13929
rect 4816 13892 5028 13920
rect 2130 13852 2136 13864
rect 2091 13824 2136 13852
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 2682 13852 2688 13864
rect 2643 13824 2688 13852
rect 2682 13812 2688 13824
rect 2740 13812 2746 13864
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 3970 13852 3976 13864
rect 3283 13824 3976 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 3970 13812 3976 13824
rect 4028 13852 4034 13864
rect 4893 13855 4951 13861
rect 4893 13852 4905 13855
rect 4028 13824 4905 13852
rect 4028 13812 4034 13824
rect 4893 13821 4905 13824
rect 4939 13821 4951 13855
rect 5000 13852 5028 13892
rect 9493 13889 9505 13923
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 5149 13855 5207 13861
rect 5149 13852 5161 13855
rect 5000 13824 5161 13852
rect 4893 13815 4951 13821
rect 5149 13821 5161 13824
rect 5195 13821 5207 13855
rect 7006 13852 7012 13864
rect 6967 13824 7012 13852
rect 5149 13815 5207 13821
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7276 13855 7334 13861
rect 7276 13821 7288 13855
rect 7322 13852 7334 13855
rect 7558 13852 7564 13864
rect 7322 13824 7564 13852
rect 7322 13821 7334 13824
rect 7276 13815 7334 13821
rect 7558 13812 7564 13824
rect 7616 13852 7622 13864
rect 9692 13852 9720 13883
rect 10226 13880 10232 13932
rect 10284 13920 10290 13932
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 10284 13892 10517 13920
rect 10284 13880 10290 13892
rect 10505 13889 10517 13892
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 10612 13852 10640 13883
rect 7616 13824 10640 13852
rect 10695 13852 10723 14028
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 12710 14056 12716 14068
rect 12176 14028 12716 14056
rect 10778 13948 10784 14000
rect 10836 13988 10842 14000
rect 12176 13988 12204 14028
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 15930 14056 15936 14068
rect 13136 14028 15936 14056
rect 13136 14016 13142 14028
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16022 14016 16028 14068
rect 16080 14056 16086 14068
rect 16482 14056 16488 14068
rect 16080 14028 16488 14056
rect 16080 14016 16086 14028
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 16945 14059 17003 14065
rect 16945 14025 16957 14059
rect 16991 14056 17003 14059
rect 17310 14056 17316 14068
rect 16991 14028 17316 14056
rect 16991 14025 17003 14028
rect 16945 14019 17003 14025
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14056 18107 14059
rect 18598 14056 18604 14068
rect 18095 14028 18604 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 19334 14056 19340 14068
rect 19295 14028 19340 14056
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 19978 14016 19984 14068
rect 20036 14016 20042 14068
rect 20162 14016 20168 14068
rect 20220 14056 20226 14068
rect 20349 14059 20407 14065
rect 20349 14056 20361 14059
rect 20220 14028 20361 14056
rect 20220 14016 20226 14028
rect 20349 14025 20361 14028
rect 20395 14025 20407 14059
rect 20349 14019 20407 14025
rect 10836 13960 12204 13988
rect 13817 13991 13875 13997
rect 10836 13948 10842 13960
rect 13817 13957 13829 13991
rect 13863 13988 13875 13991
rect 16040 13988 16068 14016
rect 17126 13988 17132 14000
rect 13863 13960 14044 13988
rect 13863 13957 13875 13960
rect 13817 13951 13875 13957
rect 11422 13920 11428 13932
rect 11383 13892 11428 13920
rect 11422 13880 11428 13892
rect 11480 13920 11486 13932
rect 11698 13920 11704 13932
rect 11480 13892 11704 13920
rect 11480 13880 11486 13892
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 11333 13855 11391 13861
rect 11333 13852 11345 13855
rect 10695 13824 11345 13852
rect 7616 13812 7622 13824
rect 11333 13821 11345 13824
rect 11379 13821 11391 13855
rect 11333 13815 11391 13821
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13852 12495 13855
rect 12526 13852 12532 13864
rect 12483 13824 12532 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 12710 13861 12716 13864
rect 12704 13852 12716 13861
rect 12671 13824 12716 13852
rect 12704 13815 12716 13824
rect 12710 13812 12716 13815
rect 12768 13812 12774 13864
rect 3510 13793 3516 13796
rect 3504 13784 3516 13793
rect 3471 13756 3516 13784
rect 3504 13747 3516 13756
rect 3510 13744 3516 13747
rect 3568 13744 3574 13796
rect 9398 13784 9404 13796
rect 9359 13756 9404 13784
rect 9398 13744 9404 13756
rect 9456 13784 9462 13796
rect 11241 13787 11299 13793
rect 11241 13784 11253 13787
rect 9456 13756 11253 13784
rect 9456 13744 9462 13756
rect 11241 13753 11253 13756
rect 11287 13753 11299 13787
rect 11241 13747 11299 13753
rect 11514 13744 11520 13796
rect 11572 13784 11578 13796
rect 14016 13784 14044 13960
rect 15304 13960 16068 13988
rect 16132 13960 17132 13988
rect 14093 13855 14151 13861
rect 14093 13821 14105 13855
rect 14139 13852 14151 13855
rect 14182 13852 14188 13864
rect 14139 13824 14188 13852
rect 14139 13821 14151 13824
rect 14093 13815 14151 13821
rect 14182 13812 14188 13824
rect 14240 13852 14246 13864
rect 15304 13852 15332 13960
rect 16132 13920 16160 13960
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 17865 13991 17923 13997
rect 17865 13957 17877 13991
rect 17911 13988 17923 13991
rect 19996 13988 20024 14016
rect 17911 13960 20024 13988
rect 17911 13957 17923 13960
rect 17865 13951 17923 13957
rect 16298 13920 16304 13932
rect 16040 13892 16160 13920
rect 16259 13892 16304 13920
rect 14240 13824 15332 13852
rect 14240 13812 14246 13824
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 16040 13852 16068 13892
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 17034 13880 17040 13932
rect 17092 13920 17098 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 17092 13892 17417 13920
rect 17092 13880 17098 13892
rect 17405 13889 17417 13892
rect 17451 13889 17463 13923
rect 17586 13920 17592 13932
rect 17547 13892 17592 13920
rect 17405 13883 17463 13889
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 18524 13929 18552 13960
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 18598 13880 18604 13932
rect 18656 13920 18662 13932
rect 18656 13892 18701 13920
rect 18656 13880 18662 13892
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 19981 13923 20039 13929
rect 19981 13920 19993 13923
rect 19484 13892 19993 13920
rect 19484 13880 19490 13892
rect 19981 13889 19993 13892
rect 20027 13920 20039 13923
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 20027 13892 20913 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 20901 13889 20913 13892
rect 20947 13889 20959 13923
rect 20901 13883 20959 13889
rect 15436 13824 16068 13852
rect 15436 13812 15442 13824
rect 14366 13793 14372 13796
rect 14360 13784 14372 13793
rect 11572 13756 13952 13784
rect 14016 13756 14372 13784
rect 11572 13744 11578 13756
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 2041 13719 2099 13725
rect 2041 13716 2053 13719
rect 1820 13688 2053 13716
rect 1820 13676 1826 13688
rect 2041 13685 2053 13688
rect 2087 13685 2099 13719
rect 9030 13716 9036 13728
rect 8991 13688 9036 13716
rect 2041 13679 2099 13685
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 10042 13716 10048 13728
rect 10003 13688 10048 13716
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 10413 13719 10471 13725
rect 10413 13685 10425 13719
rect 10459 13716 10471 13719
rect 10502 13716 10508 13728
rect 10459 13688 10508 13716
rect 10459 13685 10471 13688
rect 10413 13679 10471 13685
rect 10502 13676 10508 13688
rect 10560 13716 10566 13728
rect 13722 13716 13728 13728
rect 10560 13688 13728 13716
rect 10560 13676 10566 13688
rect 13722 13676 13728 13688
rect 13780 13676 13786 13728
rect 13924 13716 13952 13756
rect 14360 13747 14372 13756
rect 14366 13744 14372 13747
rect 14424 13744 14430 13796
rect 16040 13784 16068 13824
rect 16114 13812 16120 13864
rect 16172 13852 16178 13864
rect 19797 13855 19855 13861
rect 19797 13852 19809 13855
rect 16172 13824 19809 13852
rect 16172 13812 16178 13824
rect 19797 13821 19809 13824
rect 19843 13821 19855 13855
rect 19797 13815 19855 13821
rect 16209 13787 16267 13793
rect 16209 13784 16221 13787
rect 16040 13756 16221 13784
rect 16209 13753 16221 13756
rect 16255 13753 16267 13787
rect 16209 13747 16267 13753
rect 16390 13744 16396 13796
rect 16448 13784 16454 13796
rect 17865 13787 17923 13793
rect 17865 13784 17877 13787
rect 16448 13756 17877 13784
rect 16448 13744 16454 13756
rect 17865 13753 17877 13756
rect 17911 13753 17923 13787
rect 17865 13747 17923 13753
rect 18417 13787 18475 13793
rect 18417 13753 18429 13787
rect 18463 13784 18475 13787
rect 18690 13784 18696 13796
rect 18463 13756 18696 13784
rect 18463 13753 18475 13756
rect 18417 13747 18475 13753
rect 18690 13744 18696 13756
rect 18748 13744 18754 13796
rect 19610 13744 19616 13796
rect 19668 13784 19674 13796
rect 20809 13787 20867 13793
rect 20809 13784 20821 13787
rect 19668 13756 20821 13784
rect 19668 13744 19674 13756
rect 20809 13753 20821 13756
rect 20855 13753 20867 13787
rect 20809 13747 20867 13753
rect 15286 13716 15292 13728
rect 13924 13688 15292 13716
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 15470 13716 15476 13728
rect 15431 13688 15476 13716
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 15746 13716 15752 13728
rect 15707 13688 15752 13716
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 16080 13688 16129 13716
rect 16080 13676 16086 13688
rect 16117 13685 16129 13688
rect 16163 13685 16175 13719
rect 16117 13679 16175 13685
rect 17313 13719 17371 13725
rect 17313 13685 17325 13719
rect 17359 13716 17371 13719
rect 18782 13716 18788 13728
rect 17359 13688 18788 13716
rect 17359 13685 17371 13688
rect 17313 13679 17371 13685
rect 18782 13676 18788 13688
rect 18840 13676 18846 13728
rect 19702 13716 19708 13728
rect 19663 13688 19708 13716
rect 19702 13676 19708 13688
rect 19760 13676 19766 13728
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 20717 13719 20775 13725
rect 20717 13716 20729 13719
rect 20036 13688 20729 13716
rect 20036 13676 20042 13688
rect 20717 13685 20729 13688
rect 20763 13685 20775 13719
rect 20717 13679 20775 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 2222 13512 2228 13524
rect 2183 13484 2228 13512
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 6086 13512 6092 13524
rect 2884 13484 3648 13512
rect 6047 13484 6092 13512
rect 1765 13447 1823 13453
rect 1765 13413 1777 13447
rect 1811 13444 1823 13447
rect 2682 13444 2688 13456
rect 1811 13416 2688 13444
rect 1811 13413 1823 13416
rect 1765 13407 1823 13413
rect 2682 13404 2688 13416
rect 2740 13404 2746 13456
rect 1486 13376 1492 13388
rect 1447 13348 1492 13376
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 2590 13376 2596 13388
rect 2551 13348 2596 13376
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 2884 13376 2912 13484
rect 3142 13404 3148 13456
rect 3200 13444 3206 13456
rect 3513 13447 3571 13453
rect 3513 13444 3525 13447
rect 3200 13416 3525 13444
rect 3200 13404 3206 13416
rect 3513 13413 3525 13416
rect 3559 13413 3571 13447
rect 3620 13444 3648 13484
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 8294 13512 8300 13524
rect 6196 13484 8064 13512
rect 8255 13484 8300 13512
rect 6196 13444 6224 13484
rect 8036 13456 8064 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9030 13512 9036 13524
rect 8803 13484 9036 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 11333 13515 11391 13521
rect 11333 13481 11345 13515
rect 11379 13512 11391 13515
rect 11422 13512 11428 13524
rect 11379 13484 11428 13512
rect 11379 13481 11391 13484
rect 11333 13475 11391 13481
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12676 13484 12817 13512
rect 12676 13472 12682 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 12805 13475 12863 13481
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 13357 13515 13415 13521
rect 13357 13512 13369 13515
rect 12952 13484 13369 13512
rect 12952 13472 12958 13484
rect 13357 13481 13369 13484
rect 13403 13481 13415 13515
rect 13357 13475 13415 13481
rect 14645 13515 14703 13521
rect 14645 13481 14657 13515
rect 14691 13512 14703 13515
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 14691 13484 15485 13512
rect 14691 13481 14703 13484
rect 14645 13475 14703 13481
rect 15473 13481 15485 13484
rect 15519 13481 15531 13515
rect 15841 13515 15899 13521
rect 15841 13512 15853 13515
rect 15473 13475 15531 13481
rect 15672 13484 15853 13512
rect 3620 13416 6224 13444
rect 6549 13447 6607 13453
rect 3513 13407 3571 13413
rect 6549 13413 6561 13447
rect 6595 13444 6607 13447
rect 7098 13444 7104 13456
rect 6595 13416 7104 13444
rect 6595 13413 6607 13416
rect 6549 13407 6607 13413
rect 7098 13404 7104 13416
rect 7156 13404 7162 13456
rect 7558 13404 7564 13456
rect 7616 13404 7622 13456
rect 8018 13404 8024 13456
rect 8076 13404 8082 13456
rect 8665 13447 8723 13453
rect 8665 13413 8677 13447
rect 8711 13444 8723 13447
rect 10042 13444 10048 13456
rect 8711 13416 10048 13444
rect 8711 13413 8723 13416
rect 8665 13407 8723 13413
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 10220 13447 10278 13453
rect 10220 13413 10232 13447
rect 10266 13444 10278 13447
rect 10266 13416 11836 13444
rect 10266 13413 10278 13416
rect 10220 13407 10278 13413
rect 2700 13348 2912 13376
rect 2700 13317 2728 13348
rect 2958 13336 2964 13388
rect 3016 13376 3022 13388
rect 3237 13379 3295 13385
rect 3237 13376 3249 13379
rect 3016 13348 3249 13376
rect 3016 13336 3022 13348
rect 3237 13345 3249 13348
rect 3283 13345 3295 13379
rect 3237 13339 3295 13345
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 4709 13379 4767 13385
rect 4709 13376 4721 13379
rect 4212 13348 4721 13376
rect 4212 13336 4218 13348
rect 4709 13345 4721 13348
rect 4755 13345 4767 13379
rect 4709 13339 4767 13345
rect 4801 13379 4859 13385
rect 4801 13345 4813 13379
rect 4847 13376 4859 13379
rect 4982 13376 4988 13388
rect 4847 13348 4988 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5166 13336 5172 13388
rect 5224 13376 5230 13388
rect 5534 13376 5540 13388
rect 5224 13348 5540 13376
rect 5224 13336 5230 13348
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13376 6515 13379
rect 6914 13376 6920 13388
rect 6503 13348 6920 13376
rect 6503 13345 6515 13348
rect 6457 13339 6515 13345
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 7466 13376 7472 13388
rect 7427 13348 7472 13376
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 7576 13376 7604 13404
rect 7576 13348 7696 13376
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 2777 13311 2835 13317
rect 2777 13277 2789 13311
rect 2823 13277 2835 13311
rect 2777 13271 2835 13277
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13277 4951 13311
rect 6638 13308 6644 13320
rect 6599 13280 6644 13308
rect 4893 13271 4951 13277
rect 2314 13132 2320 13184
rect 2372 13172 2378 13184
rect 2682 13172 2688 13184
rect 2372 13144 2688 13172
rect 2372 13132 2378 13144
rect 2682 13132 2688 13144
rect 2740 13172 2746 13184
rect 2792 13172 2820 13271
rect 4908 13240 4936 13271
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7668 13317 7696 13348
rect 7834 13336 7840 13388
rect 7892 13376 7898 13388
rect 7892 13348 8984 13376
rect 7892 13336 7898 13348
rect 7561 13311 7619 13317
rect 7561 13308 7573 13311
rect 6788 13280 7573 13308
rect 6788 13268 6794 13280
rect 7561 13277 7573 13280
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 8849 13311 8907 13317
rect 8849 13308 8861 13311
rect 8444 13280 8861 13308
rect 8444 13268 8450 13280
rect 8849 13277 8861 13280
rect 8895 13277 8907 13311
rect 8956 13308 8984 13348
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9732 13348 9965 13376
rect 9732 13336 9738 13348
rect 9953 13345 9965 13348
rect 9999 13345 10011 13379
rect 11514 13376 11520 13388
rect 9953 13339 10011 13345
rect 10060 13348 11520 13376
rect 10060 13308 10088 13348
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 11698 13385 11704 13388
rect 11692 13376 11704 13385
rect 11659 13348 11704 13376
rect 11692 13339 11704 13348
rect 11698 13336 11704 13339
rect 11756 13336 11762 13388
rect 11808 13376 11836 13416
rect 11974 13404 11980 13456
rect 12032 13444 12038 13456
rect 13449 13447 13507 13453
rect 13449 13444 13461 13447
rect 12032 13416 13461 13444
rect 12032 13404 12038 13416
rect 13449 13413 13461 13416
rect 13495 13413 13507 13447
rect 13449 13407 13507 13413
rect 14553 13447 14611 13453
rect 14553 13413 14565 13447
rect 14599 13444 14611 13447
rect 15013 13447 15071 13453
rect 15013 13444 15025 13447
rect 14599 13416 15025 13444
rect 14599 13413 14611 13416
rect 14553 13407 14611 13413
rect 15013 13413 15025 13416
rect 15059 13413 15071 13447
rect 15013 13407 15071 13413
rect 15286 13404 15292 13456
rect 15344 13444 15350 13456
rect 15672 13444 15700 13484
rect 15841 13481 15853 13484
rect 15887 13512 15899 13515
rect 16390 13512 16396 13524
rect 15887 13484 16396 13512
rect 15887 13481 15899 13484
rect 15841 13475 15899 13481
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 16482 13472 16488 13524
rect 16540 13512 16546 13524
rect 16540 13484 16804 13512
rect 16540 13472 16546 13484
rect 16574 13444 16580 13456
rect 15344 13416 15700 13444
rect 15764 13416 16580 13444
rect 15344 13404 15350 13416
rect 15764 13376 15792 13416
rect 16574 13404 16580 13416
rect 16632 13404 16638 13456
rect 11808 13348 15792 13376
rect 15933 13379 15991 13385
rect 15933 13345 15945 13379
rect 15979 13376 15991 13379
rect 16666 13376 16672 13388
rect 15979 13348 16672 13376
rect 15979 13345 15991 13348
rect 15933 13339 15991 13345
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 16776 13376 16804 13484
rect 16942 13472 16948 13524
rect 17000 13512 17006 13524
rect 18690 13512 18696 13524
rect 17000 13484 18696 13512
rect 17000 13472 17006 13484
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 19794 13512 19800 13524
rect 18800 13484 19800 13512
rect 16844 13447 16902 13453
rect 16844 13413 16856 13447
rect 16890 13444 16902 13447
rect 18800 13444 18828 13484
rect 19794 13472 19800 13484
rect 19852 13512 19858 13524
rect 19981 13515 20039 13521
rect 19981 13512 19993 13515
rect 19852 13484 19993 13512
rect 19852 13472 19858 13484
rect 19981 13481 19993 13484
rect 20027 13481 20039 13515
rect 20438 13512 20444 13524
rect 20399 13484 20444 13512
rect 19981 13475 20039 13481
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 16890 13416 18828 13444
rect 18868 13447 18926 13453
rect 16890 13413 16902 13416
rect 16844 13407 16902 13413
rect 18868 13413 18880 13447
rect 18914 13444 18926 13447
rect 19426 13444 19432 13456
rect 18914 13416 19432 13444
rect 18914 13413 18926 13416
rect 18868 13407 18926 13413
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 18506 13376 18512 13388
rect 16776 13348 18512 13376
rect 18506 13336 18512 13348
rect 18564 13376 18570 13388
rect 18601 13379 18659 13385
rect 18601 13376 18613 13379
rect 18564 13348 18613 13376
rect 18564 13336 18570 13348
rect 18601 13345 18613 13348
rect 18647 13345 18659 13379
rect 18601 13339 18659 13345
rect 18690 13336 18696 13388
rect 18748 13376 18754 13388
rect 19886 13376 19892 13388
rect 18748 13348 19892 13376
rect 18748 13336 18754 13348
rect 19886 13336 19892 13348
rect 19944 13336 19950 13388
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13376 20315 13379
rect 20806 13376 20812 13388
rect 20303 13348 20812 13376
rect 20303 13345 20315 13348
rect 20257 13339 20315 13345
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 8956 13280 10088 13308
rect 11425 13311 11483 13317
rect 8849 13271 8907 13277
rect 11425 13277 11437 13311
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 5166 13240 5172 13252
rect 4908 13212 5172 13240
rect 5166 13200 5172 13212
rect 5224 13240 5230 13252
rect 6656 13240 6684 13268
rect 5224 13212 6684 13240
rect 5224 13200 5230 13212
rect 8110 13200 8116 13252
rect 8168 13240 8174 13252
rect 9766 13240 9772 13252
rect 8168 13212 9772 13240
rect 8168 13200 8174 13212
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 2740 13144 2820 13172
rect 4341 13175 4399 13181
rect 2740 13132 2746 13144
rect 4341 13141 4353 13175
rect 4387 13172 4399 13175
rect 4706 13172 4712 13184
rect 4387 13144 4712 13172
rect 4387 13141 4399 13144
rect 4341 13135 4399 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 5718 13132 5724 13184
rect 5776 13172 5782 13184
rect 6638 13172 6644 13184
rect 5776 13144 6644 13172
rect 5776 13132 5782 13144
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 7101 13175 7159 13181
rect 7101 13141 7113 13175
rect 7147 13172 7159 13175
rect 8294 13172 8300 13184
rect 7147 13144 8300 13172
rect 7147 13141 7159 13144
rect 7101 13135 7159 13141
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 11440 13172 11468 13271
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 13354 13308 13360 13320
rect 12676 13280 13360 13308
rect 12676 13268 12682 13280
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 13633 13311 13691 13317
rect 13633 13277 13645 13311
rect 13679 13308 13691 13311
rect 14366 13308 14372 13320
rect 13679 13280 14372 13308
rect 13679 13277 13691 13280
rect 13633 13271 13691 13277
rect 14366 13268 14372 13280
rect 14424 13308 14430 13320
rect 14737 13311 14795 13317
rect 14737 13308 14749 13311
rect 14424 13280 14749 13308
rect 14424 13268 14430 13280
rect 14737 13277 14749 13280
rect 14783 13277 14795 13311
rect 14737 13271 14795 13277
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13308 15071 13311
rect 15746 13308 15752 13320
rect 15059 13280 15752 13308
rect 15059 13277 15071 13280
rect 15013 13271 15071 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13308 16175 13311
rect 16298 13308 16304 13320
rect 16163 13280 16304 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 16482 13268 16488 13320
rect 16540 13308 16546 13320
rect 16577 13311 16635 13317
rect 16577 13308 16589 13311
rect 16540 13280 16589 13308
rect 16540 13268 16546 13280
rect 16577 13277 16589 13280
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 12989 13243 13047 13249
rect 12989 13209 13001 13243
rect 13035 13240 13047 13243
rect 13814 13240 13820 13252
rect 13035 13212 13820 13240
rect 13035 13209 13047 13212
rect 12989 13203 13047 13209
rect 13814 13200 13820 13212
rect 13872 13200 13878 13252
rect 14185 13243 14243 13249
rect 14185 13209 14197 13243
rect 14231 13240 14243 13243
rect 15654 13240 15660 13252
rect 14231 13212 15660 13240
rect 14231 13209 14243 13212
rect 14185 13203 14243 13209
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 12526 13172 12532 13184
rect 11440 13144 12532 13172
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 12710 13132 12716 13184
rect 12768 13172 12774 13184
rect 16114 13172 16120 13184
rect 12768 13144 16120 13172
rect 12768 13132 12774 13144
rect 16114 13132 16120 13144
rect 16172 13132 16178 13184
rect 16316 13172 16344 13268
rect 17957 13175 18015 13181
rect 17957 13172 17969 13175
rect 16316 13144 17969 13172
rect 17957 13141 17969 13144
rect 18003 13141 18015 13175
rect 17957 13135 18015 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1854 12968 1860 12980
rect 1815 12940 1860 12968
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 3605 12971 3663 12977
rect 3605 12968 3617 12971
rect 3568 12940 3617 12968
rect 3568 12928 3574 12940
rect 3605 12937 3617 12940
rect 3651 12968 3663 12971
rect 5166 12968 5172 12980
rect 3651 12940 5172 12968
rect 3651 12937 3663 12940
rect 3605 12931 3663 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7800 12940 7941 12968
rect 7800 12928 7806 12940
rect 7929 12937 7941 12940
rect 7975 12937 7987 12971
rect 7929 12931 7987 12937
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 8941 12971 8999 12977
rect 8941 12968 8953 12971
rect 8076 12940 8953 12968
rect 8076 12928 8082 12940
rect 8941 12937 8953 12940
rect 8987 12937 8999 12971
rect 8941 12931 8999 12937
rect 12621 12971 12679 12977
rect 12621 12937 12633 12971
rect 12667 12968 12679 12971
rect 14090 12968 14096 12980
rect 12667 12940 14096 12968
rect 12667 12937 12679 12940
rect 12621 12931 12679 12937
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 15654 12928 15660 12980
rect 15712 12968 15718 12980
rect 15749 12971 15807 12977
rect 15749 12968 15761 12971
rect 15712 12940 15761 12968
rect 15712 12928 15718 12940
rect 15749 12937 15761 12940
rect 15795 12937 15807 12971
rect 15749 12931 15807 12937
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 16172 12940 17785 12968
rect 16172 12928 16178 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 17862 12928 17868 12980
rect 17920 12968 17926 12980
rect 19426 12968 19432 12980
rect 17920 12940 19012 12968
rect 19387 12940 19432 12968
rect 17920 12928 17926 12940
rect 6917 12903 6975 12909
rect 6917 12869 6929 12903
rect 6963 12900 6975 12903
rect 12989 12903 13047 12909
rect 6963 12872 7687 12900
rect 6963 12869 6975 12872
rect 6917 12863 6975 12869
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 2225 12835 2283 12841
rect 2225 12832 2237 12835
rect 1636 12804 2237 12832
rect 1636 12792 1642 12804
rect 2225 12801 2237 12804
rect 2271 12801 2283 12835
rect 4154 12832 4160 12844
rect 4115 12804 4160 12832
rect 2225 12795 2283 12801
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 5166 12832 5172 12844
rect 5127 12804 5172 12832
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6604 12804 7389 12832
rect 6604 12792 6610 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7558 12832 7564 12844
rect 7519 12804 7564 12832
rect 7377 12795 7435 12801
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12733 1731 12767
rect 1673 12727 1731 12733
rect 2492 12767 2550 12773
rect 2492 12733 2504 12767
rect 2538 12764 2550 12767
rect 2774 12764 2780 12776
rect 2538 12736 2780 12764
rect 2538 12733 2550 12736
rect 2492 12727 2550 12733
rect 1688 12696 1716 12727
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 5994 12724 6000 12776
rect 6052 12764 6058 12776
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 6052 12736 7297 12764
rect 6052 12724 6058 12736
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 7392 12764 7420 12795
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 7659 12832 7687 12872
rect 12989 12869 13001 12903
rect 13035 12900 13047 12903
rect 14366 12900 14372 12912
rect 13035 12872 14372 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 15838 12860 15844 12912
rect 15896 12900 15902 12912
rect 16390 12900 16396 12912
rect 15896 12872 16396 12900
rect 15896 12860 15902 12872
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 16945 12903 17003 12909
rect 16945 12869 16957 12903
rect 16991 12900 17003 12903
rect 17954 12900 17960 12912
rect 16991 12872 17960 12900
rect 16991 12869 17003 12872
rect 16945 12863 17003 12869
rect 17954 12860 17960 12872
rect 18012 12860 18018 12912
rect 18984 12900 19012 12940
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19978 12968 19984 12980
rect 19939 12940 19984 12968
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 18984 12872 20484 12900
rect 7659 12804 7972 12832
rect 7834 12764 7840 12776
rect 7392 12736 7840 12764
rect 7285 12727 7343 12733
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 3142 12696 3148 12708
rect 1688 12668 3148 12696
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 4985 12699 5043 12705
rect 4985 12665 4997 12699
rect 5031 12696 5043 12699
rect 5166 12696 5172 12708
rect 5031 12668 5172 12696
rect 5031 12665 5043 12668
rect 4985 12659 5043 12665
rect 5166 12656 5172 12668
rect 5224 12656 5230 12708
rect 7944 12696 7972 12804
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8481 12835 8539 12841
rect 8481 12832 8493 12835
rect 8444 12804 8493 12832
rect 8444 12792 8450 12804
rect 8481 12801 8493 12804
rect 8527 12801 8539 12835
rect 8481 12795 8539 12801
rect 8662 12792 8668 12844
rect 8720 12832 8726 12844
rect 9493 12835 9551 12841
rect 9493 12832 9505 12835
rect 8720 12804 9505 12832
rect 8720 12792 8726 12804
rect 9493 12801 9505 12804
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 9582 12792 9588 12844
rect 9640 12832 9646 12844
rect 13446 12832 13452 12844
rect 9640 12804 13452 12832
rect 9640 12792 9646 12804
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 13630 12832 13636 12844
rect 13591 12804 13636 12832
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 16022 12832 16028 12844
rect 15983 12804 16028 12832
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 17494 12832 17500 12844
rect 16632 12804 17500 12832
rect 16632 12792 16638 12804
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 17773 12835 17831 12841
rect 17773 12801 17785 12835
rect 17819 12832 17831 12835
rect 17819 12804 18184 12832
rect 17819 12801 17831 12804
rect 17773 12795 17831 12801
rect 8294 12764 8300 12776
rect 8255 12736 8300 12764
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 12161 12767 12219 12773
rect 9355 12736 10916 12764
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 8389 12699 8447 12705
rect 8389 12696 8401 12699
rect 7944 12668 8401 12696
rect 8389 12665 8401 12668
rect 8435 12665 8447 12699
rect 10226 12696 10232 12708
rect 8389 12659 8447 12665
rect 9324 12668 10232 12696
rect 4614 12628 4620 12640
rect 4575 12600 4620 12628
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 5077 12631 5135 12637
rect 5077 12597 5089 12631
rect 5123 12628 5135 12631
rect 5534 12628 5540 12640
rect 5123 12600 5540 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 5534 12588 5540 12600
rect 5592 12628 5598 12640
rect 9324 12628 9352 12668
rect 10226 12656 10232 12668
rect 10284 12656 10290 12708
rect 10321 12699 10379 12705
rect 10321 12665 10333 12699
rect 10367 12696 10379 12699
rect 10410 12696 10416 12708
rect 10367 12668 10416 12696
rect 10367 12665 10379 12668
rect 10321 12659 10379 12665
rect 10410 12656 10416 12668
rect 10468 12656 10474 12708
rect 10888 12696 10916 12736
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12207 12736 12817 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14240 12736 14381 12764
rect 14240 12724 14246 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 14636 12767 14694 12773
rect 14636 12733 14648 12767
rect 14682 12764 14694 12767
rect 15470 12764 15476 12776
rect 14682 12736 15476 12764
rect 14682 12733 14694 12736
rect 14636 12727 14694 12733
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 16298 12724 16304 12776
rect 16356 12764 16362 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 16356 12736 18061 12764
rect 16356 12724 16362 12736
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18156 12764 18184 12804
rect 20346 12792 20352 12844
rect 20404 12792 20410 12844
rect 20456 12841 20484 12872
rect 20441 12835 20499 12841
rect 20441 12801 20453 12835
rect 20487 12801 20499 12835
rect 20441 12795 20499 12801
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 18305 12767 18363 12773
rect 18305 12764 18317 12767
rect 18156 12736 18317 12764
rect 18049 12727 18107 12733
rect 18305 12733 18317 12736
rect 18351 12764 18363 12767
rect 20364 12764 20392 12792
rect 20548 12764 20576 12795
rect 18351 12736 18552 12764
rect 18351 12733 18363 12736
rect 18305 12727 18363 12733
rect 12618 12696 12624 12708
rect 10888 12668 12624 12696
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 13078 12656 13084 12708
rect 13136 12696 13142 12708
rect 13449 12699 13507 12705
rect 13449 12696 13461 12699
rect 13136 12668 13461 12696
rect 13136 12656 13142 12668
rect 13449 12665 13461 12668
rect 13495 12665 13507 12699
rect 13449 12659 13507 12665
rect 13722 12656 13728 12708
rect 13780 12696 13786 12708
rect 16942 12696 16948 12708
rect 13780 12668 16948 12696
rect 13780 12656 13786 12668
rect 16942 12656 16948 12668
rect 17000 12656 17006 12708
rect 17313 12699 17371 12705
rect 17313 12665 17325 12699
rect 17359 12696 17371 12699
rect 18414 12696 18420 12708
rect 17359 12668 18420 12696
rect 17359 12665 17371 12668
rect 17313 12659 17371 12665
rect 18414 12656 18420 12668
rect 18472 12656 18478 12708
rect 18524 12696 18552 12736
rect 20272 12736 20576 12764
rect 20272 12696 20300 12736
rect 18524 12668 20300 12696
rect 20349 12699 20407 12705
rect 20349 12665 20361 12699
rect 20395 12696 20407 12699
rect 20898 12696 20904 12708
rect 20395 12668 20904 12696
rect 20395 12665 20407 12668
rect 20349 12659 20407 12665
rect 20898 12656 20904 12668
rect 20956 12656 20962 12708
rect 5592 12600 9352 12628
rect 9401 12631 9459 12637
rect 5592 12588 5598 12600
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 9674 12628 9680 12640
rect 9447 12600 9680 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11609 12631 11667 12637
rect 11609 12628 11621 12631
rect 11204 12600 11621 12628
rect 11204 12588 11210 12600
rect 11609 12597 11621 12600
rect 11655 12628 11667 12631
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 11655 12600 12173 12628
rect 11655 12597 11667 12600
rect 11609 12591 11667 12597
rect 12161 12597 12173 12600
rect 12207 12597 12219 12631
rect 13354 12628 13360 12640
rect 13315 12600 13360 12628
rect 12161 12591 12219 12597
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 17405 12631 17463 12637
rect 17405 12597 17417 12631
rect 17451 12628 17463 12631
rect 19242 12628 19248 12640
rect 17451 12600 19248 12628
rect 17451 12597 17463 12600
rect 17405 12591 17463 12597
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 2869 12427 2927 12433
rect 2869 12424 2881 12427
rect 2832 12396 2881 12424
rect 2832 12384 2838 12396
rect 2869 12393 2881 12396
rect 2915 12393 2927 12427
rect 4246 12424 4252 12436
rect 4207 12396 4252 12424
rect 2869 12387 2927 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 4617 12427 4675 12433
rect 4617 12393 4629 12427
rect 4663 12424 4675 12427
rect 4706 12424 4712 12436
rect 4663 12396 4712 12424
rect 4663 12393 4675 12396
rect 4617 12387 4675 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 5258 12424 5264 12436
rect 5040 12396 5264 12424
rect 5040 12384 5046 12396
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 9493 12427 9551 12433
rect 9493 12424 9505 12427
rect 7432 12396 9505 12424
rect 7432 12384 7438 12396
rect 9493 12393 9505 12396
rect 9539 12393 9551 12427
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9493 12387 9551 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 10045 12427 10103 12433
rect 10045 12424 10057 12427
rect 10008 12396 10057 12424
rect 10008 12384 10014 12396
rect 10045 12393 10057 12396
rect 10091 12393 10103 12427
rect 10045 12387 10103 12393
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 13078 12424 13084 12436
rect 12851 12396 13084 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13446 12384 13452 12436
rect 13504 12424 13510 12436
rect 14645 12427 14703 12433
rect 14645 12424 14657 12427
rect 13504 12396 14657 12424
rect 13504 12384 13510 12396
rect 14645 12393 14657 12396
rect 14691 12424 14703 12427
rect 16206 12424 16212 12436
rect 14691 12396 16212 12424
rect 14691 12393 14703 12396
rect 14645 12387 14703 12393
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 17681 12427 17739 12433
rect 17681 12424 17693 12427
rect 17552 12396 17693 12424
rect 17552 12384 17558 12396
rect 17681 12393 17693 12396
rect 17727 12393 17739 12427
rect 17681 12387 17739 12393
rect 17770 12384 17776 12436
rect 17828 12424 17834 12436
rect 17828 12396 19380 12424
rect 17828 12384 17834 12396
rect 1756 12359 1814 12365
rect 1756 12325 1768 12359
rect 1802 12356 1814 12359
rect 2682 12356 2688 12368
rect 1802 12328 2688 12356
rect 1802 12325 1814 12328
rect 1756 12319 1814 12325
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 15378 12356 15384 12368
rect 4120 12328 15384 12356
rect 4120 12316 4126 12328
rect 15378 12316 15384 12328
rect 15436 12316 15442 12368
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 17218 12356 17224 12368
rect 17092 12328 17224 12356
rect 17092 12316 17098 12328
rect 17218 12316 17224 12328
rect 17276 12356 17282 12368
rect 17862 12356 17868 12368
rect 17276 12328 17868 12356
rect 17276 12316 17282 12328
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 18417 12359 18475 12365
rect 18417 12325 18429 12359
rect 18463 12356 18475 12359
rect 18506 12356 18512 12368
rect 18463 12328 18512 12356
rect 18463 12325 18475 12328
rect 18417 12319 18475 12325
rect 18506 12316 18512 12328
rect 18564 12316 18570 12368
rect 19352 12365 19380 12396
rect 19610 12384 19616 12436
rect 19668 12424 19674 12436
rect 19797 12427 19855 12433
rect 19797 12424 19809 12427
rect 19668 12396 19809 12424
rect 19668 12384 19674 12396
rect 19797 12393 19809 12396
rect 19843 12393 19855 12427
rect 19797 12387 19855 12393
rect 20165 12427 20223 12433
rect 20165 12393 20177 12427
rect 20211 12424 20223 12427
rect 20714 12424 20720 12436
rect 20211 12396 20720 12424
rect 20211 12393 20223 12396
rect 20165 12387 20223 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 20898 12424 20904 12436
rect 20859 12396 20904 12424
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 19337 12359 19395 12365
rect 19337 12325 19349 12359
rect 19383 12325 19395 12359
rect 19337 12319 19395 12325
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12288 1547 12291
rect 1578 12288 1584 12300
rect 1535 12260 1584 12288
rect 1535 12257 1547 12260
rect 1489 12251 1547 12257
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 4709 12291 4767 12297
rect 4709 12288 4721 12291
rect 4672 12260 4721 12288
rect 4672 12248 4678 12260
rect 4709 12257 4721 12260
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 5885 12291 5943 12297
rect 5885 12288 5897 12291
rect 5776 12260 5897 12288
rect 5776 12248 5782 12260
rect 5885 12257 5897 12260
rect 5931 12257 5943 12291
rect 5885 12251 5943 12257
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 7064 12260 7297 12288
rect 7064 12248 7070 12260
rect 7285 12257 7297 12260
rect 7331 12257 7343 12291
rect 7552 12291 7610 12297
rect 7552 12288 7564 12291
rect 7285 12251 7343 12257
rect 7392 12260 7564 12288
rect 4798 12220 4804 12232
rect 4759 12192 4804 12220
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12189 5687 12223
rect 7392 12220 7420 12260
rect 7552 12257 7564 12260
rect 7598 12288 7610 12291
rect 7598 12260 8800 12288
rect 7598 12257 7610 12260
rect 7552 12251 7610 12257
rect 5629 12183 5687 12189
rect 7024 12192 7420 12220
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 5644 12152 5672 12183
rect 7024 12161 7052 12192
rect 4212 12124 5672 12152
rect 7009 12155 7067 12161
rect 4212 12112 4218 12124
rect 7009 12121 7021 12155
rect 7055 12121 7067 12155
rect 8662 12152 8668 12164
rect 8623 12124 8668 12152
rect 7009 12115 7067 12121
rect 8662 12112 8668 12124
rect 8720 12112 8726 12164
rect 8772 12152 8800 12260
rect 10778 12248 10784 12300
rect 10836 12288 10842 12300
rect 11140 12291 11198 12297
rect 11140 12288 11152 12291
rect 10836 12260 11152 12288
rect 10836 12248 10842 12260
rect 11140 12257 11152 12260
rect 11186 12288 11198 12291
rect 12713 12291 12771 12297
rect 12713 12288 12725 12291
rect 11186 12260 12725 12288
rect 11186 12257 11198 12260
rect 11140 12251 11198 12257
rect 12713 12257 12725 12260
rect 12759 12257 12771 12291
rect 12713 12251 12771 12257
rect 13173 12291 13231 12297
rect 13173 12257 13185 12291
rect 13219 12288 13231 12291
rect 13906 12288 13912 12300
rect 13219 12260 13912 12288
rect 13219 12257 13231 12260
rect 13173 12251 13231 12257
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14001 12291 14059 12297
rect 14001 12257 14013 12291
rect 14047 12288 14059 12291
rect 14090 12288 14096 12300
rect 14047 12260 14096 12288
rect 14047 12257 14059 12260
rect 14001 12251 14059 12257
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 14553 12291 14611 12297
rect 14553 12257 14565 12291
rect 14599 12288 14611 12291
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 14599 12260 15301 12288
rect 14599 12257 14611 12260
rect 14553 12251 14611 12257
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 16568 12291 16626 12297
rect 16568 12257 16580 12291
rect 16614 12288 16626 12291
rect 17126 12288 17132 12300
rect 16614 12260 17132 12288
rect 16614 12257 16626 12260
rect 16568 12251 16626 12257
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17954 12248 17960 12300
rect 18012 12288 18018 12300
rect 18325 12291 18383 12297
rect 18325 12288 18337 12291
rect 18012 12260 18337 12288
rect 18012 12248 18018 12260
rect 18325 12257 18337 12260
rect 18371 12257 18383 12291
rect 18325 12251 18383 12257
rect 19061 12291 19119 12297
rect 19061 12257 19073 12291
rect 19107 12257 19119 12291
rect 19061 12251 19119 12257
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12220 9551 12223
rect 9950 12220 9956 12232
rect 9539 12192 9956 12220
rect 9539 12189 9551 12192
rect 9493 12183 9551 12189
rect 9950 12180 9956 12192
rect 10008 12220 10014 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10008 12192 10149 12220
rect 10008 12180 10014 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10244 12152 10272 12183
rect 10502 12180 10508 12232
rect 10560 12220 10566 12232
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10560 12192 10885 12220
rect 10560 12180 10566 12192
rect 10873 12189 10885 12192
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 11940 12192 13277 12220
rect 11940 12180 11946 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 14182 12220 14188 12232
rect 13495 12192 14188 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 8772 12124 10272 12152
rect 12253 12155 12311 12161
rect 12253 12121 12265 12155
rect 12299 12152 12311 12155
rect 13464 12152 13492 12183
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 14642 12152 14648 12164
rect 12299 12124 13492 12152
rect 13740 12124 14648 12152
rect 12299 12121 12311 12124
rect 12253 12115 12311 12121
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 12434 12084 12440 12096
rect 4120 12056 12440 12084
rect 4120 12044 4126 12056
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12713 12087 12771 12093
rect 12713 12053 12725 12087
rect 12759 12084 12771 12087
rect 13740 12084 13768 12124
rect 14642 12112 14648 12124
rect 14700 12152 14706 12164
rect 14752 12152 14780 12183
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 16298 12220 16304 12232
rect 15804 12192 16304 12220
rect 15804 12180 15810 12192
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 18598 12220 18604 12232
rect 18559 12192 18604 12220
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 19076 12152 19104 12251
rect 20162 12180 20168 12232
rect 20220 12220 20226 12232
rect 20257 12223 20315 12229
rect 20257 12220 20269 12223
rect 20220 12192 20269 12220
rect 20220 12180 20226 12192
rect 20257 12189 20269 12192
rect 20303 12189 20315 12223
rect 20438 12220 20444 12232
rect 20399 12192 20444 12220
rect 20257 12183 20315 12189
rect 20438 12180 20444 12192
rect 20496 12180 20502 12232
rect 14700 12124 14780 12152
rect 17236 12124 19104 12152
rect 14700 12112 14706 12124
rect 12759 12056 13768 12084
rect 13817 12087 13875 12093
rect 12759 12053 12771 12056
rect 12713 12047 12771 12053
rect 13817 12053 13829 12087
rect 13863 12084 13875 12087
rect 13906 12084 13912 12096
rect 13863 12056 13912 12084
rect 13863 12053 13875 12056
rect 13817 12047 13875 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 14185 12087 14243 12093
rect 14185 12084 14197 12087
rect 14056 12056 14197 12084
rect 14056 12044 14062 12056
rect 14185 12053 14197 12056
rect 14231 12053 14243 12087
rect 14185 12047 14243 12053
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 17236 12084 17264 12124
rect 14424 12056 17264 12084
rect 17957 12087 18015 12093
rect 14424 12044 14430 12056
rect 17957 12053 17969 12087
rect 18003 12084 18015 12087
rect 19518 12084 19524 12096
rect 18003 12056 19524 12084
rect 18003 12053 18015 12056
rect 17957 12047 18015 12053
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1486 11840 1492 11892
rect 1544 11880 1550 11892
rect 2317 11883 2375 11889
rect 2317 11880 2329 11883
rect 1544 11852 2329 11880
rect 1544 11840 1550 11852
rect 2317 11849 2329 11852
rect 2363 11849 2375 11883
rect 5718 11880 5724 11892
rect 2317 11843 2375 11849
rect 2976 11852 5724 11880
rect 2976 11753 3004 11852
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7837 11883 7895 11889
rect 7837 11880 7849 11883
rect 7248 11852 7849 11880
rect 7248 11840 7254 11852
rect 7837 11849 7849 11852
rect 7883 11849 7895 11883
rect 10137 11883 10195 11889
rect 7837 11843 7895 11849
rect 8220 11852 10088 11880
rect 3326 11772 3332 11824
rect 3384 11812 3390 11824
rect 4154 11812 4160 11824
rect 3384 11784 4160 11812
rect 3384 11772 3390 11784
rect 4154 11772 4160 11784
rect 4212 11812 4218 11824
rect 4212 11784 4384 11812
rect 4212 11772 4218 11784
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 2961 11707 3019 11713
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 4246 11744 4252 11756
rect 4019 11716 4252 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 4356 11753 4384 11784
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 8220 11812 8248 11852
rect 7708 11784 8248 11812
rect 10060 11812 10088 11852
rect 10137 11849 10149 11883
rect 10183 11880 10195 11883
rect 11882 11880 11888 11892
rect 10183 11852 11888 11880
rect 10183 11849 10195 11852
rect 10137 11843 10195 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12492 11852 13400 11880
rect 12492 11840 12498 11852
rect 10870 11812 10876 11824
rect 10060 11784 10876 11812
rect 7708 11772 7714 11784
rect 10870 11772 10876 11784
rect 10928 11772 10934 11824
rect 13372 11812 13400 11852
rect 13630 11840 13636 11892
rect 13688 11880 13694 11892
rect 13817 11883 13875 11889
rect 13817 11880 13829 11883
rect 13688 11852 13829 11880
rect 13688 11840 13694 11852
rect 13817 11849 13829 11852
rect 13863 11849 13875 11883
rect 14090 11880 14096 11892
rect 14051 11852 14096 11880
rect 13817 11843 13875 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 17034 11880 17040 11892
rect 14476 11852 17040 11880
rect 13372 11784 13584 11812
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 7009 11747 7067 11753
rect 7009 11713 7021 11747
rect 7055 11744 7067 11747
rect 7466 11744 7472 11756
rect 7055 11716 7472 11744
rect 7055 11713 7067 11716
rect 7009 11707 7067 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 9950 11704 9956 11756
rect 10008 11744 10014 11756
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10008 11716 10609 11744
rect 10008 11704 10014 11716
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10778 11744 10784 11756
rect 10739 11716 10784 11744
rect 10597 11707 10655 11713
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 11882 11744 11888 11756
rect 11843 11716 11888 11744
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 13556 11744 13584 11784
rect 14476 11744 14504 11852
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 17126 11840 17132 11892
rect 17184 11880 17190 11892
rect 18969 11883 19027 11889
rect 18969 11880 18981 11883
rect 17184 11852 18981 11880
rect 17184 11840 17190 11852
rect 18969 11849 18981 11852
rect 19015 11849 19027 11883
rect 19150 11880 19156 11892
rect 19111 11852 19156 11880
rect 18969 11843 19027 11849
rect 19150 11840 19156 11852
rect 19208 11840 19214 11892
rect 19702 11840 19708 11892
rect 19760 11880 19766 11892
rect 20165 11883 20223 11889
rect 20165 11880 20177 11883
rect 19760 11852 20177 11880
rect 19760 11840 19766 11852
rect 20165 11849 20177 11852
rect 20211 11849 20223 11883
rect 20165 11843 20223 11849
rect 16117 11815 16175 11821
rect 16117 11781 16129 11815
rect 16163 11812 16175 11815
rect 19978 11812 19984 11824
rect 16163 11784 19984 11812
rect 16163 11781 16175 11784
rect 16117 11775 16175 11781
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 14642 11744 14648 11756
rect 13556 11716 14504 11744
rect 14603 11716 14648 11744
rect 14642 11704 14648 11716
rect 14700 11744 14706 11756
rect 15654 11744 15660 11756
rect 14700 11716 15660 11744
rect 14700 11704 14706 11716
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 16080 11716 16681 11744
rect 16080 11704 16086 11716
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 16758 11704 16764 11756
rect 16816 11744 16822 11756
rect 17405 11747 17463 11753
rect 17405 11744 17417 11747
rect 16816 11716 17417 11744
rect 16816 11704 16822 11716
rect 17405 11713 17417 11716
rect 17451 11713 17463 11747
rect 17405 11707 17463 11713
rect 18230 11704 18236 11756
rect 18288 11744 18294 11756
rect 18598 11744 18604 11756
rect 18288 11716 18604 11744
rect 18288 11704 18294 11716
rect 18598 11704 18604 11716
rect 18656 11744 18662 11756
rect 18693 11747 18751 11753
rect 18693 11744 18705 11747
rect 18656 11716 18705 11744
rect 18656 11704 18662 11716
rect 18693 11713 18705 11716
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11744 19027 11747
rect 19702 11744 19708 11756
rect 19015 11716 19708 11744
rect 19015 11713 19027 11716
rect 18969 11707 19027 11713
rect 19702 11704 19708 11716
rect 19760 11704 19766 11756
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 20496 11716 20729 11744
rect 20496 11704 20502 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 2498 11636 2504 11688
rect 2556 11676 2562 11688
rect 8021 11679 8079 11685
rect 2556 11648 4292 11676
rect 2556 11636 2562 11648
rect 2685 11611 2743 11617
rect 2685 11577 2697 11611
rect 2731 11608 2743 11611
rect 2731 11580 3372 11608
rect 2731 11577 2743 11580
rect 2685 11571 2743 11577
rect 1486 11540 1492 11552
rect 1447 11512 1492 11540
rect 1486 11500 1492 11512
rect 1544 11500 1550 11552
rect 2777 11543 2835 11549
rect 2777 11509 2789 11543
rect 2823 11540 2835 11543
rect 2958 11540 2964 11552
rect 2823 11512 2964 11540
rect 2823 11509 2835 11512
rect 2777 11503 2835 11509
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 3344 11549 3372 11580
rect 3329 11543 3387 11549
rect 3329 11509 3341 11543
rect 3375 11509 3387 11543
rect 3694 11540 3700 11552
rect 3655 11512 3700 11540
rect 3329 11503 3387 11509
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 3789 11543 3847 11549
rect 3789 11509 3801 11543
rect 3835 11540 3847 11543
rect 4062 11540 4068 11552
rect 3835 11512 4068 11540
rect 3835 11509 3847 11512
rect 3789 11503 3847 11509
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 4264 11540 4292 11648
rect 8021 11645 8033 11679
rect 8067 11645 8079 11679
rect 8202 11676 8208 11688
rect 8163 11648 8208 11676
rect 8021 11639 8079 11645
rect 4338 11568 4344 11620
rect 4396 11608 4402 11620
rect 4608 11611 4666 11617
rect 4608 11608 4620 11611
rect 4396 11580 4620 11608
rect 4396 11568 4402 11580
rect 4608 11577 4620 11580
rect 4654 11608 4666 11611
rect 4798 11608 4804 11620
rect 4654 11580 4804 11608
rect 4654 11577 4666 11580
rect 4608 11571 4666 11577
rect 4798 11568 4804 11580
rect 4856 11568 4862 11620
rect 5074 11568 5080 11620
rect 5132 11608 5138 11620
rect 6730 11608 6736 11620
rect 5132 11580 6736 11608
rect 5132 11568 5138 11580
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 8036 11608 8064 11639
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8472 11679 8530 11685
rect 8472 11645 8484 11679
rect 8518 11676 8530 11679
rect 8754 11676 8760 11688
rect 8518 11648 8760 11676
rect 8518 11645 8530 11648
rect 8472 11639 8530 11645
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 10042 11636 10048 11688
rect 10100 11676 10106 11688
rect 10505 11679 10563 11685
rect 10505 11676 10517 11679
rect 10100 11648 10517 11676
rect 10100 11636 10106 11648
rect 10505 11645 10517 11648
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 12250 11676 12256 11688
rect 11848 11648 12256 11676
rect 11848 11636 11854 11648
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 12400 11648 12449 11676
rect 12400 11636 12406 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 14461 11679 14519 11685
rect 14461 11645 14473 11679
rect 14507 11676 14519 11679
rect 15010 11676 15016 11688
rect 14507 11648 15016 11676
rect 14507 11645 14519 11648
rect 14461 11639 14519 11645
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 15252 11648 17233 11676
rect 15252 11636 15258 11648
rect 17221 11645 17233 11648
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 18509 11679 18567 11685
rect 18509 11645 18521 11679
rect 18555 11676 18567 11679
rect 19334 11676 19340 11688
rect 18555 11648 19340 11676
rect 18555 11645 18567 11648
rect 18509 11639 18567 11645
rect 19334 11636 19340 11648
rect 19392 11636 19398 11688
rect 19518 11676 19524 11688
rect 19479 11648 19524 11676
rect 19518 11636 19524 11648
rect 19576 11636 19582 11688
rect 11146 11608 11152 11620
rect 8036 11580 11152 11608
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 11514 11608 11520 11620
rect 11348 11580 11520 11608
rect 8662 11540 8668 11552
rect 4264 11512 8668 11540
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 11348 11549 11376 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 11701 11611 11759 11617
rect 11701 11577 11713 11611
rect 11747 11608 11759 11611
rect 12704 11611 12762 11617
rect 11747 11580 12296 11608
rect 11747 11577 11759 11580
rect 11701 11571 11759 11577
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9364 11512 9597 11540
rect 9364 11500 9370 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 11333 11543 11391 11549
rect 11333 11509 11345 11543
rect 11379 11509 11391 11543
rect 11790 11540 11796 11552
rect 11751 11512 11796 11540
rect 11333 11503 11391 11509
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12268 11540 12296 11580
rect 12704 11577 12716 11611
rect 12750 11608 12762 11611
rect 14182 11608 14188 11620
rect 12750 11580 14188 11608
rect 12750 11577 12762 11580
rect 12704 11571 12762 11577
rect 14182 11568 14188 11580
rect 14240 11568 14246 11620
rect 14553 11611 14611 11617
rect 14553 11608 14565 11611
rect 14292 11580 14565 11608
rect 12342 11540 12348 11552
rect 12268 11512 12348 11540
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 12618 11500 12624 11552
rect 12676 11540 12682 11552
rect 14292 11540 14320 11580
rect 14553 11577 14565 11580
rect 14599 11577 14611 11611
rect 14553 11571 14611 11577
rect 14642 11568 14648 11620
rect 14700 11608 14706 11620
rect 16577 11611 16635 11617
rect 16577 11608 16589 11611
rect 14700 11580 16589 11608
rect 14700 11568 14706 11580
rect 16577 11577 16589 11580
rect 16623 11577 16635 11611
rect 16577 11571 16635 11577
rect 16942 11568 16948 11620
rect 17000 11608 17006 11620
rect 17862 11608 17868 11620
rect 17000 11580 17868 11608
rect 17000 11568 17006 11580
rect 17862 11568 17868 11580
rect 17920 11568 17926 11620
rect 19613 11611 19671 11617
rect 19613 11608 19625 11611
rect 18156 11580 19625 11608
rect 15102 11540 15108 11552
rect 12676 11512 14320 11540
rect 15063 11512 15108 11540
rect 12676 11500 12682 11512
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15470 11540 15476 11552
rect 15431 11512 15476 11540
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 15565 11543 15623 11549
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 16298 11540 16304 11552
rect 15611 11512 16304 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16482 11540 16488 11552
rect 16443 11512 16488 11540
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 18156 11549 18184 11580
rect 19613 11577 19625 11580
rect 19659 11577 19671 11611
rect 20625 11611 20683 11617
rect 20625 11608 20637 11611
rect 19613 11571 19671 11577
rect 19720 11580 20637 11608
rect 18141 11543 18199 11549
rect 18141 11509 18153 11543
rect 18187 11509 18199 11543
rect 18141 11503 18199 11509
rect 18601 11543 18659 11549
rect 18601 11509 18613 11543
rect 18647 11540 18659 11543
rect 18690 11540 18696 11552
rect 18647 11512 18696 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 19720 11540 19748 11580
rect 20625 11577 20637 11580
rect 20671 11577 20683 11611
rect 20625 11571 20683 11577
rect 19576 11512 19748 11540
rect 19576 11500 19582 11512
rect 19886 11500 19892 11552
rect 19944 11540 19950 11552
rect 20533 11543 20591 11549
rect 20533 11540 20545 11543
rect 19944 11512 20545 11540
rect 19944 11500 19950 11512
rect 20533 11509 20545 11512
rect 20579 11509 20591 11543
rect 20533 11503 20591 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2590 11336 2596 11348
rect 1995 11308 2596 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 2958 11336 2964 11348
rect 2919 11308 2964 11336
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 4062 11336 4068 11348
rect 4023 11308 4068 11336
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 5537 11339 5595 11345
rect 5537 11305 5549 11339
rect 5583 11336 5595 11339
rect 5626 11336 5632 11348
rect 5583 11308 5632 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6641 11339 6699 11345
rect 6641 11305 6653 11339
rect 6687 11336 6699 11339
rect 8205 11339 8263 11345
rect 8205 11336 8217 11339
rect 6687 11308 8217 11336
rect 6687 11305 6699 11308
rect 6641 11299 6699 11305
rect 8205 11305 8217 11308
rect 8251 11305 8263 11339
rect 8205 11299 8263 11305
rect 10045 11339 10103 11345
rect 10045 11305 10057 11339
rect 10091 11336 10103 11339
rect 10226 11336 10232 11348
rect 10091 11308 10232 11336
rect 10091 11305 10103 11308
rect 10045 11299 10103 11305
rect 10226 11296 10232 11308
rect 10284 11336 10290 11348
rect 10594 11336 10600 11348
rect 10284 11308 10600 11336
rect 10284 11296 10290 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11149 11339 11207 11345
rect 11149 11336 11161 11339
rect 10928 11308 11161 11336
rect 10928 11296 10934 11308
rect 11149 11305 11161 11308
rect 11195 11305 11207 11339
rect 11149 11299 11207 11305
rect 11701 11339 11759 11345
rect 11701 11305 11713 11339
rect 11747 11336 11759 11339
rect 11790 11336 11796 11348
rect 11747 11308 11796 11336
rect 11747 11305 11759 11308
rect 11701 11299 11759 11305
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 16390 11336 16396 11348
rect 12268 11308 16396 11336
rect 2038 11228 2044 11280
rect 2096 11268 2102 11280
rect 2317 11271 2375 11277
rect 2317 11268 2329 11271
rect 2096 11240 2329 11268
rect 2096 11228 2102 11240
rect 2317 11237 2329 11240
rect 2363 11237 2375 11271
rect 2317 11231 2375 11237
rect 2406 11228 2412 11280
rect 2464 11268 2470 11280
rect 3329 11271 3387 11277
rect 2464 11240 2509 11268
rect 2464 11228 2470 11240
rect 3329 11237 3341 11271
rect 3375 11268 3387 11271
rect 3881 11271 3939 11277
rect 3881 11268 3893 11271
rect 3375 11240 3893 11268
rect 3375 11237 3387 11240
rect 3329 11231 3387 11237
rect 3881 11237 3893 11240
rect 3927 11237 3939 11271
rect 12268 11268 12296 11308
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 17126 11336 17132 11348
rect 17087 11308 17132 11336
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 17681 11339 17739 11345
rect 17681 11305 17693 11339
rect 17727 11305 17739 11339
rect 18690 11336 18696 11348
rect 17681 11299 17739 11305
rect 18064 11308 18348 11336
rect 18651 11308 18696 11336
rect 3881 11231 3939 11237
rect 4172 11240 12296 11268
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11200 1915 11203
rect 2424 11200 2452 11228
rect 4172 11200 4200 11240
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 12526 11268 12532 11280
rect 12400 11240 12532 11268
rect 12400 11228 12406 11240
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 12980 11271 13038 11277
rect 12980 11237 12992 11271
rect 13026 11268 13038 11271
rect 13630 11268 13636 11280
rect 13026 11240 13636 11268
rect 13026 11237 13038 11240
rect 12980 11231 13038 11237
rect 13630 11228 13636 11240
rect 13688 11228 13694 11280
rect 17696 11268 17724 11299
rect 18064 11268 18092 11308
rect 17696 11240 18092 11268
rect 18141 11271 18199 11277
rect 18141 11237 18153 11271
rect 18187 11268 18199 11271
rect 18320 11268 18348 11308
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 19150 11336 19156 11348
rect 19111 11308 19156 11336
rect 19150 11296 19156 11308
rect 19208 11296 19214 11348
rect 19242 11296 19248 11348
rect 19300 11336 19306 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 19300 11308 19717 11336
rect 19300 11296 19306 11308
rect 19705 11305 19717 11308
rect 19751 11305 19763 11339
rect 19705 11299 19763 11305
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20165 11339 20223 11345
rect 20165 11336 20177 11339
rect 20036 11308 20177 11336
rect 20036 11296 20042 11308
rect 20165 11305 20177 11308
rect 20211 11305 20223 11339
rect 20165 11299 20223 11305
rect 20073 11271 20131 11277
rect 20073 11268 20085 11271
rect 18187 11240 18276 11268
rect 18320 11240 20085 11268
rect 18187 11237 18199 11240
rect 18141 11231 18199 11237
rect 1903 11172 4200 11200
rect 1903 11169 1915 11172
rect 1857 11163 1915 11169
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4304 11172 4445 11200
rect 4304 11160 4310 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 4706 11200 4712 11212
rect 4571 11172 4712 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5442 11200 5448 11212
rect 5403 11172 5448 11200
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6546 11200 6552 11212
rect 6507 11172 6552 11200
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 7558 11200 7564 11212
rect 7519 11172 7564 11200
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 8478 11200 8484 11212
rect 7699 11172 8484 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 8573 11203 8631 11209
rect 8573 11169 8585 11203
rect 8619 11200 8631 11203
rect 10042 11200 10048 11212
rect 8619 11172 10048 11200
rect 8619 11169 8631 11172
rect 8573 11163 8631 11169
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10318 11200 10324 11212
rect 10192 11172 10324 11200
rect 10192 11160 10198 11172
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 10686 11200 10692 11212
rect 10428 11172 10692 11200
rect 2498 11132 2504 11144
rect 2459 11104 2504 11132
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11101 3479 11135
rect 3421 11095 3479 11101
rect 3605 11135 3663 11141
rect 3605 11101 3617 11135
rect 3651 11132 3663 11135
rect 4338 11132 4344 11144
rect 3651 11104 4344 11132
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 3436 11064 3464 11095
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 4982 11132 4988 11144
rect 4663 11104 4988 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4982 11092 4988 11104
rect 5040 11132 5046 11144
rect 5721 11135 5779 11141
rect 5721 11132 5733 11135
rect 5040 11104 5733 11132
rect 5040 11092 5046 11104
rect 5721 11101 5733 11104
rect 5767 11132 5779 11135
rect 6730 11132 6736 11144
rect 5767 11104 6736 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 7745 11135 7803 11141
rect 7745 11132 7757 11135
rect 7524 11104 7757 11132
rect 7524 11092 7530 11104
rect 7745 11101 7757 11104
rect 7791 11101 7803 11135
rect 7745 11095 7803 11101
rect 8665 11135 8723 11141
rect 8665 11101 8677 11135
rect 8711 11101 8723 11135
rect 8665 11095 8723 11101
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11101 8815 11135
rect 8757 11095 8815 11101
rect 6181 11067 6239 11073
rect 6181 11064 6193 11067
rect 3436 11036 6193 11064
rect 6181 11033 6193 11036
rect 6227 11033 6239 11067
rect 6181 11027 6239 11033
rect 6822 11024 6828 11076
rect 6880 11064 6886 11076
rect 7193 11067 7251 11073
rect 7193 11064 7205 11067
rect 6880 11036 7205 11064
rect 6880 11024 6886 11036
rect 7193 11033 7205 11036
rect 7239 11033 7251 11067
rect 7193 11027 7251 11033
rect 7650 11024 7656 11076
rect 7708 11064 7714 11076
rect 8680 11064 8708 11095
rect 7708 11036 8708 11064
rect 7708 11024 7714 11036
rect 3881 10999 3939 11005
rect 3881 10965 3893 10999
rect 3927 10996 3939 10999
rect 5077 10999 5135 11005
rect 5077 10996 5089 10999
rect 3927 10968 5089 10996
rect 3927 10965 3939 10968
rect 3881 10959 3939 10965
rect 5077 10965 5089 10968
rect 5123 10965 5135 10999
rect 5077 10959 5135 10965
rect 6270 10956 6276 11008
rect 6328 10996 6334 11008
rect 8772 10996 8800 11095
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 9364 11104 10241 11132
rect 9364 11092 9370 11104
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 10042 11024 10048 11076
rect 10100 11064 10106 11076
rect 10428 11064 10456 11172
rect 10686 11160 10692 11172
rect 10744 11200 10750 11212
rect 11057 11203 11115 11209
rect 11057 11200 11069 11203
rect 10744 11172 11069 11200
rect 10744 11160 10750 11172
rect 11057 11169 11069 11172
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 12069 11203 12127 11209
rect 12069 11169 12081 11203
rect 12115 11200 12127 11203
rect 12618 11200 12624 11212
rect 12115 11172 12624 11200
rect 12115 11169 12127 11172
rect 12069 11163 12127 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 13964 11172 15669 11200
rect 13964 11160 13970 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11200 15807 11203
rect 15838 11200 15844 11212
rect 15795 11172 15844 11200
rect 15795 11169 15807 11172
rect 15749 11163 15807 11169
rect 11330 11132 11336 11144
rect 11291 11104 11336 11132
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11101 12219 11135
rect 12342 11132 12348 11144
rect 12303 11104 12348 11132
rect 12161 11095 12219 11101
rect 10100 11036 10456 11064
rect 10689 11067 10747 11073
rect 10100 11024 10106 11036
rect 10689 11033 10701 11067
rect 10735 11064 10747 11067
rect 12176 11064 12204 11095
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12434 11092 12440 11144
rect 12492 11092 12498 11144
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 15764 11132 15792 11163
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 16022 11209 16028 11212
rect 16016 11200 16028 11209
rect 15983 11172 16028 11200
rect 16016 11163 16028 11172
rect 16022 11160 16028 11163
rect 16080 11160 16086 11212
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11169 18107 11203
rect 18248 11200 18276 11240
rect 20073 11237 20085 11240
rect 20119 11237 20131 11271
rect 20073 11231 20131 11237
rect 18598 11200 18604 11212
rect 18248 11172 18604 11200
rect 18049 11163 18107 11169
rect 15427 11104 15792 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 12452 11064 12480 11092
rect 12728 11064 12756 11095
rect 14090 11064 14096 11076
rect 10735 11036 12204 11064
rect 12360 11036 12756 11064
rect 14051 11036 14096 11064
rect 10735 11033 10747 11036
rect 10689 11027 10747 11033
rect 6328 10968 8800 10996
rect 9677 10999 9735 11005
rect 6328 10956 6334 10968
rect 9677 10965 9689 10999
rect 9723 10996 9735 10999
rect 10134 10996 10140 11008
rect 9723 10968 10140 10996
rect 9723 10965 9735 10968
rect 9677 10959 9735 10965
rect 10134 10956 10140 10968
rect 10192 10956 10198 11008
rect 10502 10956 10508 11008
rect 10560 10996 10566 11008
rect 12360 10996 12388 11036
rect 14090 11024 14096 11036
rect 14148 11024 14154 11076
rect 18064 11064 18092 11163
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 18690 11160 18696 11212
rect 18748 11200 18754 11212
rect 19061 11203 19119 11209
rect 19061 11200 19073 11203
rect 18748 11172 19073 11200
rect 18748 11160 18754 11172
rect 19061 11169 19073 11172
rect 19107 11200 19119 11203
rect 19610 11200 19616 11212
rect 19107 11172 19616 11200
rect 19107 11169 19119 11172
rect 19061 11163 19119 11169
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 18230 11132 18236 11144
rect 18191 11104 18236 11132
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 19242 11132 19248 11144
rect 19203 11104 19248 11132
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 19702 11092 19708 11144
rect 19760 11132 19766 11144
rect 20257 11135 20315 11141
rect 20257 11132 20269 11135
rect 19760 11104 20269 11132
rect 19760 11092 19766 11104
rect 20257 11101 20269 11104
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 19058 11064 19064 11076
rect 15304 11036 15608 11064
rect 18064 11036 19064 11064
rect 10560 10968 12388 10996
rect 10560 10956 10566 10968
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 15304 10996 15332 11036
rect 12492 10968 15332 10996
rect 15381 10999 15439 11005
rect 12492 10956 12498 10968
rect 15381 10965 15393 10999
rect 15427 10996 15439 10999
rect 15473 10999 15531 11005
rect 15473 10996 15485 10999
rect 15427 10968 15485 10996
rect 15427 10965 15439 10968
rect 15381 10959 15439 10965
rect 15473 10965 15485 10968
rect 15519 10965 15531 10999
rect 15580 10996 15608 11036
rect 19058 11024 19064 11036
rect 19116 11024 19122 11076
rect 17310 10996 17316 11008
rect 15580 10968 17316 10996
rect 15473 10959 15531 10965
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 2682 10752 2688 10804
rect 2740 10792 2746 10804
rect 2869 10795 2927 10801
rect 2869 10792 2881 10795
rect 2740 10764 2881 10792
rect 2740 10752 2746 10764
rect 2869 10761 2881 10764
rect 2915 10761 2927 10795
rect 2869 10755 2927 10761
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 4798 10792 4804 10804
rect 3384 10764 4384 10792
rect 4759 10764 4804 10792
rect 3384 10752 3390 10764
rect 4356 10724 4384 10764
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5721 10795 5779 10801
rect 5721 10761 5733 10795
rect 5767 10792 5779 10795
rect 6546 10792 6552 10804
rect 5767 10764 6552 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 7558 10792 7564 10804
rect 7519 10764 7564 10792
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 12618 10792 12624 10804
rect 8128 10764 11560 10792
rect 12579 10764 12624 10792
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 4356 10696 5089 10724
rect 5077 10693 5089 10696
rect 5123 10693 5135 10727
rect 7006 10724 7012 10736
rect 5077 10687 5135 10693
rect 5276 10696 7012 10724
rect 1489 10591 1547 10597
rect 1489 10557 1501 10591
rect 1535 10588 1547 10591
rect 1578 10588 1584 10600
rect 1535 10560 1584 10588
rect 1535 10557 1547 10560
rect 1489 10551 1547 10557
rect 1578 10548 1584 10560
rect 1636 10548 1642 10600
rect 1756 10591 1814 10597
rect 1756 10557 1768 10591
rect 1802 10588 1814 10591
rect 2498 10588 2504 10600
rect 1802 10560 2504 10588
rect 1802 10557 1814 10560
rect 1756 10551 1814 10557
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10557 3479 10591
rect 3688 10591 3746 10597
rect 3688 10588 3700 10591
rect 3421 10551 3479 10557
rect 3620 10560 3700 10588
rect 1596 10520 1624 10548
rect 3326 10520 3332 10532
rect 1596 10492 3332 10520
rect 3326 10480 3332 10492
rect 3384 10520 3390 10532
rect 3436 10520 3464 10551
rect 3620 10532 3648 10560
rect 3688 10557 3700 10560
rect 3734 10588 3746 10591
rect 4982 10588 4988 10600
rect 3734 10560 4988 10588
rect 3734 10557 3746 10560
rect 3688 10551 3746 10557
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 5276 10597 5304 10696
rect 7006 10684 7012 10696
rect 7064 10684 7070 10736
rect 6270 10656 6276 10668
rect 6231 10628 6276 10656
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10656 6883 10659
rect 8128 10656 8156 10764
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 9582 10724 9588 10736
rect 8536 10696 9588 10724
rect 8536 10684 8542 10696
rect 9582 10684 9588 10696
rect 9640 10684 9646 10736
rect 6871 10628 8156 10656
rect 8205 10659 8263 10665
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 8205 10625 8217 10659
rect 8251 10656 8263 10659
rect 8294 10656 8300 10668
rect 8251 10628 8300 10656
rect 8251 10625 8263 10628
rect 8205 10619 8263 10625
rect 8294 10616 8300 10628
rect 8352 10616 8358 10668
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 9364 10628 10057 10656
rect 9364 10616 9370 10628
rect 10045 10625 10057 10628
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6362 10588 6368 10600
rect 6135 10560 6368 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 7190 10588 7196 10600
rect 7151 10560 7196 10588
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10588 7987 10591
rect 8478 10588 8484 10600
rect 7975 10560 8484 10588
rect 7975 10557 7987 10560
rect 7929 10551 7987 10557
rect 8478 10548 8484 10560
rect 8536 10548 8542 10600
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10588 9919 10591
rect 9950 10588 9956 10600
rect 9907 10560 9956 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 10502 10588 10508 10600
rect 10463 10560 10508 10588
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 11532 10588 11560 10764
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 13354 10752 13360 10804
rect 13412 10792 13418 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 13412 10764 13645 10792
rect 13412 10752 13418 10764
rect 13633 10761 13645 10764
rect 13679 10761 13691 10795
rect 16022 10792 16028 10804
rect 15983 10764 16028 10792
rect 13633 10755 13691 10761
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 16301 10795 16359 10801
rect 16301 10761 16313 10795
rect 16347 10792 16359 10795
rect 16482 10792 16488 10804
rect 16347 10764 16488 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 18598 10792 18604 10804
rect 18559 10764 18604 10792
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19392 10764 19625 10792
rect 19392 10752 19398 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 19702 10752 19708 10804
rect 19760 10792 19766 10804
rect 20254 10792 20260 10804
rect 19760 10764 20260 10792
rect 19760 10752 19766 10764
rect 20254 10752 20260 10764
rect 20312 10752 20318 10804
rect 11698 10684 11704 10736
rect 11756 10724 11762 10736
rect 12434 10724 12440 10736
rect 11756 10696 12440 10724
rect 11756 10684 11762 10696
rect 12434 10684 12440 10696
rect 12492 10684 12498 10736
rect 13262 10656 13268 10668
rect 13223 10628 13268 10656
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 14182 10656 14188 10668
rect 14143 10628 14188 10656
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 11532 10560 13093 10588
rect 13081 10557 13093 10560
rect 13127 10588 13139 10591
rect 13170 10588 13176 10600
rect 13127 10560 13176 10588
rect 13127 10557 13139 10560
rect 13081 10551 13139 10557
rect 13170 10548 13176 10560
rect 13228 10548 13234 10600
rect 13998 10588 14004 10600
rect 13959 10560 14004 10588
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 14645 10591 14703 10597
rect 14645 10588 14657 10591
rect 14608 10560 14657 10588
rect 14608 10548 14614 10560
rect 14645 10557 14657 10560
rect 14691 10557 14703 10591
rect 16761 10591 16819 10597
rect 16761 10588 16773 10591
rect 14645 10551 14703 10557
rect 14752 10560 16773 10588
rect 3384 10492 3464 10520
rect 3384 10480 3390 10492
rect 3602 10480 3608 10532
rect 3660 10480 3666 10532
rect 4062 10480 4068 10532
rect 4120 10520 4126 10532
rect 10594 10520 10600 10532
rect 4120 10492 10600 10520
rect 4120 10480 4126 10492
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 10772 10523 10830 10529
rect 10772 10489 10784 10523
rect 10818 10520 10830 10523
rect 11146 10520 11152 10532
rect 10818 10492 11152 10520
rect 10818 10489 10830 10492
rect 10772 10483 10830 10489
rect 11146 10480 11152 10492
rect 11204 10480 11210 10532
rect 14752 10520 14780 10560
rect 16761 10557 16773 10560
rect 16807 10557 16819 10591
rect 16761 10551 16819 10557
rect 11716 10492 14780 10520
rect 14912 10523 14970 10529
rect 6181 10455 6239 10461
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6227 10424 6837 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 6825 10415 6883 10421
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 8021 10455 8079 10461
rect 8021 10452 8033 10455
rect 7156 10424 8033 10452
rect 7156 10412 7162 10424
rect 8021 10421 8033 10424
rect 8067 10421 8079 10455
rect 9490 10452 9496 10464
rect 9451 10424 9496 10452
rect 8021 10415 8079 10421
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 9953 10455 10011 10461
rect 9953 10452 9965 10455
rect 9916 10424 9965 10452
rect 9916 10412 9922 10424
rect 9953 10421 9965 10424
rect 9999 10452 10011 10455
rect 11716 10452 11744 10492
rect 14912 10489 14924 10523
rect 14958 10520 14970 10523
rect 15010 10520 15016 10532
rect 14958 10492 15016 10520
rect 14958 10489 14970 10492
rect 14912 10483 14970 10489
rect 15010 10480 15016 10492
rect 15068 10520 15074 10532
rect 16868 10520 16896 10619
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 18012 10628 18061 10656
rect 18012 10616 18018 10628
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 18598 10616 18604 10668
rect 18656 10656 18662 10668
rect 19150 10656 19156 10668
rect 18656 10628 19012 10656
rect 19111 10628 19156 10656
rect 18656 10616 18662 10628
rect 17034 10548 17040 10600
rect 17092 10588 17098 10600
rect 18690 10588 18696 10600
rect 17092 10560 18696 10588
rect 17092 10548 17098 10560
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 18984 10597 19012 10628
rect 19150 10616 19156 10628
rect 19208 10656 19214 10668
rect 20165 10659 20223 10665
rect 20165 10656 20177 10659
rect 19208 10628 20177 10656
rect 19208 10616 19214 10628
rect 20165 10625 20177 10628
rect 20211 10625 20223 10659
rect 20806 10656 20812 10668
rect 20767 10628 20812 10656
rect 20165 10619 20223 10625
rect 20806 10616 20812 10628
rect 20864 10616 20870 10668
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10557 19027 10591
rect 18969 10551 19027 10557
rect 19242 10548 19248 10600
rect 19300 10588 19306 10600
rect 19610 10588 19616 10600
rect 19300 10560 19616 10588
rect 19300 10548 19306 10560
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 20622 10588 20628 10600
rect 20583 10560 20628 10588
rect 20622 10548 20628 10560
rect 20680 10548 20686 10600
rect 17494 10520 17500 10532
rect 15068 10492 17500 10520
rect 15068 10480 15074 10492
rect 17494 10480 17500 10492
rect 17552 10480 17558 10532
rect 19518 10520 19524 10532
rect 18616 10492 19524 10520
rect 11882 10452 11888 10464
rect 9999 10424 11744 10452
rect 11795 10424 11888 10452
rect 9999 10421 10011 10424
rect 9953 10415 10011 10421
rect 11882 10412 11888 10424
rect 11940 10452 11946 10464
rect 12342 10452 12348 10464
rect 11940 10424 12348 10452
rect 11940 10412 11946 10424
rect 12342 10412 12348 10424
rect 12400 10412 12406 10464
rect 12989 10455 13047 10461
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 13998 10452 14004 10464
rect 13035 10424 14004 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14093 10455 14151 10461
rect 14093 10421 14105 10455
rect 14139 10452 14151 10455
rect 15102 10452 15108 10464
rect 14139 10424 15108 10452
rect 14139 10421 14151 10424
rect 14093 10415 14151 10421
rect 15102 10412 15108 10424
rect 15160 10412 15166 10464
rect 16669 10455 16727 10461
rect 16669 10421 16681 10455
rect 16715 10452 16727 10455
rect 18616 10452 18644 10492
rect 19518 10480 19524 10492
rect 19576 10480 19582 10532
rect 19981 10523 20039 10529
rect 19981 10489 19993 10523
rect 20027 10520 20039 10523
rect 20162 10520 20168 10532
rect 20027 10492 20168 10520
rect 20027 10489 20039 10492
rect 19981 10483 20039 10489
rect 20162 10480 20168 10492
rect 20220 10480 20226 10532
rect 20254 10480 20260 10532
rect 20312 10520 20318 10532
rect 20990 10520 20996 10532
rect 20312 10492 20996 10520
rect 20312 10480 20318 10492
rect 20990 10480 20996 10492
rect 21048 10480 21054 10532
rect 18690 10452 18696 10464
rect 16715 10424 18696 10452
rect 16715 10421 16727 10424
rect 16669 10415 16727 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 19061 10455 19119 10461
rect 19061 10421 19073 10455
rect 19107 10452 19119 10455
rect 19334 10452 19340 10464
rect 19107 10424 19340 10452
rect 19107 10421 19119 10424
rect 19061 10415 19119 10421
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 20073 10455 20131 10461
rect 20073 10421 20085 10455
rect 20119 10452 20131 10455
rect 20346 10452 20352 10464
rect 20119 10424 20352 10452
rect 20119 10421 20131 10424
rect 20073 10415 20131 10421
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2130 10248 2136 10260
rect 1995 10220 2136 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 2961 10251 3019 10257
rect 2961 10217 2973 10251
rect 3007 10248 3019 10251
rect 3694 10248 3700 10260
rect 3007 10220 3700 10248
rect 3007 10217 3019 10220
rect 2961 10211 3019 10217
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 5442 10248 5448 10260
rect 4663 10220 5448 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 5537 10251 5595 10257
rect 5537 10217 5549 10251
rect 5583 10248 5595 10251
rect 5994 10248 6000 10260
rect 5583 10220 6000 10248
rect 5583 10217 5595 10220
rect 5537 10211 5595 10217
rect 5994 10208 6000 10220
rect 6052 10248 6058 10260
rect 6178 10248 6184 10260
rect 6052 10220 6184 10248
rect 6052 10208 6058 10220
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6788 10220 7021 10248
rect 6788 10208 6794 10220
rect 7009 10217 7021 10220
rect 7055 10217 7067 10251
rect 7009 10211 7067 10217
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 9309 10251 9367 10257
rect 9309 10248 9321 10251
rect 7524 10220 9321 10248
rect 7524 10208 7530 10220
rect 9309 10217 9321 10220
rect 9355 10217 9367 10251
rect 9309 10211 9367 10217
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 9548 10220 10057 10248
rect 9548 10208 9554 10220
rect 10045 10217 10057 10220
rect 10091 10217 10103 10251
rect 10045 10211 10103 10217
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 12066 10248 12072 10260
rect 10192 10220 10237 10248
rect 10336 10220 12072 10248
rect 10192 10208 10198 10220
rect 2409 10183 2467 10189
rect 2409 10149 2421 10183
rect 2455 10180 2467 10183
rect 2774 10180 2780 10192
rect 2455 10152 2780 10180
rect 2455 10149 2467 10152
rect 2409 10143 2467 10149
rect 2774 10140 2780 10152
rect 2832 10140 2838 10192
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 8196 10183 8254 10189
rect 4120 10152 7972 10180
rect 4120 10140 4126 10152
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10112 2375 10115
rect 3329 10115 3387 10121
rect 2363 10084 3280 10112
rect 2363 10081 2375 10084
rect 2317 10075 2375 10081
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 1581 9979 1639 9985
rect 1581 9945 1593 9979
rect 1627 9976 1639 9979
rect 2866 9976 2872 9988
rect 1627 9948 2872 9976
rect 1627 9945 1639 9948
rect 1581 9939 1639 9945
rect 2866 9936 2872 9948
rect 2924 9936 2930 9988
rect 3252 9908 3280 10084
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 4157 10115 4215 10121
rect 4157 10112 4169 10115
rect 3375 10084 4169 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 4157 10081 4169 10084
rect 4203 10081 4215 10115
rect 4157 10075 4215 10081
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10112 5043 10115
rect 5896 10115 5954 10121
rect 5896 10112 5908 10115
rect 5031 10084 5212 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3602 10044 3608 10056
rect 3563 10016 3608 10044
rect 3421 10007 3479 10013
rect 3436 9976 3464 10007
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 3694 10004 3700 10056
rect 3752 10044 3758 10056
rect 5074 10044 5080 10056
rect 3752 10016 5080 10044
rect 3752 10004 3758 10016
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 4154 9976 4160 9988
rect 3436 9948 4160 9976
rect 4154 9936 4160 9948
rect 4212 9936 4218 9988
rect 5184 9976 5212 10084
rect 5276 10084 5908 10112
rect 5276 10053 5304 10084
rect 5896 10081 5908 10084
rect 5942 10112 5954 10115
rect 6270 10112 6276 10124
rect 5942 10084 6276 10112
rect 5942 10081 5954 10084
rect 5896 10075 5954 10081
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 7064 10084 7849 10112
rect 7064 10072 7070 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 7944 10112 7972 10152
rect 8196 10149 8208 10183
rect 8242 10180 8254 10183
rect 8294 10180 8300 10192
rect 8242 10152 8300 10180
rect 8242 10149 8254 10152
rect 8196 10143 8254 10149
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 9950 10140 9956 10192
rect 10008 10180 10014 10192
rect 10336 10180 10364 10220
rect 10008 10152 10364 10180
rect 11140 10183 11198 10189
rect 10008 10140 10014 10152
rect 11140 10149 11152 10183
rect 11186 10180 11198 10183
rect 11882 10180 11888 10192
rect 11186 10152 11888 10180
rect 11186 10149 11198 10152
rect 11140 10143 11198 10149
rect 11882 10140 11888 10152
rect 11940 10140 11946 10192
rect 11698 10112 11704 10124
rect 7944 10084 11704 10112
rect 7837 10075 7895 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11992 10112 12020 10220
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 17494 10248 17500 10260
rect 17455 10220 17500 10248
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 17770 10208 17776 10260
rect 17828 10248 17834 10260
rect 17865 10251 17923 10257
rect 17865 10248 17877 10251
rect 17828 10220 17877 10248
rect 17828 10208 17834 10220
rect 17865 10217 17877 10220
rect 17911 10217 17923 10251
rect 17865 10211 17923 10217
rect 18049 10251 18107 10257
rect 18049 10217 18061 10251
rect 18095 10248 18107 10251
rect 18506 10248 18512 10260
rect 18095 10220 18512 10248
rect 18095 10217 18107 10220
rect 18049 10211 18107 10217
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19245 10251 19303 10257
rect 19245 10248 19257 10251
rect 19116 10220 19257 10248
rect 19116 10208 19122 10220
rect 19245 10217 19257 10220
rect 19291 10217 19303 10251
rect 19245 10211 19303 10217
rect 13722 10180 13728 10192
rect 13683 10152 13728 10180
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 13817 10183 13875 10189
rect 13817 10149 13829 10183
rect 13863 10180 13875 10183
rect 15746 10180 15752 10192
rect 13863 10152 15752 10180
rect 13863 10149 13875 10152
rect 13817 10143 13875 10149
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 16384 10183 16442 10189
rect 16384 10149 16396 10183
rect 16430 10180 16442 10183
rect 16574 10180 16580 10192
rect 16430 10152 16580 10180
rect 16430 10149 16442 10152
rect 16384 10143 16442 10149
rect 16574 10140 16580 10152
rect 16632 10140 16638 10192
rect 16850 10140 16856 10192
rect 16908 10180 16914 10192
rect 17310 10180 17316 10192
rect 16908 10152 17316 10180
rect 16908 10140 16914 10152
rect 17310 10140 17316 10152
rect 17368 10140 17374 10192
rect 17512 10180 17540 10208
rect 19150 10180 19156 10192
rect 17512 10152 19156 10180
rect 11992 10084 18092 10112
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10013 5687 10047
rect 7926 10044 7932 10056
rect 5629 10007 5687 10013
rect 7668 10016 7932 10044
rect 5445 9979 5503 9985
rect 5445 9976 5457 9979
rect 5184 9948 5457 9976
rect 5445 9945 5457 9948
rect 5491 9945 5503 9979
rect 5445 9939 5503 9945
rect 5166 9908 5172 9920
rect 3252 9880 5172 9908
rect 5166 9868 5172 9880
rect 5224 9868 5230 9920
rect 5644 9908 5672 10007
rect 7668 9917 7696 10016
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 9456 10016 10241 10044
rect 9456 10004 9462 10016
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 10502 10004 10508 10056
rect 10560 10044 10566 10056
rect 10870 10044 10876 10056
rect 10560 10016 10876 10044
rect 10560 10004 10566 10016
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 12710 10044 12716 10056
rect 12671 10016 12716 10044
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 13909 10047 13967 10053
rect 13909 10044 13921 10047
rect 13320 10016 13921 10044
rect 13320 10004 13326 10016
rect 13909 10013 13921 10016
rect 13955 10044 13967 10047
rect 14090 10044 14096 10056
rect 13955 10016 14096 10044
rect 13955 10013 13967 10016
rect 13909 10007 13967 10013
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 14550 10004 14556 10056
rect 14608 10044 14614 10056
rect 15194 10044 15200 10056
rect 14608 10016 15200 10044
rect 14608 10004 14614 10016
rect 15194 10004 15200 10016
rect 15252 10044 15258 10056
rect 15838 10044 15844 10056
rect 15252 10016 15844 10044
rect 15252 10004 15258 10016
rect 15838 10004 15844 10016
rect 15896 10044 15902 10056
rect 16114 10044 16120 10056
rect 15896 10016 16120 10044
rect 15896 10004 15902 10016
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 9582 9936 9588 9988
rect 9640 9976 9646 9988
rect 9677 9979 9735 9985
rect 9677 9976 9689 9979
rect 9640 9948 9689 9976
rect 9640 9936 9646 9948
rect 9677 9945 9689 9948
rect 9723 9945 9735 9979
rect 9677 9939 9735 9945
rect 12544 9948 13492 9976
rect 7653 9911 7711 9917
rect 7653 9908 7665 9911
rect 5644 9880 7665 9908
rect 7653 9877 7665 9880
rect 7699 9877 7711 9911
rect 7653 9871 7711 9877
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 11882 9908 11888 9920
rect 7892 9880 11888 9908
rect 7892 9868 7898 9880
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12250 9868 12256 9920
rect 12308 9908 12314 9920
rect 12308 9880 12353 9908
rect 12308 9868 12314 9880
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12544 9908 12572 9948
rect 13354 9908 13360 9920
rect 12492 9880 12572 9908
rect 13315 9880 13360 9908
rect 12492 9868 12498 9880
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 13464 9908 13492 9948
rect 13998 9936 14004 9988
rect 14056 9976 14062 9988
rect 14642 9976 14648 9988
rect 14056 9948 14648 9976
rect 14056 9936 14062 9948
rect 14642 9936 14648 9948
rect 14700 9936 14706 9988
rect 17954 9976 17960 9988
rect 17052 9948 17960 9976
rect 17052 9908 17080 9948
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 13464 9880 17080 9908
rect 18064 9908 18092 10084
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 18288 10084 18429 10112
rect 18288 10072 18294 10084
rect 18417 10081 18429 10084
rect 18463 10081 18475 10115
rect 18417 10075 18475 10081
rect 18138 10004 18144 10056
rect 18196 10044 18202 10056
rect 18616 10053 18644 10152
rect 19150 10140 19156 10152
rect 19208 10140 19214 10192
rect 19705 10183 19763 10189
rect 19705 10149 19717 10183
rect 19751 10180 19763 10183
rect 19794 10180 19800 10192
rect 19751 10152 19800 10180
rect 19751 10149 19763 10152
rect 19705 10143 19763 10149
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 19058 10072 19064 10124
rect 19116 10112 19122 10124
rect 19334 10112 19340 10124
rect 19116 10084 19340 10112
rect 19116 10072 19122 10084
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19613 10115 19671 10121
rect 19613 10081 19625 10115
rect 19659 10112 19671 10115
rect 19978 10112 19984 10124
rect 19659 10084 19984 10112
rect 19659 10081 19671 10084
rect 19613 10075 19671 10081
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 18196 10016 18521 10044
rect 18196 10004 18202 10016
rect 18509 10013 18521 10016
rect 18555 10013 18567 10047
rect 18509 10007 18567 10013
rect 18601 10047 18659 10053
rect 18601 10013 18613 10047
rect 18647 10013 18659 10047
rect 19702 10044 19708 10056
rect 18601 10007 18659 10013
rect 18708 10016 19708 10044
rect 18524 9976 18552 10007
rect 18708 9976 18736 10016
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 19797 10047 19855 10053
rect 19797 10013 19809 10047
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 18524 9948 18736 9976
rect 19150 9936 19156 9988
rect 19208 9976 19214 9988
rect 19812 9976 19840 10007
rect 19208 9948 19840 9976
rect 19208 9936 19214 9948
rect 18782 9908 18788 9920
rect 18064 9880 18788 9908
rect 18782 9868 18788 9880
rect 18840 9868 18846 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 7009 9707 7067 9713
rect 3016 9676 4016 9704
rect 3016 9664 3022 9676
rect 1762 9636 1768 9648
rect 1723 9608 1768 9636
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 2498 9568 2504 9580
rect 2455 9540 2504 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 1486 9460 1492 9512
rect 1544 9500 1550 9512
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 1544 9472 2145 9500
rect 1544 9460 1550 9472
rect 2133 9469 2145 9472
rect 2179 9469 2191 9503
rect 2133 9463 2191 9469
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 3988 9500 4016 9676
rect 7009 9673 7021 9707
rect 7055 9704 7067 9707
rect 7098 9704 7104 9716
rect 7055 9676 7104 9704
rect 7055 9673 7067 9676
rect 7009 9667 7067 9673
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 7834 9704 7840 9716
rect 7208 9676 7840 9704
rect 4157 9639 4215 9645
rect 4157 9605 4169 9639
rect 4203 9605 4215 9639
rect 4157 9599 4215 9605
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 4706 9636 4712 9648
rect 4571 9608 4712 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 4172 9568 4200 9599
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 4798 9596 4804 9648
rect 4856 9636 4862 9648
rect 5442 9636 5448 9648
rect 4856 9608 5448 9636
rect 4856 9596 4862 9608
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 5626 9636 5632 9648
rect 5587 9608 5632 9636
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 4172 9540 5181 9568
rect 5169 9537 5181 9540
rect 5215 9568 5227 9571
rect 6270 9568 6276 9580
rect 5215 9540 6276 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5552 9512 5580 9540
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 3988 9472 5396 9500
rect 2777 9463 2835 9469
rect 1578 9392 1584 9444
rect 1636 9432 1642 9444
rect 2792 9432 2820 9463
rect 1636 9404 2820 9432
rect 1636 9392 1642 9404
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 3022 9435 3080 9441
rect 3022 9432 3034 9435
rect 2924 9404 3034 9432
rect 2924 9392 2930 9404
rect 3022 9401 3034 9404
rect 3068 9401 3080 9435
rect 4706 9432 4712 9444
rect 3022 9395 3080 9401
rect 3896 9404 4712 9432
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 3896 9364 3924 9404
rect 4706 9392 4712 9404
rect 4764 9392 4770 9444
rect 4798 9392 4804 9444
rect 4856 9432 4862 9444
rect 4985 9435 5043 9441
rect 4985 9432 4997 9435
rect 4856 9404 4997 9432
rect 4856 9392 4862 9404
rect 4985 9401 4997 9404
rect 5031 9401 5043 9435
rect 4985 9395 5043 9401
rect 2271 9336 3924 9364
rect 4893 9367 4951 9373
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 4893 9333 4905 9367
rect 4939 9364 4951 9367
rect 5166 9364 5172 9376
rect 4939 9336 5172 9364
rect 4939 9333 4951 9336
rect 4893 9327 4951 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5368 9364 5396 9472
rect 5534 9460 5540 9512
rect 5592 9460 5598 9512
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 6052 9472 6101 9500
rect 6052 9460 6058 9472
rect 6089 9469 6101 9472
rect 6135 9500 6147 9503
rect 7208 9500 7236 9676
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 9398 9704 9404 9716
rect 8352 9676 9404 9704
rect 8352 9664 8358 9676
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 12158 9704 12164 9716
rect 9508 9676 12164 9704
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9568 7711 9571
rect 7699 9540 8156 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 6135 9472 7236 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7984 9472 8033 9500
rect 7984 9460 7990 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 8128 9500 8156 9540
rect 8277 9503 8335 9509
rect 8277 9500 8289 9503
rect 8128 9472 8289 9500
rect 8021 9463 8079 9469
rect 8277 9469 8289 9472
rect 8323 9500 8335 9503
rect 9306 9500 9312 9512
rect 8323 9472 9312 9500
rect 8323 9469 8335 9472
rect 8277 9463 8335 9469
rect 5442 9392 5448 9444
rect 5500 9432 5506 9444
rect 7469 9435 7527 9441
rect 7469 9432 7481 9435
rect 5500 9404 7481 9432
rect 5500 9392 5506 9404
rect 7469 9401 7481 9404
rect 7515 9401 7527 9435
rect 7469 9395 7527 9401
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 5368 9336 6009 9364
rect 5997 9333 6009 9336
rect 6043 9364 6055 9367
rect 7098 9364 7104 9376
rect 6043 9336 7104 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7374 9364 7380 9376
rect 7335 9336 7380 9364
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 8036 9364 8064 9463
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 8202 9364 8208 9376
rect 8036 9336 8208 9364
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 9416 9373 9444 9664
rect 9508 9580 9536 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12360 9676 12664 9704
rect 10870 9596 10876 9648
rect 10928 9636 10934 9648
rect 12069 9639 12127 9645
rect 12069 9636 12081 9639
rect 10928 9608 12081 9636
rect 10928 9596 10934 9608
rect 12069 9605 12081 9608
rect 12115 9636 12127 9639
rect 12360 9636 12388 9676
rect 12115 9608 12388 9636
rect 12437 9639 12495 9645
rect 12115 9605 12127 9608
rect 12069 9599 12127 9605
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 12526 9636 12532 9648
rect 12483 9608 12532 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 12636 9636 12664 9676
rect 16390 9664 16396 9716
rect 16448 9704 16454 9716
rect 18506 9704 18512 9716
rect 16448 9676 18512 9704
rect 16448 9664 16454 9676
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 20530 9664 20536 9716
rect 20588 9704 20594 9716
rect 21082 9704 21088 9716
rect 20588 9676 21088 9704
rect 20588 9664 20594 9676
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 16574 9636 16580 9648
rect 12636 9608 13584 9636
rect 16535 9608 16580 9636
rect 9490 9528 9496 9580
rect 9548 9528 9554 9580
rect 10318 9568 10324 9580
rect 10279 9540 10324 9568
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10502 9568 10508 9580
rect 10463 9540 10508 9568
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 13556 9577 13584 9608
rect 16574 9596 16580 9608
rect 16632 9636 16638 9648
rect 18877 9639 18935 9645
rect 16632 9608 17448 9636
rect 16632 9596 16638 9608
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12400 9540 13001 9568
rect 12400 9528 12406 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9537 13599 9571
rect 13541 9531 13599 9537
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 14700 9540 15332 9568
rect 14700 9528 14706 9540
rect 10226 9500 10232 9512
rect 10187 9472 10232 9500
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 11882 9432 11888 9444
rect 9548 9404 11888 9432
rect 9548 9392 9554 9404
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 9401 9367 9459 9373
rect 9401 9333 9413 9367
rect 9447 9333 9459 9367
rect 9858 9364 9864 9376
rect 9819 9336 9864 9364
rect 9401 9327 9459 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 12268 9364 12296 9463
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12768 9472 12817 9500
rect 12768 9460 12774 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 13354 9500 13360 9512
rect 12943 9472 13360 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 15194 9500 15200 9512
rect 15155 9472 15200 9500
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 15304 9500 15332 9540
rect 16206 9528 16212 9580
rect 16264 9568 16270 9580
rect 17034 9568 17040 9580
rect 16264 9540 17040 9568
rect 16264 9528 16270 9540
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 17420 9577 17448 9608
rect 18877 9605 18889 9639
rect 18923 9636 18935 9639
rect 20622 9636 20628 9648
rect 18923 9608 20628 9636
rect 18923 9605 18935 9608
rect 18877 9599 18935 9605
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 17405 9571 17463 9577
rect 17405 9537 17417 9571
rect 17451 9537 17463 9571
rect 17405 9531 17463 9537
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 20533 9571 20591 9577
rect 20533 9537 20545 9571
rect 20579 9537 20591 9571
rect 20533 9531 20591 9537
rect 16390 9500 16396 9512
rect 15304 9472 16396 9500
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 16850 9460 16856 9512
rect 16908 9500 16914 9512
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 16908 9472 18153 9500
rect 16908 9460 16914 9472
rect 18141 9469 18153 9472
rect 18187 9469 18199 9503
rect 18141 9463 18199 9469
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 19337 9503 19395 9509
rect 19337 9500 19349 9503
rect 19300 9472 19349 9500
rect 19300 9460 19306 9472
rect 19337 9469 19349 9472
rect 19383 9469 19395 9503
rect 19536 9500 19564 9531
rect 19610 9500 19616 9512
rect 19536 9472 19616 9500
rect 19337 9463 19395 9469
rect 19610 9460 19616 9472
rect 19668 9460 19674 9512
rect 20548 9500 20576 9531
rect 20548 9472 20668 9500
rect 20640 9444 20668 9472
rect 13814 9441 13820 9444
rect 13808 9432 13820 9441
rect 13775 9404 13820 9432
rect 13808 9395 13820 9404
rect 13814 9392 13820 9395
rect 13872 9392 13878 9444
rect 15010 9432 15016 9444
rect 14923 9404 15016 9432
rect 13906 9364 13912 9376
rect 12268 9336 13912 9364
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 14936 9373 14964 9404
rect 15010 9392 15016 9404
rect 15068 9432 15074 9444
rect 15464 9435 15522 9441
rect 15464 9432 15476 9435
rect 15068 9404 15476 9432
rect 15068 9392 15074 9404
rect 15464 9401 15476 9404
rect 15510 9432 15522 9435
rect 15838 9432 15844 9444
rect 15510 9404 15844 9432
rect 15510 9401 15522 9404
rect 15464 9395 15522 9401
rect 15838 9392 15844 9404
rect 15896 9392 15902 9444
rect 16022 9392 16028 9444
rect 16080 9432 16086 9444
rect 17313 9435 17371 9441
rect 17313 9432 17325 9435
rect 16080 9404 17325 9432
rect 16080 9392 16086 9404
rect 17313 9401 17325 9404
rect 17359 9401 17371 9435
rect 17313 9395 17371 9401
rect 18417 9435 18475 9441
rect 18417 9401 18429 9435
rect 18463 9432 18475 9435
rect 20070 9432 20076 9444
rect 18463 9404 20076 9432
rect 18463 9401 18475 9404
rect 18417 9395 18475 9401
rect 20070 9392 20076 9404
rect 20128 9392 20134 9444
rect 20257 9435 20315 9441
rect 20257 9401 20269 9435
rect 20303 9432 20315 9435
rect 20530 9432 20536 9444
rect 20303 9404 20536 9432
rect 20303 9401 20315 9404
rect 20257 9395 20315 9401
rect 20530 9392 20536 9404
rect 20588 9392 20594 9444
rect 20622 9392 20628 9444
rect 20680 9392 20686 9444
rect 14921 9367 14979 9373
rect 14921 9333 14933 9367
rect 14967 9333 14979 9367
rect 14921 9327 14979 9333
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 17218 9364 17224 9376
rect 16908 9336 16953 9364
rect 17179 9336 17224 9364
rect 16908 9324 16914 9336
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 19245 9367 19303 9373
rect 19245 9333 19257 9367
rect 19291 9364 19303 9367
rect 19518 9364 19524 9376
rect 19291 9336 19524 9364
rect 19291 9333 19303 9336
rect 19245 9327 19303 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 19886 9364 19892 9376
rect 19847 9336 19892 9364
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 20162 9324 20168 9376
rect 20220 9364 20226 9376
rect 20349 9367 20407 9373
rect 20349 9364 20361 9367
rect 20220 9336 20361 9364
rect 20220 9324 20226 9336
rect 20349 9333 20361 9336
rect 20395 9333 20407 9367
rect 20349 9327 20407 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1118 9120 1124 9172
rect 1176 9160 1182 9172
rect 3602 9160 3608 9172
rect 1176 9132 3608 9160
rect 1176 9120 1182 9132
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 4246 9160 4252 9172
rect 4207 9132 4252 9160
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 4617 9163 4675 9169
rect 4617 9129 4629 9163
rect 4663 9160 4675 9163
rect 4982 9160 4988 9172
rect 4663 9132 4988 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 5718 9120 5724 9172
rect 5776 9160 5782 9172
rect 6086 9160 6092 9172
rect 5776 9132 6092 9160
rect 5776 9120 5782 9132
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 8478 9160 8484 9172
rect 8439 9132 8484 9160
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 9858 9120 9864 9172
rect 9916 9160 9922 9172
rect 9916 9132 12480 9160
rect 9916 9120 9922 9132
rect 1394 9052 1400 9104
rect 1452 9092 1458 9104
rect 1765 9095 1823 9101
rect 1765 9092 1777 9095
rect 1452 9064 1777 9092
rect 1452 9052 1458 9064
rect 1765 9061 1777 9064
rect 1811 9061 1823 9095
rect 1765 9055 1823 9061
rect 3142 9052 3148 9104
rect 3200 9092 3206 9104
rect 3513 9095 3571 9101
rect 3513 9092 3525 9095
rect 3200 9064 3525 9092
rect 3200 9052 3206 9064
rect 3513 9061 3525 9064
rect 3559 9061 3571 9095
rect 5258 9092 5264 9104
rect 3513 9055 3571 9061
rect 4724 9064 5264 9092
rect 1489 9027 1547 9033
rect 1489 8993 1501 9027
rect 1535 8993 1547 9027
rect 1489 8987 1547 8993
rect 1504 8820 1532 8987
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 2593 9027 2651 9033
rect 2593 9024 2605 9027
rect 1912 8996 2605 9024
rect 1912 8984 1918 8996
rect 2593 8993 2605 8996
rect 2639 8993 2651 9027
rect 2593 8987 2651 8993
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 8993 3295 9027
rect 3237 8987 3295 8993
rect 2682 8956 2688 8968
rect 2643 8928 2688 8956
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 2225 8891 2283 8897
rect 2225 8857 2237 8891
rect 2271 8888 2283 8891
rect 3252 8888 3280 8987
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 4724 8965 4752 9064
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 5442 9052 5448 9104
rect 5500 9092 5506 9104
rect 7374 9092 7380 9104
rect 5500 9064 7380 9092
rect 5500 9052 5506 9064
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 7837 9095 7895 9101
rect 7837 9061 7849 9095
rect 7883 9092 7895 9095
rect 8570 9092 8576 9104
rect 7883 9064 8576 9092
rect 7883 9061 7895 9064
rect 7837 9055 7895 9061
rect 8570 9052 8576 9064
rect 8628 9092 8634 9104
rect 9490 9092 9496 9104
rect 8628 9064 9496 9092
rect 8628 9052 8634 9064
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 10312 9095 10370 9101
rect 10312 9061 10324 9095
rect 10358 9092 10370 9095
rect 11790 9092 11796 9104
rect 10358 9064 11796 9092
rect 10358 9061 10370 9064
rect 10312 9055 10370 9061
rect 11790 9052 11796 9064
rect 11848 9092 11854 9104
rect 12250 9092 12256 9104
rect 11848 9064 12256 9092
rect 11848 9052 11854 9064
rect 12250 9052 12256 9064
rect 12308 9052 12314 9104
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 5132 8996 5641 9024
rect 5132 8984 5138 8996
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 7929 9027 7987 9033
rect 6788 8996 7696 9024
rect 6788 8984 6794 8996
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 3660 8928 4721 8956
rect 3660 8916 3666 8928
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8956 4951 8959
rect 5534 8956 5540 8968
rect 4939 8928 5540 8956
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5718 8956 5724 8968
rect 5679 8928 5724 8956
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 6914 8956 6920 8968
rect 5951 8928 6920 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 2271 8860 3280 8888
rect 2271 8857 2283 8860
rect 2225 8851 2283 8857
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 7668 8888 7696 8996
rect 7929 8993 7941 9027
rect 7975 9024 7987 9027
rect 8294 9024 8300 9036
rect 7975 8996 8300 9024
rect 7975 8993 7987 8996
rect 7929 8987 7987 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 12066 9024 12072 9036
rect 10928 8996 12072 9024
rect 10928 8984 10934 8996
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 12342 9033 12348 9036
rect 12336 9024 12348 9033
rect 12303 8996 12348 9024
rect 12336 8987 12348 8996
rect 12342 8984 12348 8987
rect 12400 8984 12406 9036
rect 12452 9024 12480 9132
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 13722 9160 13728 9172
rect 12584 9132 13728 9160
rect 12584 9120 12590 9132
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9160 14243 9163
rect 16022 9160 16028 9172
rect 14231 9132 16028 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 16758 9160 16764 9172
rect 16719 9132 16764 9160
rect 16758 9120 16764 9132
rect 16816 9120 16822 9172
rect 16850 9120 16856 9172
rect 16908 9160 16914 9172
rect 17218 9160 17224 9172
rect 16908 9132 17224 9160
rect 16908 9120 16914 9132
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 20070 9120 20076 9172
rect 20128 9160 20134 9172
rect 20346 9160 20352 9172
rect 20128 9132 20352 9160
rect 20128 9120 20134 9132
rect 20346 9120 20352 9132
rect 20404 9120 20410 9172
rect 12710 9052 12716 9104
rect 12768 9092 12774 9104
rect 19610 9092 19616 9104
rect 12768 9064 19616 9092
rect 12768 9052 12774 9064
rect 19610 9052 19616 9064
rect 19668 9092 19674 9104
rect 19668 9064 19932 9092
rect 19668 9052 19674 9064
rect 14458 9024 14464 9036
rect 12452 8996 14464 9024
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 14553 9027 14611 9033
rect 14553 8993 14565 9027
rect 14599 9024 14611 9027
rect 15286 9024 15292 9036
rect 14599 8996 15292 9024
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15396 8996 15669 9024
rect 8018 8956 8024 8968
rect 7979 8928 8024 8956
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 8260 8928 10057 8956
rect 8260 8916 8266 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 14090 8916 14096 8968
rect 14148 8956 14154 8968
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 14148 8928 14657 8956
rect 14148 8916 14154 8928
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 14645 8919 14703 8925
rect 14829 8959 14887 8965
rect 14829 8925 14841 8959
rect 14875 8956 14887 8959
rect 15010 8956 15016 8968
rect 14875 8928 15016 8956
rect 14875 8925 14887 8928
rect 14829 8919 14887 8925
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 9950 8888 9956 8900
rect 4120 8860 7604 8888
rect 7668 8860 9956 8888
rect 4120 8848 4126 8860
rect 5261 8823 5319 8829
rect 5261 8820 5273 8823
rect 1504 8792 5273 8820
rect 5261 8789 5273 8792
rect 5307 8789 5319 8823
rect 5261 8783 5319 8789
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 7469 8823 7527 8829
rect 7469 8820 7481 8823
rect 5592 8792 7481 8820
rect 5592 8780 5598 8792
rect 7469 8789 7481 8792
rect 7515 8789 7527 8823
rect 7576 8820 7604 8860
rect 9950 8848 9956 8860
rect 10008 8848 10014 8900
rect 13446 8888 13452 8900
rect 10980 8860 11744 8888
rect 13407 8860 13452 8888
rect 10980 8820 11008 8860
rect 7576 8792 11008 8820
rect 11425 8823 11483 8829
rect 7469 8783 7527 8789
rect 11425 8789 11437 8823
rect 11471 8820 11483 8823
rect 11606 8820 11612 8832
rect 11471 8792 11612 8820
rect 11471 8789 11483 8792
rect 11425 8783 11483 8789
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 11716 8820 11744 8860
rect 13446 8848 13452 8860
rect 13504 8888 13510 8900
rect 13814 8888 13820 8900
rect 13504 8860 13820 8888
rect 13504 8848 13510 8860
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 14274 8848 14280 8900
rect 14332 8888 14338 8900
rect 15396 8888 15424 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 15746 8984 15752 9036
rect 15804 9024 15810 9036
rect 16117 9027 16175 9033
rect 16117 9024 16129 9027
rect 15804 8996 16129 9024
rect 15804 8984 15810 8996
rect 16117 8993 16129 8996
rect 16163 8993 16175 9027
rect 16117 8987 16175 8993
rect 16669 9027 16727 9033
rect 16669 8993 16681 9027
rect 16715 9024 16727 9027
rect 17313 9027 17371 9033
rect 17313 9024 17325 9027
rect 16715 8996 17325 9024
rect 16715 8993 16727 8996
rect 16669 8987 16727 8993
rect 17313 8993 17325 8996
rect 17359 8993 17371 9027
rect 17313 8987 17371 8993
rect 18776 9027 18834 9033
rect 18776 8993 18788 9027
rect 18822 9024 18834 9027
rect 19334 9024 19340 9036
rect 18822 8996 19340 9024
rect 18822 8993 18834 8996
rect 18776 8987 18834 8993
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 15933 8959 15991 8965
rect 15933 8956 15945 8959
rect 15764 8928 15945 8956
rect 14332 8860 15424 8888
rect 14332 8848 14338 8860
rect 15654 8848 15660 8900
rect 15712 8888 15718 8900
rect 15764 8888 15792 8928
rect 15933 8925 15945 8928
rect 15979 8956 15991 8959
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 15979 8928 16865 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 18509 8959 18567 8965
rect 18509 8956 18521 8959
rect 17920 8928 18521 8956
rect 17920 8916 17926 8928
rect 18509 8925 18521 8928
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 15712 8860 15792 8888
rect 16117 8891 16175 8897
rect 15712 8848 15718 8860
rect 16117 8857 16129 8891
rect 16163 8888 16175 8891
rect 17494 8888 17500 8900
rect 16163 8860 17500 8888
rect 16163 8857 16175 8860
rect 16117 8851 16175 8857
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 19904 8897 19932 9064
rect 19889 8891 19947 8897
rect 19889 8857 19901 8891
rect 19935 8857 19947 8891
rect 19889 8851 19947 8857
rect 14182 8820 14188 8832
rect 11716 8792 14188 8820
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 15289 8823 15347 8829
rect 15289 8789 15301 8823
rect 15335 8820 15347 8823
rect 15746 8820 15752 8832
rect 15335 8792 15752 8820
rect 15335 8789 15347 8792
rect 15289 8783 15347 8789
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 16298 8820 16304 8832
rect 16259 8792 16304 8820
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 16390 8780 16396 8832
rect 16448 8820 16454 8832
rect 19794 8820 19800 8832
rect 16448 8792 19800 8820
rect 16448 8780 16454 8792
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3053 8619 3111 8625
rect 3053 8616 3065 8619
rect 2924 8588 3065 8616
rect 2924 8576 2930 8588
rect 3053 8585 3065 8588
rect 3099 8585 3111 8619
rect 3053 8579 3111 8585
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4617 8619 4675 8625
rect 4617 8616 4629 8619
rect 4212 8588 4629 8616
rect 4212 8576 4218 8588
rect 4617 8585 4629 8588
rect 4663 8585 4675 8619
rect 5718 8616 5724 8628
rect 5679 8588 5724 8616
rect 4617 8579 4675 8585
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 12434 8616 12440 8628
rect 6052 8588 12440 8616
rect 6052 8576 6058 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 14090 8616 14096 8628
rect 12676 8588 13400 8616
rect 14051 8588 14096 8616
rect 12676 8576 12682 8588
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 4338 8548 4344 8560
rect 3651 8520 4344 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 8018 8548 8024 8560
rect 5736 8520 8024 8548
rect 2682 8440 2688 8492
rect 2740 8480 2746 8492
rect 3970 8480 3976 8492
rect 2740 8452 3976 8480
rect 2740 8440 2746 8452
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4154 8480 4160 8492
rect 4115 8452 4160 8480
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5626 8480 5632 8492
rect 5307 8452 5632 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 1578 8372 1584 8424
rect 1636 8412 1642 8424
rect 1673 8415 1731 8421
rect 1673 8412 1685 8415
rect 1636 8384 1685 8412
rect 1636 8372 1642 8384
rect 1673 8381 1685 8384
rect 1719 8381 1731 8415
rect 1673 8375 1731 8381
rect 4430 8372 4436 8424
rect 4488 8412 4494 8424
rect 5077 8415 5135 8421
rect 5077 8412 5089 8415
rect 4488 8384 5089 8412
rect 4488 8372 4494 8384
rect 5077 8381 5089 8384
rect 5123 8412 5135 8415
rect 5442 8412 5448 8424
rect 5123 8384 5448 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 1940 8347 1998 8353
rect 1940 8313 1952 8347
rect 1986 8344 1998 8347
rect 2314 8344 2320 8356
rect 1986 8316 2320 8344
rect 1986 8313 1998 8316
rect 1940 8307 1998 8313
rect 2314 8304 2320 8316
rect 2372 8304 2378 8356
rect 2498 8304 2504 8356
rect 2556 8344 2562 8356
rect 3694 8344 3700 8356
rect 2556 8316 3700 8344
rect 2556 8304 2562 8316
rect 3694 8304 3700 8316
rect 3752 8344 3758 8356
rect 3973 8347 4031 8353
rect 3973 8344 3985 8347
rect 3752 8316 3985 8344
rect 3752 8304 3758 8316
rect 3973 8313 3985 8316
rect 4019 8313 4031 8347
rect 3973 8307 4031 8313
rect 4154 8304 4160 8356
rect 4212 8344 4218 8356
rect 4338 8344 4344 8356
rect 4212 8316 4344 8344
rect 4212 8304 4218 8316
rect 4338 8304 4344 8316
rect 4396 8344 4402 8356
rect 5736 8344 5764 8520
rect 8018 8508 8024 8520
rect 8076 8548 8082 8560
rect 8570 8548 8576 8560
rect 8076 8520 8576 8548
rect 8076 8508 8082 8520
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 11054 8548 11060 8560
rect 10704 8520 11060 8548
rect 6273 8483 6331 8489
rect 6273 8480 6285 8483
rect 4396 8316 5764 8344
rect 6012 8452 6285 8480
rect 4396 8304 4402 8316
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 3786 8276 3792 8288
rect 2832 8248 3792 8276
rect 2832 8236 2838 8248
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4065 8279 4123 8285
rect 4065 8245 4077 8279
rect 4111 8276 4123 8279
rect 4614 8276 4620 8288
rect 4111 8248 4620 8276
rect 4111 8245 4123 8248
rect 4065 8239 4123 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 4985 8279 5043 8285
rect 4985 8276 4997 8279
rect 4764 8248 4997 8276
rect 4764 8236 4770 8248
rect 4985 8245 4997 8248
rect 5031 8245 5043 8279
rect 4985 8239 5043 8245
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 6012 8276 6040 8452
rect 6273 8449 6285 8452
rect 6319 8449 6331 8483
rect 6273 8443 6331 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 7699 8452 8708 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 6181 8415 6239 8421
rect 6181 8381 6193 8415
rect 6227 8412 6239 8415
rect 8202 8412 8208 8424
rect 6227 8384 8208 8412
rect 6227 8381 6239 8384
rect 6181 8375 6239 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8381 8631 8415
rect 8680 8412 8708 8452
rect 9950 8440 9956 8492
rect 10008 8480 10014 8492
rect 10704 8489 10732 8520
rect 11054 8508 11060 8520
rect 11112 8508 11118 8560
rect 13372 8548 13400 8588
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 14182 8576 14188 8628
rect 14240 8616 14246 8628
rect 15470 8616 15476 8628
rect 14240 8588 15476 8616
rect 14240 8576 14246 8588
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 16666 8616 16672 8628
rect 15620 8588 16672 8616
rect 15620 8576 15626 8588
rect 16666 8576 16672 8588
rect 16724 8616 16730 8628
rect 17402 8616 17408 8628
rect 16724 8588 17408 8616
rect 16724 8576 16730 8588
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 17552 8588 19012 8616
rect 17552 8576 17558 8588
rect 16577 8551 16635 8557
rect 13372 8520 15976 8548
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 10008 8452 10701 8480
rect 10008 8440 10014 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 11606 8480 11612 8492
rect 10827 8452 11612 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 8829 8415 8887 8421
rect 8829 8412 8841 8415
rect 8680 8384 8841 8412
rect 8573 8375 8631 8381
rect 8829 8381 8841 8384
rect 8875 8412 8887 8415
rect 10796 8412 10824 8443
rect 11606 8440 11612 8452
rect 11664 8480 11670 8492
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11664 8452 11805 8480
rect 11664 8440 11670 8452
rect 11793 8449 11805 8452
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 13446 8440 13452 8492
rect 13504 8480 13510 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 13504 8452 14749 8480
rect 13504 8440 13510 8452
rect 14737 8449 14749 8452
rect 14783 8480 14795 8483
rect 15654 8480 15660 8492
rect 14783 8452 15660 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 15654 8440 15660 8452
rect 15712 8480 15718 8492
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 15712 8452 15853 8480
rect 15712 8440 15718 8452
rect 15841 8449 15853 8452
rect 15887 8449 15899 8483
rect 15948 8480 15976 8520
rect 16577 8517 16589 8551
rect 16623 8548 16635 8551
rect 18046 8548 18052 8560
rect 16623 8520 18052 8548
rect 16623 8517 16635 8520
rect 16577 8511 16635 8517
rect 18046 8508 18052 8520
rect 18104 8508 18110 8560
rect 18984 8548 19012 8588
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 19392 8588 19441 8616
rect 19392 8576 19398 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 20070 8548 20076 8560
rect 18984 8520 20076 8548
rect 20070 8508 20076 8520
rect 20128 8508 20134 8560
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 15948 8452 17049 8480
rect 15841 8443 15899 8449
rect 17037 8449 17049 8452
rect 17083 8449 17095 8483
rect 17218 8480 17224 8492
rect 17179 8452 17224 8480
rect 17037 8443 17095 8449
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 20441 8483 20499 8489
rect 20441 8449 20453 8483
rect 20487 8480 20499 8483
rect 20622 8480 20628 8492
rect 20487 8452 20628 8480
rect 20487 8449 20499 8452
rect 20441 8443 20499 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 11698 8412 11704 8424
rect 8875 8384 10824 8412
rect 11659 8384 11704 8412
rect 8875 8381 8887 8384
rect 8829 8375 8887 8381
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8344 6147 8347
rect 7190 8344 7196 8356
rect 6135 8316 7196 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 8110 8344 8116 8356
rect 7616 8316 8116 8344
rect 7616 8304 7622 8316
rect 8110 8304 8116 8316
rect 8168 8344 8174 8356
rect 8588 8344 8616 8375
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 12066 8372 12072 8424
rect 12124 8412 12130 8424
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 12124 8384 12449 8412
rect 12124 8372 12130 8384
rect 12437 8381 12449 8384
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 16942 8412 16948 8424
rect 14599 8384 14688 8412
rect 16903 8384 16948 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 8168 8316 8616 8344
rect 10597 8347 10655 8353
rect 8168 8304 8174 8316
rect 10597 8313 10609 8347
rect 10643 8344 10655 8347
rect 10962 8344 10968 8356
rect 10643 8316 10968 8344
rect 10643 8313 10655 8316
rect 10597 8307 10655 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 11609 8347 11667 8353
rect 11609 8344 11621 8347
rect 11204 8316 11621 8344
rect 11204 8304 11210 8316
rect 11609 8313 11621 8316
rect 11655 8344 11667 8347
rect 12250 8344 12256 8356
rect 11655 8316 12256 8344
rect 11655 8313 11667 8316
rect 11609 8307 11667 8313
rect 12250 8304 12256 8316
rect 12308 8304 12314 8356
rect 12710 8353 12716 8356
rect 12704 8344 12716 8353
rect 12671 8316 12716 8344
rect 12704 8307 12716 8316
rect 12710 8304 12716 8307
rect 12768 8304 12774 8356
rect 14461 8347 14519 8353
rect 14461 8313 14473 8347
rect 14507 8313 14519 8347
rect 14461 8307 14519 8313
rect 7006 8276 7012 8288
rect 5776 8248 6040 8276
rect 6967 8248 7012 8276
rect 5776 8236 5782 8248
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 7098 8236 7104 8288
rect 7156 8276 7162 8288
rect 7377 8279 7435 8285
rect 7377 8276 7389 8279
rect 7156 8248 7389 8276
rect 7156 8236 7162 8248
rect 7377 8245 7389 8248
rect 7423 8245 7435 8279
rect 7377 8239 7435 8245
rect 7469 8279 7527 8285
rect 7469 8245 7481 8279
rect 7515 8276 7527 8279
rect 8846 8276 8852 8288
rect 7515 8248 8852 8276
rect 7515 8245 7527 8248
rect 7469 8239 7527 8245
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 9950 8276 9956 8288
rect 9911 8248 9956 8276
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 10226 8276 10232 8288
rect 10187 8248 10232 8276
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 10318 8236 10324 8288
rect 10376 8276 10382 8288
rect 11241 8279 11299 8285
rect 11241 8276 11253 8279
rect 10376 8248 11253 8276
rect 10376 8236 10382 8248
rect 11241 8245 11253 8248
rect 11287 8245 11299 8279
rect 11241 8239 11299 8245
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 13817 8279 13875 8285
rect 13817 8276 13829 8279
rect 13320 8248 13829 8276
rect 13320 8236 13326 8248
rect 13817 8245 13829 8248
rect 13863 8245 13875 8279
rect 13817 8239 13875 8245
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 14476 8276 14504 8307
rect 13964 8248 14504 8276
rect 14660 8276 14688 8384
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 17126 8372 17132 8424
rect 17184 8412 17190 8424
rect 17862 8412 17868 8424
rect 17184 8384 17868 8412
rect 17184 8372 17190 8384
rect 17862 8372 17868 8384
rect 17920 8412 17926 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17920 8384 18061 8412
rect 17920 8372 17926 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20036 8384 20300 8412
rect 20036 8372 20042 8384
rect 18316 8347 18374 8353
rect 18316 8313 18328 8347
rect 18362 8344 18374 8347
rect 18598 8344 18604 8356
rect 18362 8316 18604 8344
rect 18362 8313 18374 8316
rect 18316 8307 18374 8313
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 19150 8304 19156 8356
rect 19208 8344 19214 8356
rect 20165 8347 20223 8353
rect 20165 8344 20177 8347
rect 19208 8316 20177 8344
rect 19208 8304 19214 8316
rect 20165 8313 20177 8316
rect 20211 8313 20223 8347
rect 20165 8307 20223 8313
rect 15010 8276 15016 8288
rect 14660 8248 15016 8276
rect 13964 8236 13970 8248
rect 15010 8236 15016 8248
rect 15068 8236 15074 8288
rect 15286 8276 15292 8288
rect 15247 8248 15292 8276
rect 15286 8236 15292 8248
rect 15344 8236 15350 8288
rect 15562 8236 15568 8288
rect 15620 8276 15626 8288
rect 15657 8279 15715 8285
rect 15657 8276 15669 8279
rect 15620 8248 15669 8276
rect 15620 8236 15626 8248
rect 15657 8245 15669 8248
rect 15703 8245 15715 8279
rect 15657 8239 15715 8245
rect 15749 8279 15807 8285
rect 15749 8245 15761 8279
rect 15795 8276 15807 8279
rect 16390 8276 16396 8288
rect 15795 8248 16396 8276
rect 15795 8245 15807 8248
rect 15749 8239 15807 8245
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 19610 8236 19616 8288
rect 19668 8276 19674 8288
rect 20272 8285 20300 8384
rect 20346 8304 20352 8356
rect 20404 8344 20410 8356
rect 20809 8347 20867 8353
rect 20809 8344 20821 8347
rect 20404 8316 20821 8344
rect 20404 8304 20410 8316
rect 20809 8313 20821 8316
rect 20855 8313 20867 8347
rect 20809 8307 20867 8313
rect 19797 8279 19855 8285
rect 19797 8276 19809 8279
rect 19668 8248 19809 8276
rect 19668 8236 19674 8248
rect 19797 8245 19809 8248
rect 19843 8245 19855 8279
rect 19797 8239 19855 8245
rect 20257 8279 20315 8285
rect 20257 8245 20269 8279
rect 20303 8276 20315 8279
rect 20714 8276 20720 8288
rect 20303 8248 20720 8276
rect 20303 8245 20315 8248
rect 20257 8239 20315 8245
rect 20714 8236 20720 8248
rect 20772 8236 20778 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 1854 8072 1860 8084
rect 1811 8044 1860 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 1854 8032 1860 8044
rect 1912 8032 1918 8084
rect 2225 8075 2283 8081
rect 2225 8041 2237 8075
rect 2271 8072 2283 8075
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2271 8044 2789 8072
rect 2271 8041 2283 8044
rect 2225 8035 2283 8041
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 2777 8035 2835 8041
rect 3878 8032 3884 8084
rect 3936 8072 3942 8084
rect 4430 8072 4436 8084
rect 3936 8044 4436 8072
rect 3936 8032 3942 8044
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 5491 8044 6132 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 3602 8004 3608 8016
rect 3160 7976 3608 8004
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2774 7936 2780 7948
rect 2179 7908 2780 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 2866 7896 2872 7948
rect 2924 7936 2930 7948
rect 3160 7945 3188 7976
rect 3602 7964 3608 7976
rect 3660 7964 3666 8016
rect 4985 8007 5043 8013
rect 4985 7973 4997 8007
rect 5031 8004 5043 8007
rect 5994 8004 6000 8016
rect 5031 7976 6000 8004
rect 5031 7973 5043 7976
rect 4985 7967 5043 7973
rect 5994 7964 6000 7976
rect 6052 7964 6058 8016
rect 6104 8004 6132 8044
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7064 8044 7757 8072
rect 7064 8032 7070 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 8294 8072 8300 8084
rect 8255 8044 8300 8072
rect 7745 8035 7803 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9122 8072 9128 8084
rect 8803 8044 9128 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9122 8032 9128 8044
rect 9180 8072 9186 8084
rect 9582 8072 9588 8084
rect 9180 8044 9588 8072
rect 9180 8032 9186 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 10226 8072 10232 8084
rect 10183 8044 10232 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 15010 8072 15016 8084
rect 10735 8044 15016 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 16298 8072 16304 8084
rect 15703 8044 16304 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 18046 8032 18052 8084
rect 18104 8072 18110 8084
rect 19153 8075 19211 8081
rect 19153 8072 19165 8075
rect 18104 8044 19165 8072
rect 18104 8032 18110 8044
rect 19153 8041 19165 8044
rect 19199 8041 19211 8075
rect 19153 8035 19211 8041
rect 20165 8075 20223 8081
rect 20165 8041 20177 8075
rect 20211 8072 20223 8075
rect 20346 8072 20352 8084
rect 20211 8044 20352 8072
rect 20211 8041 20223 8044
rect 20165 8035 20223 8041
rect 20346 8032 20352 8044
rect 20404 8032 20410 8084
rect 9950 8004 9956 8016
rect 6104 7976 9956 8004
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 2924 7908 3157 7936
rect 2924 7896 2930 7908
rect 3145 7905 3157 7908
rect 3191 7905 3203 7939
rect 3145 7899 3203 7905
rect 3237 7939 3295 7945
rect 3237 7905 3249 7939
rect 3283 7936 3295 7939
rect 4154 7936 4160 7948
rect 3283 7908 4160 7936
rect 3283 7905 3295 7908
rect 3237 7899 3295 7905
rect 4154 7896 4160 7908
rect 4212 7936 4218 7948
rect 4798 7936 4804 7948
rect 4212 7908 4804 7936
rect 4212 7896 4218 7908
rect 4798 7896 4804 7908
rect 4856 7896 4862 7948
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 5885 7939 5943 7945
rect 5885 7936 5897 7939
rect 5776 7908 5897 7936
rect 5776 7896 5782 7908
rect 5885 7905 5897 7908
rect 5931 7905 5943 7939
rect 5885 7899 5943 7905
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 6328 7908 7665 7936
rect 6328 7896 6334 7908
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 7653 7899 7711 7905
rect 2314 7868 2320 7880
rect 2275 7840 2320 7868
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 3384 7840 3433 7868
rect 3384 7828 3390 7840
rect 3421 7837 3433 7840
rect 3467 7868 3479 7871
rect 4338 7868 4344 7880
rect 3467 7840 4344 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 5077 7871 5135 7877
rect 5077 7868 5089 7871
rect 4764 7840 5089 7868
rect 4764 7828 4770 7840
rect 5077 7837 5089 7840
rect 5123 7837 5135 7871
rect 5258 7868 5264 7880
rect 5171 7840 5264 7868
rect 5077 7831 5135 7837
rect 5258 7828 5264 7840
rect 5316 7868 5322 7880
rect 5445 7871 5503 7877
rect 5445 7868 5457 7871
rect 5316 7840 5457 7868
rect 5316 7828 5322 7840
rect 5445 7837 5457 7840
rect 5491 7837 5503 7871
rect 5626 7868 5632 7880
rect 5587 7840 5632 7868
rect 5445 7831 5503 7837
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8036 7868 8064 7976
rect 9950 7964 9956 7976
rect 10008 7964 10014 8016
rect 10045 8007 10103 8013
rect 10045 7973 10057 8007
rect 10091 8004 10103 8007
rect 10318 8004 10324 8016
rect 10091 7976 10324 8004
rect 10091 7973 10103 7976
rect 10045 7967 10103 7973
rect 10318 7964 10324 7976
rect 10376 7964 10382 8016
rect 11057 8007 11115 8013
rect 11057 8004 11069 8007
rect 10980 7976 11069 8004
rect 10980 7948 11008 7976
rect 11057 7973 11069 7976
rect 11103 7973 11115 8007
rect 11057 7967 11115 7973
rect 12526 7964 12532 8016
rect 12584 8004 12590 8016
rect 15378 8004 15384 8016
rect 12584 7976 15384 8004
rect 12584 7964 12590 7976
rect 15378 7964 15384 7976
rect 15436 7964 15442 8016
rect 15746 8004 15752 8016
rect 15707 7976 15752 8004
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 17218 7964 17224 8016
rect 17276 8013 17282 8016
rect 17276 8007 17340 8013
rect 17276 7973 17294 8007
rect 17328 7973 17340 8007
rect 20254 8004 20260 8016
rect 20215 7976 20260 8004
rect 17276 7967 17340 7973
rect 17276 7964 17282 7967
rect 20254 7964 20260 7976
rect 20312 7964 20318 8016
rect 8665 7939 8723 7945
rect 8665 7905 8677 7939
rect 8711 7936 8723 7939
rect 8711 7908 10916 7936
rect 8711 7905 8723 7908
rect 8665 7899 8723 7905
rect 7975 7840 8064 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 8904 7840 8949 7868
rect 8904 7828 8910 7840
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 10008 7840 10241 7868
rect 10008 7828 10014 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10888 7868 10916 7908
rect 10962 7896 10968 7948
rect 11020 7896 11026 7948
rect 11974 7936 11980 7948
rect 11072 7908 11980 7936
rect 11072 7868 11100 7908
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 12986 7936 12992 7948
rect 12947 7908 12992 7936
rect 12986 7896 12992 7908
rect 13044 7896 13050 7948
rect 18966 7896 18972 7948
rect 19024 7936 19030 7948
rect 19061 7939 19119 7945
rect 19061 7936 19073 7939
rect 19024 7908 19073 7936
rect 19024 7896 19030 7908
rect 19061 7905 19073 7908
rect 19107 7905 19119 7939
rect 19061 7899 19119 7905
rect 10888 7840 11100 7868
rect 10229 7831 10287 7837
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11333 7871 11391 7877
rect 11204 7840 11249 7868
rect 11204 7828 11210 7840
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 4120 7772 5580 7800
rect 4120 7760 4126 7772
rect 4617 7735 4675 7741
rect 4617 7701 4629 7735
rect 4663 7732 4675 7735
rect 5442 7732 5448 7744
rect 4663 7704 5448 7732
rect 4663 7701 4675 7704
rect 4617 7695 4675 7701
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 5552 7732 5580 7772
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7009 7803 7067 7809
rect 7009 7800 7021 7803
rect 6972 7772 7021 7800
rect 6972 7760 6978 7772
rect 7009 7769 7021 7772
rect 7055 7769 7067 7803
rect 7009 7763 7067 7769
rect 7190 7760 7196 7812
rect 7248 7800 7254 7812
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 7248 7772 7297 7800
rect 7248 7760 7254 7772
rect 7285 7769 7297 7772
rect 7331 7769 7343 7803
rect 7285 7763 7343 7769
rect 8202 7760 8208 7812
rect 8260 7800 8266 7812
rect 9677 7803 9735 7809
rect 9677 7800 9689 7803
rect 8260 7772 9689 7800
rect 8260 7760 8266 7772
rect 9677 7769 9689 7772
rect 9723 7769 9735 7803
rect 11348 7800 11376 7831
rect 11698 7828 11704 7880
rect 11756 7868 11762 7880
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 11756 7840 13093 7868
rect 11756 7828 11762 7840
rect 13081 7837 13093 7840
rect 13127 7837 13139 7871
rect 13262 7868 13268 7880
rect 13223 7840 13268 7868
rect 13081 7831 13139 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 15838 7868 15844 7880
rect 15799 7840 15844 7868
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 17034 7868 17040 7880
rect 16995 7840 17040 7868
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 18708 7840 19349 7868
rect 12342 7800 12348 7812
rect 11348 7772 12348 7800
rect 9677 7763 9735 7769
rect 12342 7760 12348 7772
rect 12400 7800 12406 7812
rect 13280 7800 13308 7828
rect 12400 7772 13308 7800
rect 15289 7803 15347 7809
rect 12400 7760 12406 7772
rect 15289 7769 15301 7803
rect 15335 7800 15347 7803
rect 16850 7800 16856 7812
rect 15335 7772 16856 7800
rect 15335 7769 15347 7772
rect 15289 7763 15347 7769
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 18598 7800 18604 7812
rect 18511 7772 18604 7800
rect 18598 7760 18604 7772
rect 18656 7800 18662 7812
rect 18708 7800 18736 7840
rect 19337 7837 19349 7840
rect 19383 7868 19395 7871
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 19383 7840 20453 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 20441 7837 20453 7840
rect 20487 7868 20499 7871
rect 20622 7868 20628 7880
rect 20487 7840 20628 7868
rect 20487 7837 20499 7840
rect 20441 7831 20499 7837
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 18656 7772 18736 7800
rect 18656 7760 18662 7772
rect 12526 7732 12532 7744
rect 5552 7704 12532 7732
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 12621 7735 12679 7741
rect 12621 7701 12633 7735
rect 12667 7732 12679 7735
rect 13906 7732 13912 7744
rect 12667 7704 13912 7732
rect 12667 7701 12679 7704
rect 12621 7695 12679 7701
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 15930 7692 15936 7744
rect 15988 7732 15994 7744
rect 17954 7732 17960 7744
rect 15988 7704 17960 7732
rect 15988 7692 15994 7704
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18417 7735 18475 7741
rect 18417 7701 18429 7735
rect 18463 7732 18475 7735
rect 18616 7732 18644 7760
rect 18463 7704 18644 7732
rect 18693 7735 18751 7741
rect 18463 7701 18475 7704
rect 18417 7695 18475 7701
rect 18693 7701 18705 7735
rect 18739 7732 18751 7735
rect 19702 7732 19708 7744
rect 18739 7704 19708 7732
rect 18739 7701 18751 7704
rect 18693 7695 18751 7701
rect 19702 7692 19708 7704
rect 19760 7692 19766 7744
rect 19797 7735 19855 7741
rect 19797 7701 19809 7735
rect 19843 7732 19855 7735
rect 20622 7732 20628 7744
rect 19843 7704 20628 7732
rect 19843 7701 19855 7704
rect 19797 7695 19855 7701
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 5626 7528 5632 7540
rect 3620 7500 5632 7528
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 2317 7327 2375 7333
rect 2317 7324 2329 7327
rect 1636 7296 2329 7324
rect 1636 7284 1642 7296
rect 2317 7293 2329 7296
rect 2363 7293 2375 7327
rect 2317 7287 2375 7293
rect 2584 7327 2642 7333
rect 2584 7293 2596 7327
rect 2630 7324 2642 7327
rect 3326 7324 3332 7336
rect 2630 7296 3332 7324
rect 2630 7293 2642 7296
rect 2584 7287 2642 7293
rect 2332 7256 2360 7287
rect 3326 7284 3332 7296
rect 3384 7284 3390 7336
rect 3620 7256 3648 7500
rect 3697 7463 3755 7469
rect 3697 7429 3709 7463
rect 3743 7429 3755 7463
rect 3970 7460 3976 7472
rect 3931 7432 3976 7460
rect 3697 7423 3755 7429
rect 2332 7228 3648 7256
rect 3712 7392 3740 7423
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 4525 7395 4583 7401
rect 4525 7392 4537 7395
rect 3712 7364 4537 7392
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 3712 7188 3740 7364
rect 4525 7361 4537 7364
rect 4571 7361 4583 7395
rect 4632 7392 4660 7500
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 17678 7528 17684 7540
rect 6012 7500 17684 7528
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4632 7364 4997 7392
rect 4525 7355 4583 7361
rect 4985 7361 4997 7364
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 4341 7327 4399 7333
rect 4341 7324 4353 7327
rect 4304 7296 4353 7324
rect 4304 7284 4310 7296
rect 4341 7293 4353 7296
rect 4387 7293 4399 7327
rect 6012 7324 6040 7500
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 18049 7531 18107 7537
rect 18049 7497 18061 7531
rect 18095 7528 18107 7531
rect 18966 7528 18972 7540
rect 18095 7500 18972 7528
rect 18095 7497 18107 7500
rect 18049 7491 18107 7497
rect 18966 7488 18972 7500
rect 19024 7488 19030 7540
rect 19242 7528 19248 7540
rect 19203 7500 19248 7528
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 20257 7531 20315 7537
rect 20257 7528 20269 7531
rect 19576 7500 20269 7528
rect 19576 7488 19582 7500
rect 20257 7497 20269 7500
rect 20303 7497 20315 7531
rect 20257 7491 20315 7497
rect 9861 7463 9919 7469
rect 9861 7429 9873 7463
rect 9907 7429 9919 7463
rect 9861 7423 9919 7429
rect 4341 7287 4399 7293
rect 4448 7296 6040 7324
rect 6825 7327 6883 7333
rect 4062 7216 4068 7268
rect 4120 7256 4126 7268
rect 4448 7256 4476 7296
rect 6825 7293 6837 7327
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 5258 7265 5264 7268
rect 5252 7256 5264 7265
rect 4120 7228 4476 7256
rect 5219 7228 5264 7256
rect 4120 7216 4126 7228
rect 5252 7219 5264 7228
rect 5258 7216 5264 7219
rect 5316 7216 5322 7268
rect 6840 7256 6868 7287
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7081 7327 7139 7333
rect 7081 7324 7093 7327
rect 6972 7296 7093 7324
rect 6972 7284 6978 7296
rect 7081 7293 7093 7296
rect 7127 7293 7139 7327
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 7081 7287 7139 7293
rect 7576 7296 8493 7324
rect 7576 7268 7604 7296
rect 8481 7293 8493 7296
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 9876 7324 9904 7423
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 19058 7460 19064 7472
rect 13044 7432 19064 7460
rect 13044 7420 13050 7432
rect 19058 7420 19064 7432
rect 19116 7420 19122 7472
rect 19334 7420 19340 7472
rect 19392 7460 19398 7472
rect 19392 7432 20852 7460
rect 19392 7420 19398 7432
rect 17218 7352 17224 7404
rect 17276 7392 17282 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17276 7364 18613 7392
rect 17276 7352 17282 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 19702 7392 19708 7404
rect 19663 7364 19708 7392
rect 18601 7355 18659 7361
rect 19702 7352 19708 7364
rect 19760 7352 19766 7404
rect 19812 7401 19840 7432
rect 19797 7395 19855 7401
rect 19797 7361 19809 7395
rect 19843 7361 19855 7395
rect 19797 7355 19855 7361
rect 19886 7352 19892 7404
rect 19944 7392 19950 7404
rect 20824 7401 20852 7432
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 19944 7364 20729 7392
rect 19944 7352 19950 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 20809 7395 20867 7401
rect 20809 7361 20821 7395
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 8628 7296 9904 7324
rect 18417 7327 18475 7333
rect 8628 7284 8634 7296
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18506 7324 18512 7336
rect 18463 7296 18512 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18506 7284 18512 7296
rect 18564 7324 18570 7336
rect 18966 7324 18972 7336
rect 18564 7296 18972 7324
rect 18564 7284 18570 7296
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 19610 7324 19616 7336
rect 19571 7296 19616 7324
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 20622 7324 20628 7336
rect 20583 7296 20628 7324
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 7558 7256 7564 7268
rect 6840 7228 7564 7256
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 8748 7259 8806 7265
rect 8748 7256 8760 7259
rect 8220 7228 8760 7256
rect 2372 7160 3740 7188
rect 4433 7191 4491 7197
rect 2372 7148 2378 7160
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 5534 7188 5540 7200
rect 4479 7160 5540 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 5718 7148 5724 7200
rect 5776 7188 5782 7200
rect 8220 7197 8248 7228
rect 8748 7225 8760 7228
rect 8794 7256 8806 7259
rect 8846 7256 8852 7268
rect 8794 7228 8852 7256
rect 8794 7225 8806 7228
rect 8748 7219 8806 7225
rect 8846 7216 8852 7228
rect 8904 7216 8910 7268
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 5776 7160 6377 7188
rect 5776 7148 5782 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 8205 7191 8263 7197
rect 8205 7157 8217 7191
rect 8251 7157 8263 7191
rect 8205 7151 8263 7157
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7188 18567 7191
rect 18690 7188 18696 7200
rect 18555 7160 18696 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 18690 7148 18696 7160
rect 18748 7188 18754 7200
rect 18874 7188 18880 7200
rect 18748 7160 18880 7188
rect 18748 7148 18754 7160
rect 18874 7148 18880 7160
rect 18932 7148 18938 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 2832 6956 2877 6984
rect 2832 6944 2838 6956
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 17957 6987 18015 6993
rect 17957 6984 17969 6987
rect 17276 6956 17969 6984
rect 17276 6944 17282 6956
rect 17957 6953 17969 6956
rect 18003 6953 18015 6987
rect 17957 6947 18015 6953
rect 5258 6876 5264 6928
rect 5316 6916 5322 6928
rect 17034 6916 17040 6928
rect 5316 6888 5580 6916
rect 5316 6876 5322 6888
rect 3142 6848 3148 6860
rect 3103 6820 3148 6848
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 3878 6848 3884 6860
rect 3252 6820 3884 6848
rect 3252 6792 3280 6820
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 5040 6820 5365 6848
rect 5040 6808 5046 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 3234 6780 3240 6792
rect 3195 6752 3240 6780
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 3384 6752 3429 6780
rect 3384 6740 3390 6752
rect 5166 6740 5172 6792
rect 5224 6780 5230 6792
rect 5552 6789 5580 6888
rect 16592 6888 17040 6916
rect 5994 6848 6000 6860
rect 5955 6820 6000 6848
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 16592 6857 16620 6888
rect 17034 6876 17040 6888
rect 17092 6916 17098 6928
rect 17092 6888 18828 6916
rect 17092 6876 17098 6888
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6817 16635 6851
rect 16577 6811 16635 6817
rect 16844 6851 16902 6857
rect 16844 6817 16856 6851
rect 16890 6848 16902 6851
rect 16890 6820 18736 6848
rect 16890 6817 16902 6820
rect 16844 6811 16902 6817
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5224 6752 5457 6780
rect 5224 6740 5230 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 4798 6672 4804 6724
rect 4856 6712 4862 6724
rect 14274 6712 14280 6724
rect 4856 6684 14280 6712
rect 4856 6672 4862 6684
rect 14274 6672 14280 6684
rect 14332 6672 14338 6724
rect 4985 6647 5043 6653
rect 4985 6613 4997 6647
rect 5031 6644 5043 6647
rect 5534 6644 5540 6656
rect 5031 6616 5540 6644
rect 5031 6613 5043 6616
rect 4985 6607 5043 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 8938 6604 8944 6656
rect 8996 6644 9002 6656
rect 17954 6644 17960 6656
rect 8996 6616 17960 6644
rect 8996 6604 9002 6616
rect 17954 6604 17960 6616
rect 18012 6604 18018 6656
rect 18708 6644 18736 6820
rect 18800 6792 18828 6888
rect 19052 6851 19110 6857
rect 19052 6817 19064 6851
rect 19098 6848 19110 6851
rect 19426 6848 19432 6860
rect 19098 6820 19432 6848
rect 19098 6817 19110 6820
rect 19052 6811 19110 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 18840 6752 18885 6780
rect 18840 6740 18846 6752
rect 20070 6644 20076 6656
rect 18708 6616 20076 6644
rect 20070 6604 20076 6616
rect 20128 6604 20134 6656
rect 20165 6647 20223 6653
rect 20165 6613 20177 6647
rect 20211 6644 20223 6647
rect 20346 6644 20352 6656
rect 20211 6616 20352 6644
rect 20211 6613 20223 6616
rect 20165 6607 20223 6613
rect 20346 6604 20352 6616
rect 20404 6604 20410 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2961 6443 3019 6449
rect 2961 6409 2973 6443
rect 3007 6440 3019 6443
rect 3050 6440 3056 6452
rect 3007 6412 3056 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 5074 6440 5080 6452
rect 5035 6412 5080 6440
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 18506 6440 18512 6452
rect 12308 6412 18512 6440
rect 12308 6400 12314 6412
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 20070 6400 20076 6452
rect 20128 6440 20134 6452
rect 20438 6440 20444 6452
rect 20128 6412 20444 6440
rect 20128 6400 20134 6412
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 12158 6372 12164 6384
rect 4120 6344 12164 6372
rect 4120 6332 4126 6344
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 1578 6304 1584 6316
rect 1539 6276 1584 6304
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 3142 6264 3148 6316
rect 3200 6304 3206 6316
rect 3237 6307 3295 6313
rect 3237 6304 3249 6307
rect 3200 6276 3249 6304
rect 3200 6264 3206 6276
rect 3237 6273 3249 6276
rect 3283 6273 3295 6307
rect 5534 6304 5540 6316
rect 5495 6276 5540 6304
rect 3237 6267 3295 6273
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 5718 6304 5724 6316
rect 5679 6276 5724 6304
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 13630 6264 13636 6316
rect 13688 6304 13694 6316
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 13688 6276 18521 6304
rect 13688 6264 13694 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 18782 6264 18788 6316
rect 18840 6304 18846 6316
rect 19061 6307 19119 6313
rect 19061 6304 19073 6307
rect 18840 6276 19073 6304
rect 18840 6264 18846 6276
rect 19061 6273 19073 6276
rect 19107 6273 19119 6307
rect 19061 6267 19119 6273
rect 5442 6236 5448 6248
rect 5403 6208 5448 6236
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 18325 6239 18383 6245
rect 18325 6205 18337 6239
rect 18371 6205 18383 6239
rect 18325 6199 18383 6205
rect 1848 6171 1906 6177
rect 1848 6137 1860 6171
rect 1894 6168 1906 6171
rect 2222 6168 2228 6180
rect 1894 6140 2228 6168
rect 1894 6137 1906 6140
rect 1848 6131 1906 6137
rect 2222 6128 2228 6140
rect 2280 6128 2286 6180
rect 18340 6100 18368 6199
rect 19794 6196 19800 6248
rect 19852 6236 19858 6248
rect 20070 6236 20076 6248
rect 19852 6208 20076 6236
rect 19852 6196 19858 6208
rect 20070 6196 20076 6208
rect 20128 6196 20134 6248
rect 19328 6171 19386 6177
rect 19328 6137 19340 6171
rect 19374 6168 19386 6171
rect 20346 6168 20352 6180
rect 19374 6140 20352 6168
rect 19374 6137 19386 6140
rect 19328 6131 19386 6137
rect 20346 6128 20352 6140
rect 20404 6128 20410 6180
rect 19702 6100 19708 6112
rect 18340 6072 19708 6100
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 20530 6060 20536 6112
rect 20588 6100 20594 6112
rect 20717 6103 20775 6109
rect 20717 6100 20729 6103
rect 20588 6072 20729 6100
rect 20588 6060 20594 6072
rect 20717 6069 20729 6072
rect 20763 6069 20775 6103
rect 20717 6063 20775 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 19628 5732 20177 5760
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 19628 5633 19656 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 20254 5692 20260 5704
rect 20215 5664 20260 5692
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20404 5664 20449 5692
rect 20404 5652 20410 5664
rect 19613 5627 19671 5633
rect 19613 5624 19625 5627
rect 4120 5596 19625 5624
rect 4120 5584 4126 5596
rect 19613 5593 19625 5596
rect 19659 5593 19671 5627
rect 19613 5587 19671 5593
rect 19794 5556 19800 5568
rect 19755 5528 19800 5556
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 17954 5352 17960 5364
rect 5960 5324 17960 5352
rect 5960 5312 5966 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 19702 5312 19708 5364
rect 19760 5352 19766 5364
rect 19797 5355 19855 5361
rect 19797 5352 19809 5355
rect 19760 5324 19809 5352
rect 19760 5312 19766 5324
rect 19797 5321 19809 5324
rect 19843 5321 19855 5355
rect 19797 5315 19855 5321
rect 3970 5244 3976 5296
rect 4028 5284 4034 5296
rect 5350 5284 5356 5296
rect 4028 5256 5356 5284
rect 4028 5244 4034 5256
rect 5350 5244 5356 5256
rect 5408 5244 5414 5296
rect 19794 5176 19800 5228
rect 19852 5216 19858 5228
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 19852 5188 20269 5216
rect 19852 5176 19858 5188
rect 20257 5185 20269 5188
rect 20303 5185 20315 5219
rect 20438 5216 20444 5228
rect 20399 5188 20444 5216
rect 20257 5179 20315 5185
rect 20438 5176 20444 5188
rect 20496 5176 20502 5228
rect 20165 5151 20223 5157
rect 20165 5117 20177 5151
rect 20211 5148 20223 5151
rect 20530 5148 20536 5160
rect 20211 5120 20536 5148
rect 20211 5117 20223 5120
rect 20165 5111 20223 5117
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 7466 4128 7472 4140
rect 6788 4100 7472 4128
rect 6788 4088 6794 4100
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 4890 3040 4896 3052
rect 4851 3012 4896 3040
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 20438 3040 20444 3052
rect 5460 3012 20444 3040
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 5460 2972 5488 3012
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 4663 2944 5488 2972
rect 5537 2975 5595 2981
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 5537 2941 5549 2975
rect 5583 2972 5595 2975
rect 11146 2972 11152 2984
rect 5583 2944 11152 2972
rect 5583 2941 5595 2944
rect 5537 2935 5595 2941
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2972 15255 2975
rect 15838 2972 15844 2984
rect 15243 2944 15844 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 15838 2932 15844 2944
rect 15896 2932 15902 2984
rect 5813 2907 5871 2913
rect 5813 2873 5825 2907
rect 5859 2904 5871 2907
rect 6086 2904 6092 2916
rect 5859 2876 6092 2904
rect 5859 2873 5871 2876
rect 5813 2867 5871 2873
rect 6086 2864 6092 2876
rect 6144 2864 6150 2916
rect 9766 2864 9772 2916
rect 9824 2904 9830 2916
rect 15473 2907 15531 2913
rect 15473 2904 15485 2907
rect 9824 2876 15485 2904
rect 9824 2864 9830 2876
rect 15473 2873 15485 2876
rect 15519 2873 15531 2907
rect 15473 2867 15531 2873
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 2958 1164 2964 1216
rect 3016 1204 3022 1216
rect 6270 1204 6276 1216
rect 3016 1176 6276 1204
rect 3016 1164 3022 1176
rect 6270 1164 6276 1176
rect 6328 1164 6334 1216
<< via1 >>
rect 4068 20952 4120 21004
rect 5724 20952 5776 21004
rect 9772 20680 9824 20732
rect 10324 20680 10376 20732
rect 14372 20612 14424 20664
rect 19616 20612 19668 20664
rect 12256 20544 12308 20596
rect 16672 20544 16724 20596
rect 15660 20408 15712 20460
rect 17868 20408 17920 20460
rect 10232 20340 10284 20392
rect 17684 20340 17736 20392
rect 14556 20272 14608 20324
rect 17040 20272 17092 20324
rect 15108 20204 15160 20256
rect 19156 20204 19208 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2780 20000 2832 20052
rect 10232 20043 10284 20052
rect 10232 20009 10241 20043
rect 10241 20009 10275 20043
rect 10275 20009 10284 20043
rect 10232 20000 10284 20009
rect 14372 20000 14424 20052
rect 15108 20000 15160 20052
rect 15660 20043 15712 20052
rect 15660 20009 15669 20043
rect 15669 20009 15703 20043
rect 15703 20009 15712 20043
rect 15660 20000 15712 20009
rect 17500 20000 17552 20052
rect 18512 20043 18564 20052
rect 18512 20009 18521 20043
rect 18521 20009 18555 20043
rect 18555 20009 18564 20043
rect 18512 20000 18564 20009
rect 19064 20043 19116 20052
rect 19064 20009 19073 20043
rect 19073 20009 19107 20043
rect 19107 20009 19116 20043
rect 19064 20000 19116 20009
rect 19248 20000 19300 20052
rect 8484 19932 8536 19984
rect 15568 19932 15620 19984
rect 3700 19864 3752 19916
rect 7748 19864 7800 19916
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 12164 19864 12216 19916
rect 12992 19907 13044 19916
rect 12992 19873 13001 19907
rect 13001 19873 13035 19907
rect 13035 19873 13044 19907
rect 12992 19864 13044 19873
rect 13544 19864 13596 19916
rect 14004 19864 14056 19916
rect 14832 19907 14884 19916
rect 14832 19873 14841 19907
rect 14841 19873 14875 19907
rect 14875 19873 14884 19907
rect 14832 19864 14884 19873
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 16856 19932 16908 19984
rect 16672 19864 16724 19916
rect 18512 19864 18564 19916
rect 19524 19864 19576 19916
rect 20260 19864 20312 19916
rect 4988 19796 5040 19848
rect 7564 19839 7616 19848
rect 7564 19805 7573 19839
rect 7573 19805 7607 19839
rect 7607 19805 7616 19839
rect 7564 19796 7616 19805
rect 9128 19839 9180 19848
rect 6920 19728 6972 19780
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 10232 19796 10284 19848
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 13084 19839 13136 19848
rect 10324 19796 10376 19805
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 14556 19728 14608 19780
rect 18788 19796 18840 19848
rect 18328 19728 18380 19780
rect 19432 19728 19484 19780
rect 20168 19771 20220 19780
rect 20168 19737 20177 19771
rect 20177 19737 20211 19771
rect 20211 19737 20220 19771
rect 20168 19728 20220 19737
rect 2596 19703 2648 19712
rect 2596 19669 2605 19703
rect 2605 19669 2639 19703
rect 2639 19669 2648 19703
rect 2596 19660 2648 19669
rect 7472 19660 7524 19712
rect 9588 19660 9640 19712
rect 12256 19660 12308 19712
rect 13820 19660 13872 19712
rect 13912 19703 13964 19712
rect 13912 19669 13921 19703
rect 13921 19669 13955 19703
rect 13955 19669 13964 19703
rect 13912 19660 13964 19669
rect 17960 19660 18012 19712
rect 20628 19660 20680 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 3516 19499 3568 19508
rect 3516 19465 3525 19499
rect 3525 19465 3559 19499
rect 3559 19465 3568 19499
rect 3516 19456 3568 19465
rect 5724 19499 5776 19508
rect 5724 19465 5733 19499
rect 5733 19465 5767 19499
rect 5767 19465 5776 19499
rect 5724 19456 5776 19465
rect 7564 19456 7616 19508
rect 7932 19456 7984 19508
rect 13084 19456 13136 19508
rect 13912 19456 13964 19508
rect 19616 19499 19668 19508
rect 7748 19388 7800 19440
rect 14832 19388 14884 19440
rect 204 19252 256 19304
rect 2044 19159 2096 19168
rect 2044 19125 2053 19159
rect 2053 19125 2087 19159
rect 2087 19125 2096 19159
rect 2044 19116 2096 19125
rect 2872 19184 2924 19236
rect 10232 19320 10284 19372
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 5172 19252 5224 19304
rect 6092 19252 6144 19304
rect 6184 19252 6236 19304
rect 6828 19252 6880 19304
rect 7012 19295 7064 19304
rect 7012 19261 7021 19295
rect 7021 19261 7055 19295
rect 7055 19261 7064 19295
rect 7012 19252 7064 19261
rect 7564 19184 7616 19236
rect 6368 19116 6420 19168
rect 7288 19116 7340 19168
rect 9588 19295 9640 19304
rect 8116 19184 8168 19236
rect 9312 19184 9364 19236
rect 9588 19261 9597 19295
rect 9597 19261 9631 19295
rect 9631 19261 9640 19295
rect 9588 19252 9640 19261
rect 9772 19252 9824 19304
rect 9956 19252 10008 19304
rect 13268 19320 13320 19372
rect 17500 19363 17552 19372
rect 17500 19329 17509 19363
rect 17509 19329 17543 19363
rect 17543 19329 17552 19363
rect 17500 19320 17552 19329
rect 10968 19252 11020 19304
rect 11060 19252 11112 19304
rect 11980 19252 12032 19304
rect 12256 19252 12308 19304
rect 9680 19184 9732 19236
rect 10416 19184 10468 19236
rect 10784 19184 10836 19236
rect 12808 19184 12860 19236
rect 13820 19252 13872 19304
rect 15108 19252 15160 19304
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 16580 19252 16632 19304
rect 17408 19252 17460 19304
rect 18788 19252 18840 19304
rect 14096 19184 14148 19236
rect 15476 19184 15528 19236
rect 16672 19184 16724 19236
rect 16764 19184 16816 19236
rect 17684 19184 17736 19236
rect 19616 19465 19625 19499
rect 19625 19465 19659 19499
rect 19659 19465 19668 19499
rect 19616 19456 19668 19465
rect 19616 19252 19668 19304
rect 20076 19252 20128 19304
rect 7748 19116 7800 19168
rect 10048 19116 10100 19168
rect 10232 19116 10284 19168
rect 11520 19116 11572 19168
rect 11980 19116 12032 19168
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 12900 19116 12952 19125
rect 13084 19116 13136 19168
rect 15384 19116 15436 19168
rect 15752 19116 15804 19168
rect 16948 19116 17000 19168
rect 17224 19159 17276 19168
rect 17224 19125 17233 19159
rect 17233 19125 17267 19159
rect 17267 19125 17276 19159
rect 17224 19116 17276 19125
rect 18604 19116 18656 19168
rect 22100 19184 22152 19236
rect 20168 19159 20220 19168
rect 20168 19125 20177 19159
rect 20177 19125 20211 19159
rect 20211 19125 20220 19159
rect 20168 19116 20220 19125
rect 20536 19116 20588 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1952 18912 2004 18964
rect 2964 18912 3016 18964
rect 3056 18912 3108 18964
rect 3608 18912 3660 18964
rect 8208 18912 8260 18964
rect 9036 18912 9088 18964
rect 1032 18844 1084 18896
rect 2044 18776 2096 18828
rect 2136 18708 2188 18760
rect 2688 18844 2740 18896
rect 3240 18776 3292 18828
rect 3792 18776 3844 18828
rect 6920 18844 6972 18896
rect 8392 18776 8444 18828
rect 8852 18776 8904 18828
rect 5356 18640 5408 18692
rect 3148 18572 3200 18624
rect 5448 18572 5500 18624
rect 6552 18751 6604 18760
rect 6552 18717 6561 18751
rect 6561 18717 6595 18751
rect 6595 18717 6604 18751
rect 6552 18708 6604 18717
rect 7564 18708 7616 18760
rect 8300 18708 8352 18760
rect 8668 18751 8720 18760
rect 8668 18717 8677 18751
rect 8677 18717 8711 18751
rect 8711 18717 8720 18751
rect 8668 18708 8720 18717
rect 7564 18572 7616 18624
rect 7748 18572 7800 18624
rect 8208 18615 8260 18624
rect 8208 18581 8217 18615
rect 8217 18581 8251 18615
rect 8251 18581 8260 18615
rect 8208 18572 8260 18581
rect 8392 18640 8444 18692
rect 10784 18912 10836 18964
rect 10968 18912 11020 18964
rect 11520 18912 11572 18964
rect 12716 18912 12768 18964
rect 13176 18912 13228 18964
rect 17408 18912 17460 18964
rect 17500 18912 17552 18964
rect 10048 18844 10100 18896
rect 10324 18844 10376 18896
rect 11980 18887 12032 18896
rect 11980 18853 12014 18887
rect 12014 18853 12032 18887
rect 11980 18844 12032 18853
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 10416 18776 10468 18828
rect 15568 18844 15620 18896
rect 16948 18844 17000 18896
rect 14188 18776 14240 18828
rect 15752 18776 15804 18828
rect 17040 18776 17092 18828
rect 17960 18844 18012 18896
rect 18696 18844 18748 18896
rect 18972 18776 19024 18828
rect 19708 18776 19760 18828
rect 11520 18708 11572 18760
rect 12716 18708 12768 18760
rect 13176 18708 13228 18760
rect 19340 18751 19392 18760
rect 14740 18683 14792 18692
rect 14740 18649 14749 18683
rect 14749 18649 14783 18683
rect 14783 18649 14792 18683
rect 19340 18717 19349 18751
rect 19349 18717 19383 18751
rect 19383 18717 19392 18751
rect 19340 18708 19392 18717
rect 19984 18708 20036 18760
rect 20720 18708 20772 18760
rect 14740 18640 14792 18649
rect 18788 18640 18840 18692
rect 9588 18572 9640 18624
rect 9864 18572 9916 18624
rect 14464 18572 14516 18624
rect 15660 18572 15712 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2780 18368 2832 18420
rect 2228 18300 2280 18352
rect 3516 18368 3568 18420
rect 3976 18300 4028 18352
rect 1860 18232 1912 18284
rect 8668 18368 8720 18420
rect 9128 18368 9180 18420
rect 9588 18368 9640 18420
rect 10416 18368 10468 18420
rect 11152 18368 11204 18420
rect 11704 18368 11756 18420
rect 12992 18368 13044 18420
rect 13176 18368 13228 18420
rect 15016 18368 15068 18420
rect 8576 18300 8628 18352
rect 10876 18300 10928 18352
rect 12716 18300 12768 18352
rect 12900 18300 12952 18352
rect 6092 18275 6144 18284
rect 6092 18241 6101 18275
rect 6101 18241 6135 18275
rect 6135 18241 6144 18275
rect 6092 18232 6144 18241
rect 6552 18232 6604 18284
rect 8484 18275 8536 18284
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 2964 18164 3016 18216
rect 3884 18164 3936 18216
rect 6736 18164 6788 18216
rect 4804 18096 4856 18148
rect 5356 18096 5408 18148
rect 1400 18028 1452 18080
rect 2872 18028 2924 18080
rect 3608 18071 3660 18080
rect 3608 18037 3617 18071
rect 3617 18037 3651 18071
rect 3651 18037 3660 18071
rect 3608 18028 3660 18037
rect 5908 18028 5960 18080
rect 8484 18241 8493 18275
rect 8493 18241 8527 18275
rect 8527 18241 8536 18275
rect 8484 18232 8536 18241
rect 10048 18275 10100 18284
rect 10048 18241 10057 18275
rect 10057 18241 10091 18275
rect 10091 18241 10100 18275
rect 10048 18232 10100 18241
rect 10140 18232 10192 18284
rect 13268 18232 13320 18284
rect 11796 18164 11848 18216
rect 11980 18164 12032 18216
rect 14740 18164 14792 18216
rect 9220 18096 9272 18148
rect 10600 18096 10652 18148
rect 11152 18096 11204 18148
rect 13084 18096 13136 18148
rect 13176 18096 13228 18148
rect 13636 18096 13688 18148
rect 15016 18096 15068 18148
rect 6920 18028 6972 18080
rect 8300 18028 8352 18080
rect 9312 18028 9364 18080
rect 9772 18028 9824 18080
rect 10048 18028 10100 18080
rect 11428 18071 11480 18080
rect 11428 18037 11437 18071
rect 11437 18037 11471 18071
rect 11471 18037 11480 18071
rect 11428 18028 11480 18037
rect 12992 18071 13044 18080
rect 12992 18037 13001 18071
rect 13001 18037 13035 18071
rect 13035 18037 13044 18071
rect 17040 18368 17092 18420
rect 17776 18368 17828 18420
rect 19524 18368 19576 18420
rect 19708 18411 19760 18420
rect 19708 18377 19717 18411
rect 19717 18377 19751 18411
rect 19751 18377 19760 18411
rect 19708 18368 19760 18377
rect 19248 18232 19300 18284
rect 15752 18207 15804 18216
rect 15752 18173 15761 18207
rect 15761 18173 15795 18207
rect 15795 18173 15804 18207
rect 15752 18164 15804 18173
rect 16304 18164 16356 18216
rect 17960 18164 18012 18216
rect 18604 18164 18656 18216
rect 18788 18164 18840 18216
rect 20996 18164 21048 18216
rect 15844 18096 15896 18148
rect 17500 18096 17552 18148
rect 20812 18096 20864 18148
rect 12992 18028 13044 18037
rect 19248 18028 19300 18080
rect 20628 18028 20680 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 3516 17824 3568 17876
rect 7012 17824 7064 17876
rect 7472 17867 7524 17876
rect 7472 17833 7481 17867
rect 7481 17833 7515 17867
rect 7515 17833 7524 17867
rect 7472 17824 7524 17833
rect 8208 17824 8260 17876
rect 8392 17824 8444 17876
rect 9864 17867 9916 17876
rect 9864 17833 9873 17867
rect 9873 17833 9907 17867
rect 9907 17833 9916 17867
rect 9864 17824 9916 17833
rect 11428 17824 11480 17876
rect 13268 17824 13320 17876
rect 14556 17824 14608 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15660 17867 15712 17876
rect 15660 17833 15669 17867
rect 15669 17833 15703 17867
rect 15703 17833 15712 17867
rect 15660 17824 15712 17833
rect 16764 17824 16816 17876
rect 16948 17824 17000 17876
rect 17224 17824 17276 17876
rect 20720 17824 20772 17876
rect 20812 17824 20864 17876
rect 2320 17756 2372 17808
rect 9588 17756 9640 17808
rect 1676 17731 1728 17740
rect 1676 17697 1685 17731
rect 1685 17697 1719 17731
rect 1719 17697 1728 17731
rect 1676 17688 1728 17697
rect 2136 17620 2188 17672
rect 3332 17688 3384 17740
rect 5080 17731 5132 17740
rect 5080 17697 5089 17731
rect 5089 17697 5123 17731
rect 5123 17697 5132 17731
rect 5080 17688 5132 17697
rect 7012 17620 7064 17672
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 8484 17731 8536 17740
rect 8484 17697 8493 17731
rect 8493 17697 8527 17731
rect 8527 17697 8536 17731
rect 8484 17688 8536 17697
rect 8944 17620 8996 17672
rect 9128 17688 9180 17740
rect 10232 17688 10284 17740
rect 10968 17688 11020 17740
rect 11888 17688 11940 17740
rect 12716 17688 12768 17740
rect 14924 17688 14976 17740
rect 10048 17620 10100 17672
rect 10324 17620 10376 17672
rect 12624 17663 12676 17672
rect 12624 17629 12633 17663
rect 12633 17629 12667 17663
rect 12667 17629 12676 17663
rect 12624 17620 12676 17629
rect 5816 17552 5868 17604
rect 1768 17484 1820 17536
rect 3332 17484 3384 17536
rect 3424 17484 3476 17536
rect 6920 17484 6972 17536
rect 7196 17484 7248 17536
rect 9312 17552 9364 17604
rect 10232 17552 10284 17604
rect 11796 17595 11848 17604
rect 11796 17561 11805 17595
rect 11805 17561 11839 17595
rect 11839 17561 11848 17595
rect 11796 17552 11848 17561
rect 12164 17552 12216 17604
rect 13636 17620 13688 17672
rect 15016 17620 15068 17672
rect 17132 17688 17184 17740
rect 18512 17688 18564 17740
rect 19248 17756 19300 17808
rect 21732 17756 21784 17808
rect 20260 17731 20312 17740
rect 20260 17697 20269 17731
rect 20269 17697 20303 17731
rect 20303 17697 20312 17731
rect 20260 17688 20312 17697
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 12256 17484 12308 17536
rect 13452 17484 13504 17536
rect 17040 17663 17092 17672
rect 17040 17629 17049 17663
rect 17049 17629 17083 17663
rect 17083 17629 17092 17663
rect 17040 17620 17092 17629
rect 18604 17663 18656 17672
rect 18604 17629 18613 17663
rect 18613 17629 18647 17663
rect 18647 17629 18656 17663
rect 18604 17620 18656 17629
rect 18788 17484 18840 17536
rect 19800 17484 19852 17536
rect 19984 17527 20036 17536
rect 19984 17493 19993 17527
rect 19993 17493 20027 17527
rect 20027 17493 20036 17527
rect 19984 17484 20036 17493
rect 20444 17527 20496 17536
rect 20444 17493 20453 17527
rect 20453 17493 20487 17527
rect 20487 17493 20496 17527
rect 20444 17484 20496 17493
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 2780 17280 2832 17332
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 3148 17280 3200 17332
rect 5080 17280 5132 17332
rect 5816 17280 5868 17332
rect 8024 17280 8076 17332
rect 2872 17212 2924 17264
rect 10784 17280 10836 17332
rect 11152 17280 11204 17332
rect 4712 17144 4764 17196
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 6920 17144 6972 17196
rect 7472 17187 7524 17196
rect 1860 17076 1912 17128
rect 3424 17119 3476 17128
rect 2412 17008 2464 17060
rect 3424 17085 3433 17119
rect 3433 17085 3467 17119
rect 3467 17085 3476 17119
rect 3424 17076 3476 17085
rect 6276 17076 6328 17128
rect 7196 17119 7248 17128
rect 7196 17085 7205 17119
rect 7205 17085 7239 17119
rect 7239 17085 7248 17119
rect 7196 17076 7248 17085
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 7564 17144 7616 17196
rect 8944 17144 8996 17196
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 4804 16983 4856 16992
rect 4804 16949 4813 16983
rect 4813 16949 4847 16983
rect 4847 16949 4856 16983
rect 4804 16940 4856 16949
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 5816 16983 5868 16992
rect 4896 16940 4948 16949
rect 5816 16949 5825 16983
rect 5825 16949 5859 16983
rect 5859 16949 5868 16983
rect 5816 16940 5868 16949
rect 6828 16983 6880 16992
rect 6828 16949 6837 16983
rect 6837 16949 6871 16983
rect 6871 16949 6880 16983
rect 6828 16940 6880 16949
rect 8668 17076 8720 17128
rect 9680 17076 9732 17128
rect 10968 17212 11020 17264
rect 12624 17280 12676 17332
rect 17868 17280 17920 17332
rect 9864 17144 9916 17196
rect 11060 17144 11112 17196
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 14188 17212 14240 17264
rect 12808 17144 12860 17196
rect 13728 17187 13780 17196
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 13728 17144 13780 17153
rect 13452 17119 13504 17128
rect 8300 17008 8352 17060
rect 10968 17008 11020 17060
rect 8576 16940 8628 16992
rect 8668 16940 8720 16992
rect 10232 16940 10284 16992
rect 10784 16940 10836 16992
rect 11428 17008 11480 17060
rect 13452 17085 13461 17119
rect 13461 17085 13495 17119
rect 13495 17085 13504 17119
rect 13452 17076 13504 17085
rect 14556 17212 14608 17264
rect 16028 17144 16080 17196
rect 11244 16983 11296 16992
rect 11244 16949 11253 16983
rect 11253 16949 11287 16983
rect 11287 16949 11296 16983
rect 11244 16940 11296 16949
rect 11888 16940 11940 16992
rect 13084 16983 13136 16992
rect 13084 16949 13093 16983
rect 13093 16949 13127 16983
rect 13127 16949 13136 16983
rect 13084 16940 13136 16949
rect 13912 17008 13964 17060
rect 14004 17008 14056 17060
rect 14924 17008 14976 17060
rect 15200 17008 15252 17060
rect 17500 17212 17552 17264
rect 19156 17212 19208 17264
rect 20996 17212 21048 17264
rect 16580 17187 16632 17196
rect 16580 17153 16589 17187
rect 16589 17153 16623 17187
rect 16623 17153 16632 17187
rect 16580 17144 16632 17153
rect 16856 17076 16908 17128
rect 18328 17144 18380 17196
rect 18880 17144 18932 17196
rect 19248 17144 19300 17196
rect 13636 16940 13688 16992
rect 14096 16940 14148 16992
rect 15568 16940 15620 16992
rect 19524 17076 19576 17128
rect 20536 17119 20588 17128
rect 20536 17085 20545 17119
rect 20545 17085 20579 17119
rect 20579 17085 20588 17119
rect 20536 17076 20588 17085
rect 17224 17008 17276 17060
rect 17960 17008 18012 17060
rect 19156 16940 19208 16992
rect 19524 16983 19576 16992
rect 19524 16949 19533 16983
rect 19533 16949 19567 16983
rect 19567 16949 19576 16983
rect 19524 16940 19576 16949
rect 19708 16940 19760 16992
rect 20352 16940 20404 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 3240 16736 3292 16788
rect 5540 16736 5592 16788
rect 572 16668 624 16720
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 2872 16600 2924 16652
rect 4712 16668 4764 16720
rect 6828 16736 6880 16788
rect 6000 16668 6052 16720
rect 7472 16668 7524 16720
rect 8576 16736 8628 16788
rect 10508 16736 10560 16788
rect 15016 16736 15068 16788
rect 17500 16736 17552 16788
rect 17868 16779 17920 16788
rect 17868 16745 17877 16779
rect 17877 16745 17911 16779
rect 17911 16745 17920 16779
rect 17868 16736 17920 16745
rect 18604 16779 18656 16788
rect 18604 16745 18613 16779
rect 18613 16745 18647 16779
rect 18647 16745 18656 16779
rect 18604 16736 18656 16745
rect 18880 16736 18932 16788
rect 10232 16668 10284 16720
rect 13912 16668 13964 16720
rect 14648 16668 14700 16720
rect 18328 16668 18380 16720
rect 3332 16532 3384 16584
rect 3608 16532 3660 16584
rect 5540 16532 5592 16584
rect 5908 16575 5960 16584
rect 5908 16541 5917 16575
rect 5917 16541 5951 16575
rect 5951 16541 5960 16575
rect 5908 16532 5960 16541
rect 7196 16600 7248 16652
rect 8300 16600 8352 16652
rect 8392 16600 8444 16652
rect 10324 16600 10376 16652
rect 1952 16507 2004 16516
rect 1952 16473 1961 16507
rect 1961 16473 1995 16507
rect 1995 16473 2004 16507
rect 1952 16464 2004 16473
rect 9036 16532 9088 16584
rect 11244 16600 11296 16652
rect 13084 16600 13136 16652
rect 15108 16600 15160 16652
rect 15752 16600 15804 16652
rect 15936 16600 15988 16652
rect 19064 16600 19116 16652
rect 19248 16643 19300 16652
rect 19248 16609 19282 16643
rect 19282 16609 19300 16643
rect 19248 16600 19300 16609
rect 12164 16575 12216 16584
rect 2044 16396 2096 16448
rect 7288 16439 7340 16448
rect 7288 16405 7297 16439
rect 7297 16405 7331 16439
rect 7331 16405 7340 16439
rect 9680 16507 9732 16516
rect 9680 16473 9689 16507
rect 9689 16473 9723 16507
rect 9723 16473 9732 16507
rect 9680 16464 9732 16473
rect 11060 16464 11112 16516
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 12164 16532 12216 16541
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 13636 16575 13688 16584
rect 12256 16532 12308 16541
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 14556 16575 14608 16584
rect 14556 16541 14565 16575
rect 14565 16541 14599 16575
rect 14599 16541 14608 16575
rect 14556 16532 14608 16541
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 18788 16532 18840 16584
rect 14004 16507 14056 16516
rect 7288 16396 7340 16405
rect 12348 16396 12400 16448
rect 14004 16473 14013 16507
rect 14013 16473 14047 16507
rect 14047 16473 14056 16507
rect 14004 16464 14056 16473
rect 14280 16396 14332 16448
rect 14648 16396 14700 16448
rect 17776 16396 17828 16448
rect 17868 16396 17920 16448
rect 19984 16396 20036 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 4804 16192 4856 16244
rect 5264 16192 5316 16244
rect 5724 16192 5776 16244
rect 5908 16192 5960 16244
rect 7472 16192 7524 16244
rect 9404 16192 9456 16244
rect 10324 16192 10376 16244
rect 12164 16192 12216 16244
rect 12348 16192 12400 16244
rect 15568 16192 15620 16244
rect 16028 16235 16080 16244
rect 16028 16201 16037 16235
rect 16037 16201 16071 16235
rect 16071 16201 16080 16235
rect 16028 16192 16080 16201
rect 16212 16192 16264 16244
rect 16856 16235 16908 16244
rect 16856 16201 16865 16235
rect 16865 16201 16899 16235
rect 16899 16201 16908 16235
rect 16856 16192 16908 16201
rect 17040 16192 17092 16244
rect 4712 16124 4764 16176
rect 5172 16124 5224 16176
rect 5264 16056 5316 16108
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 3056 16031 3108 16040
rect 3056 15997 3065 16031
rect 3065 15997 3099 16031
rect 3099 15997 3108 16031
rect 3056 15988 3108 15997
rect 3608 15988 3660 16040
rect 5448 16031 5500 16040
rect 5448 15997 5457 16031
rect 5457 15997 5491 16031
rect 5491 15997 5500 16031
rect 5448 15988 5500 15997
rect 8484 16056 8536 16108
rect 11336 16124 11388 16176
rect 12900 16124 12952 16176
rect 11060 16056 11112 16108
rect 11704 16056 11756 16108
rect 11980 16056 12032 16108
rect 14004 16056 14056 16108
rect 3148 15920 3200 15972
rect 3424 15920 3476 15972
rect 3976 15920 4028 15972
rect 6644 15920 6696 15972
rect 1952 15895 2004 15904
rect 1952 15861 1961 15895
rect 1961 15861 1995 15895
rect 1995 15861 2004 15895
rect 1952 15852 2004 15861
rect 2504 15895 2556 15904
rect 2504 15861 2513 15895
rect 2513 15861 2547 15895
rect 2547 15861 2556 15895
rect 2504 15852 2556 15861
rect 5080 15852 5132 15904
rect 6920 15988 6972 16040
rect 9036 16031 9088 16040
rect 9036 15997 9070 16031
rect 9070 15997 9088 16031
rect 9036 15988 9088 15997
rect 10968 16031 11020 16040
rect 10968 15997 10977 16031
rect 10977 15997 11011 16031
rect 11011 15997 11020 16031
rect 10968 15988 11020 15997
rect 12348 15988 12400 16040
rect 7288 15920 7340 15972
rect 8944 15920 8996 15972
rect 9312 15920 9364 15972
rect 10232 15920 10284 15972
rect 10784 15920 10836 15972
rect 13636 15988 13688 16040
rect 13912 15920 13964 15972
rect 7196 15852 7248 15904
rect 8484 15895 8536 15904
rect 8484 15861 8493 15895
rect 8493 15861 8527 15895
rect 8527 15861 8536 15895
rect 8484 15852 8536 15861
rect 12900 15852 12952 15904
rect 17224 15988 17276 16040
rect 18052 16056 18104 16108
rect 19248 16192 19300 16244
rect 18420 15988 18472 16040
rect 18788 15988 18840 16040
rect 14556 15920 14608 15972
rect 15200 15920 15252 15972
rect 17040 15920 17092 15972
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 14372 15852 14424 15861
rect 18604 15920 18656 15972
rect 19616 15920 19668 15972
rect 19984 15988 20036 16040
rect 21088 15988 21140 16040
rect 20168 15920 20220 15972
rect 20996 15920 21048 15972
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 18512 15895 18564 15904
rect 17316 15852 17368 15861
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 18512 15852 18564 15861
rect 20628 15852 20680 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 3240 15691 3292 15700
rect 3240 15657 3249 15691
rect 3249 15657 3283 15691
rect 3283 15657 3292 15691
rect 3240 15648 3292 15657
rect 3516 15580 3568 15632
rect 5540 15648 5592 15700
rect 5816 15648 5868 15700
rect 11888 15648 11940 15700
rect 6644 15580 6696 15632
rect 8668 15580 8720 15632
rect 3608 15512 3660 15564
rect 4988 15555 5040 15564
rect 4988 15521 4997 15555
rect 4997 15521 5031 15555
rect 5031 15521 5040 15555
rect 4988 15512 5040 15521
rect 5172 15512 5224 15564
rect 3424 15487 3476 15496
rect 3424 15453 3433 15487
rect 3433 15453 3467 15487
rect 3467 15453 3476 15487
rect 5264 15487 5316 15496
rect 3424 15444 3476 15453
rect 4896 15376 4948 15428
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 8300 15512 8352 15564
rect 11336 15580 11388 15632
rect 12348 15648 12400 15700
rect 14280 15648 14332 15700
rect 10876 15555 10928 15564
rect 10876 15521 10910 15555
rect 10910 15521 10928 15555
rect 10876 15512 10928 15521
rect 16028 15580 16080 15632
rect 14280 15555 14332 15564
rect 7564 15487 7616 15496
rect 7564 15453 7573 15487
rect 7573 15453 7607 15487
rect 7607 15453 7616 15487
rect 7564 15444 7616 15453
rect 8944 15444 8996 15496
rect 8392 15376 8444 15428
rect 1952 15351 2004 15360
rect 1952 15317 1961 15351
rect 1961 15317 1995 15351
rect 1995 15317 2004 15351
rect 1952 15308 2004 15317
rect 2320 15308 2372 15360
rect 3976 15308 4028 15360
rect 4160 15308 4212 15360
rect 6276 15308 6328 15360
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 15936 15512 15988 15564
rect 17960 15648 18012 15700
rect 17500 15623 17552 15632
rect 17500 15589 17509 15623
rect 17509 15589 17543 15623
rect 17543 15589 17552 15623
rect 18696 15648 18748 15700
rect 19524 15648 19576 15700
rect 17500 15580 17552 15589
rect 19708 15580 19760 15632
rect 20536 15580 20588 15632
rect 16580 15376 16632 15428
rect 12624 15308 12676 15360
rect 13636 15351 13688 15360
rect 13636 15317 13645 15351
rect 13645 15317 13679 15351
rect 13679 15317 13688 15351
rect 13636 15308 13688 15317
rect 15752 15308 15804 15360
rect 17040 15351 17092 15360
rect 17040 15317 17049 15351
rect 17049 15317 17083 15351
rect 17083 15317 17092 15351
rect 17040 15308 17092 15317
rect 17224 15308 17276 15360
rect 17592 15308 17644 15360
rect 19340 15512 19392 15564
rect 19892 15512 19944 15564
rect 20076 15555 20128 15564
rect 20076 15521 20085 15555
rect 20085 15521 20119 15555
rect 20119 15521 20128 15555
rect 20076 15512 20128 15521
rect 19248 15444 19300 15496
rect 17776 15376 17828 15428
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 18880 15308 18932 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 7012 15104 7064 15156
rect 8300 15104 8352 15156
rect 10876 15104 10928 15156
rect 11888 15104 11940 15156
rect 3424 15036 3476 15088
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 3056 14900 3108 14952
rect 3976 14900 4028 14952
rect 4988 14968 5040 15020
rect 6644 14968 6696 15020
rect 7012 14968 7064 15020
rect 7196 14968 7248 15020
rect 8760 14968 8812 15020
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 9680 15036 9732 15088
rect 14280 15104 14332 15156
rect 14096 15079 14148 15088
rect 11704 14968 11756 15020
rect 14096 15045 14105 15079
rect 14105 15045 14139 15079
rect 14139 15045 14148 15079
rect 14096 15036 14148 15045
rect 13820 15011 13872 15020
rect 5448 14900 5500 14952
rect 6276 14900 6328 14952
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 3240 14832 3292 14884
rect 4252 14832 4304 14884
rect 8668 14832 8720 14884
rect 8944 14832 8996 14884
rect 11704 14875 11756 14884
rect 11704 14841 11713 14875
rect 11713 14841 11747 14875
rect 11747 14841 11756 14875
rect 11704 14832 11756 14841
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 4712 14764 4764 14816
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 8300 14764 8352 14816
rect 9036 14764 9088 14816
rect 11520 14764 11572 14816
rect 11796 14807 11848 14816
rect 11796 14773 11805 14807
rect 11805 14773 11839 14807
rect 11839 14773 11848 14807
rect 11796 14764 11848 14773
rect 12992 14832 13044 14884
rect 17592 15036 17644 15088
rect 14372 14968 14424 15020
rect 15844 14968 15896 15020
rect 18052 15036 18104 15088
rect 19616 15104 19668 15156
rect 15016 14900 15068 14952
rect 13912 14832 13964 14884
rect 15844 14764 15896 14816
rect 16028 14764 16080 14816
rect 16580 14943 16632 14952
rect 16580 14909 16614 14943
rect 16614 14909 16632 14943
rect 16580 14900 16632 14909
rect 17500 14832 17552 14884
rect 19064 14968 19116 15020
rect 18788 14900 18840 14952
rect 17960 14832 18012 14884
rect 17868 14764 17920 14816
rect 18696 14764 18748 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1676 14560 1728 14612
rect 4160 14560 4212 14612
rect 4620 14560 4672 14612
rect 4712 14603 4764 14612
rect 4712 14569 4721 14603
rect 4721 14569 4755 14603
rect 4755 14569 4764 14603
rect 4712 14560 4764 14569
rect 6920 14560 6972 14612
rect 3332 14492 3384 14544
rect 6092 14492 6144 14544
rect 7104 14492 7156 14544
rect 1676 14424 1728 14476
rect 3608 14424 3660 14476
rect 3976 14424 4028 14476
rect 5448 14424 5500 14476
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 8116 14424 8168 14476
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 2780 14356 2832 14408
rect 3424 14399 3476 14408
rect 2964 14288 3016 14340
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 4804 14356 4856 14408
rect 7012 14356 7064 14408
rect 9772 14560 9824 14612
rect 10232 14492 10284 14544
rect 11704 14560 11756 14612
rect 12532 14560 12584 14612
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 15108 14560 15160 14612
rect 17868 14560 17920 14612
rect 17960 14560 18012 14612
rect 18880 14603 18932 14612
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 20076 14560 20128 14612
rect 11060 14424 11112 14476
rect 16120 14492 16172 14544
rect 12440 14424 12492 14476
rect 12992 14424 13044 14476
rect 14096 14467 14148 14476
rect 14096 14433 14105 14467
rect 14105 14433 14139 14467
rect 14139 14433 14148 14467
rect 14096 14424 14148 14433
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 17776 14492 17828 14544
rect 20168 14492 20220 14544
rect 17592 14424 17644 14476
rect 18696 14467 18748 14476
rect 18696 14433 18705 14467
rect 18705 14433 18739 14467
rect 18739 14433 18748 14467
rect 18696 14424 18748 14433
rect 20076 14424 20128 14476
rect 10784 14356 10836 14408
rect 10876 14356 10928 14408
rect 3516 14220 3568 14272
rect 12716 14356 12768 14408
rect 7564 14220 7616 14272
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 11980 14220 12032 14272
rect 12624 14220 12676 14272
rect 12900 14263 12952 14272
rect 12900 14229 12909 14263
rect 12909 14229 12943 14263
rect 12943 14229 12952 14263
rect 12900 14220 12952 14229
rect 13820 14356 13872 14408
rect 15476 14288 15528 14340
rect 16028 14356 16080 14408
rect 19340 14356 19392 14408
rect 19800 14399 19852 14408
rect 19800 14365 19809 14399
rect 19809 14365 19843 14399
rect 19843 14365 19852 14399
rect 19800 14356 19852 14365
rect 18696 14288 18748 14340
rect 16304 14220 16356 14272
rect 17684 14220 17736 14272
rect 20444 14263 20496 14272
rect 20444 14229 20453 14263
rect 20453 14229 20487 14263
rect 20487 14229 20496 14263
rect 20444 14220 20496 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 1676 14059 1728 14068
rect 1676 14025 1685 14059
rect 1685 14025 1719 14059
rect 1719 14025 1728 14059
rect 1676 14016 1728 14025
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 5540 14016 5592 14068
rect 8116 14016 8168 14068
rect 8392 14059 8444 14068
rect 8392 14025 8401 14059
rect 8401 14025 8435 14059
rect 8435 14025 8444 14059
rect 8392 14016 8444 14025
rect 4804 13948 4856 14000
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 9588 14016 9640 14068
rect 10876 14059 10928 14068
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 2688 13855 2740 13864
rect 2688 13821 2697 13855
rect 2697 13821 2731 13855
rect 2731 13821 2740 13855
rect 2688 13812 2740 13821
rect 3976 13812 4028 13864
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 7564 13812 7616 13864
rect 10232 13880 10284 13932
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 10784 13948 10836 14000
rect 12716 14016 12768 14068
rect 13084 14016 13136 14068
rect 15936 14016 15988 14068
rect 16028 14016 16080 14068
rect 16488 14016 16540 14068
rect 17316 14016 17368 14068
rect 18604 14016 18656 14068
rect 19340 14059 19392 14068
rect 19340 14025 19349 14059
rect 19349 14025 19383 14059
rect 19383 14025 19392 14059
rect 19340 14016 19392 14025
rect 19984 14016 20036 14068
rect 20168 14016 20220 14068
rect 11428 13923 11480 13932
rect 11428 13889 11437 13923
rect 11437 13889 11471 13923
rect 11471 13889 11480 13923
rect 11428 13880 11480 13889
rect 11704 13880 11756 13932
rect 12532 13812 12584 13864
rect 12716 13855 12768 13864
rect 12716 13821 12750 13855
rect 12750 13821 12768 13855
rect 12716 13812 12768 13821
rect 3516 13787 3568 13796
rect 3516 13753 3550 13787
rect 3550 13753 3568 13787
rect 3516 13744 3568 13753
rect 9404 13787 9456 13796
rect 9404 13753 9413 13787
rect 9413 13753 9447 13787
rect 9447 13753 9456 13787
rect 9404 13744 9456 13753
rect 11520 13744 11572 13796
rect 14188 13812 14240 13864
rect 17132 13948 17184 14000
rect 16304 13923 16356 13932
rect 15384 13812 15436 13864
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16304 13880 16356 13889
rect 17040 13880 17092 13932
rect 17592 13923 17644 13932
rect 17592 13889 17601 13923
rect 17601 13889 17635 13923
rect 17635 13889 17644 13923
rect 17592 13880 17644 13889
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 19432 13880 19484 13932
rect 14372 13787 14424 13796
rect 1768 13676 1820 13728
rect 9036 13719 9088 13728
rect 9036 13685 9045 13719
rect 9045 13685 9079 13719
rect 9079 13685 9088 13719
rect 9036 13676 9088 13685
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 10508 13676 10560 13728
rect 13728 13676 13780 13728
rect 14372 13753 14406 13787
rect 14406 13753 14424 13787
rect 14372 13744 14424 13753
rect 16120 13812 16172 13864
rect 16396 13744 16448 13796
rect 18696 13744 18748 13796
rect 19616 13744 19668 13796
rect 15292 13676 15344 13728
rect 15476 13719 15528 13728
rect 15476 13685 15485 13719
rect 15485 13685 15519 13719
rect 15519 13685 15528 13719
rect 15476 13676 15528 13685
rect 15752 13719 15804 13728
rect 15752 13685 15761 13719
rect 15761 13685 15795 13719
rect 15795 13685 15804 13719
rect 15752 13676 15804 13685
rect 16028 13676 16080 13728
rect 18788 13676 18840 13728
rect 19708 13719 19760 13728
rect 19708 13685 19717 13719
rect 19717 13685 19751 13719
rect 19751 13685 19760 13719
rect 19708 13676 19760 13685
rect 19984 13676 20036 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 2228 13515 2280 13524
rect 2228 13481 2237 13515
rect 2237 13481 2271 13515
rect 2271 13481 2280 13515
rect 2228 13472 2280 13481
rect 6092 13515 6144 13524
rect 2688 13404 2740 13456
rect 1492 13379 1544 13388
rect 1492 13345 1501 13379
rect 1501 13345 1535 13379
rect 1535 13345 1544 13379
rect 1492 13336 1544 13345
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 3148 13404 3200 13456
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 9036 13472 9088 13524
rect 11428 13472 11480 13524
rect 12624 13472 12676 13524
rect 12900 13472 12952 13524
rect 7104 13404 7156 13456
rect 7564 13404 7616 13456
rect 8024 13404 8076 13456
rect 10048 13404 10100 13456
rect 2964 13336 3016 13388
rect 4160 13336 4212 13388
rect 4988 13336 5040 13388
rect 5172 13336 5224 13388
rect 5540 13336 5592 13388
rect 6920 13336 6972 13388
rect 7472 13379 7524 13388
rect 7472 13345 7481 13379
rect 7481 13345 7515 13379
rect 7515 13345 7524 13379
rect 7472 13336 7524 13345
rect 6644 13311 6696 13320
rect 2320 13132 2372 13184
rect 2688 13132 2740 13184
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 6736 13268 6788 13320
rect 7840 13336 7892 13388
rect 8392 13268 8444 13320
rect 9680 13336 9732 13388
rect 11520 13336 11572 13388
rect 11704 13379 11756 13388
rect 11704 13345 11738 13379
rect 11738 13345 11756 13379
rect 11704 13336 11756 13345
rect 11980 13404 12032 13456
rect 15292 13404 15344 13456
rect 16396 13472 16448 13524
rect 16488 13472 16540 13524
rect 16580 13404 16632 13456
rect 16672 13336 16724 13388
rect 16948 13472 17000 13524
rect 18696 13472 18748 13524
rect 19800 13472 19852 13524
rect 20444 13515 20496 13524
rect 20444 13481 20453 13515
rect 20453 13481 20487 13515
rect 20487 13481 20496 13515
rect 20444 13472 20496 13481
rect 19432 13404 19484 13456
rect 18512 13336 18564 13388
rect 18696 13336 18748 13388
rect 19892 13336 19944 13388
rect 20812 13336 20864 13388
rect 5172 13200 5224 13252
rect 8116 13200 8168 13252
rect 9772 13200 9824 13252
rect 4712 13132 4764 13184
rect 5724 13132 5776 13184
rect 6644 13132 6696 13184
rect 8300 13132 8352 13184
rect 12624 13268 12676 13320
rect 13360 13268 13412 13320
rect 14372 13268 14424 13320
rect 15752 13268 15804 13320
rect 16304 13268 16356 13320
rect 16488 13268 16540 13320
rect 13820 13200 13872 13252
rect 15660 13200 15712 13252
rect 12532 13132 12584 13184
rect 12716 13132 12768 13184
rect 16120 13132 16172 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1860 12971 1912 12980
rect 1860 12937 1869 12971
rect 1869 12937 1903 12971
rect 1903 12937 1912 12971
rect 1860 12928 1912 12937
rect 3516 12928 3568 12980
rect 5172 12928 5224 12980
rect 7748 12928 7800 12980
rect 8024 12928 8076 12980
rect 14096 12928 14148 12980
rect 15660 12928 15712 12980
rect 16120 12928 16172 12980
rect 17868 12928 17920 12980
rect 19432 12971 19484 12980
rect 1584 12792 1636 12844
rect 4160 12835 4212 12844
rect 4160 12801 4169 12835
rect 4169 12801 4203 12835
rect 4203 12801 4212 12835
rect 4160 12792 4212 12801
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 6552 12792 6604 12844
rect 7564 12835 7616 12844
rect 2780 12724 2832 12776
rect 6000 12724 6052 12776
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 14372 12860 14424 12912
rect 15844 12860 15896 12912
rect 16396 12860 16448 12912
rect 17960 12860 18012 12912
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 19984 12971 20036 12980
rect 19984 12937 19993 12971
rect 19993 12937 20027 12971
rect 20027 12937 20036 12971
rect 19984 12928 20036 12937
rect 7840 12724 7892 12776
rect 3148 12656 3200 12708
rect 5172 12656 5224 12708
rect 8392 12792 8444 12844
rect 8668 12792 8720 12844
rect 9588 12792 9640 12844
rect 13452 12792 13504 12844
rect 13636 12835 13688 12844
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 16028 12835 16080 12844
rect 16028 12801 16037 12835
rect 16037 12801 16071 12835
rect 16071 12801 16080 12835
rect 16028 12792 16080 12801
rect 16580 12792 16632 12844
rect 17500 12835 17552 12844
rect 17500 12801 17509 12835
rect 17509 12801 17543 12835
rect 17543 12801 17552 12835
rect 17500 12792 17552 12801
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 4620 12631 4672 12640
rect 4620 12597 4629 12631
rect 4629 12597 4663 12631
rect 4663 12597 4672 12631
rect 4620 12588 4672 12597
rect 5540 12588 5592 12640
rect 10232 12656 10284 12708
rect 10416 12656 10468 12708
rect 14188 12724 14240 12776
rect 15476 12724 15528 12776
rect 16304 12724 16356 12776
rect 20352 12792 20404 12844
rect 12624 12656 12676 12708
rect 13084 12656 13136 12708
rect 13728 12656 13780 12708
rect 16948 12656 17000 12708
rect 18420 12656 18472 12708
rect 20904 12656 20956 12708
rect 9680 12588 9732 12640
rect 11152 12588 11204 12640
rect 13360 12631 13412 12640
rect 13360 12597 13369 12631
rect 13369 12597 13403 12631
rect 13403 12597 13412 12631
rect 13360 12588 13412 12597
rect 19248 12588 19300 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2780 12384 2832 12436
rect 4252 12427 4304 12436
rect 4252 12393 4261 12427
rect 4261 12393 4295 12427
rect 4295 12393 4304 12427
rect 4252 12384 4304 12393
rect 4712 12384 4764 12436
rect 4988 12384 5040 12436
rect 5264 12384 5316 12436
rect 7380 12384 7432 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 9956 12384 10008 12436
rect 13084 12384 13136 12436
rect 13452 12384 13504 12436
rect 16212 12384 16264 12436
rect 17500 12384 17552 12436
rect 17776 12384 17828 12436
rect 2688 12316 2740 12368
rect 4068 12316 4120 12368
rect 15384 12316 15436 12368
rect 17040 12316 17092 12368
rect 17224 12316 17276 12368
rect 17868 12316 17920 12368
rect 18512 12316 18564 12368
rect 19616 12384 19668 12436
rect 20720 12384 20772 12436
rect 20904 12427 20956 12436
rect 20904 12393 20913 12427
rect 20913 12393 20947 12427
rect 20947 12393 20956 12427
rect 20904 12384 20956 12393
rect 1584 12248 1636 12300
rect 4620 12248 4672 12300
rect 5724 12248 5776 12300
rect 7012 12248 7064 12300
rect 4804 12223 4856 12232
rect 4804 12189 4813 12223
rect 4813 12189 4847 12223
rect 4847 12189 4856 12223
rect 4804 12180 4856 12189
rect 4160 12112 4212 12164
rect 8668 12155 8720 12164
rect 8668 12121 8677 12155
rect 8677 12121 8711 12155
rect 8711 12121 8720 12155
rect 8668 12112 8720 12121
rect 10784 12248 10836 12300
rect 13912 12248 13964 12300
rect 14096 12248 14148 12300
rect 17132 12248 17184 12300
rect 17960 12248 18012 12300
rect 9956 12180 10008 12232
rect 10508 12180 10560 12232
rect 11888 12180 11940 12232
rect 14188 12180 14240 12232
rect 4068 12044 4120 12096
rect 12440 12044 12492 12096
rect 14648 12112 14700 12164
rect 15752 12180 15804 12232
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 18604 12223 18656 12232
rect 18604 12189 18613 12223
rect 18613 12189 18647 12223
rect 18647 12189 18656 12223
rect 18604 12180 18656 12189
rect 20168 12180 20220 12232
rect 20444 12223 20496 12232
rect 20444 12189 20453 12223
rect 20453 12189 20487 12223
rect 20487 12189 20496 12223
rect 20444 12180 20496 12189
rect 13912 12044 13964 12096
rect 14004 12044 14056 12096
rect 14372 12044 14424 12096
rect 19524 12044 19576 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 1492 11840 1544 11892
rect 5724 11883 5776 11892
rect 5724 11849 5733 11883
rect 5733 11849 5767 11883
rect 5767 11849 5776 11883
rect 5724 11840 5776 11849
rect 7196 11840 7248 11892
rect 3332 11772 3384 11824
rect 4160 11772 4212 11824
rect 4252 11704 4304 11756
rect 7656 11772 7708 11824
rect 11888 11840 11940 11892
rect 12440 11840 12492 11892
rect 10876 11772 10928 11824
rect 13636 11840 13688 11892
rect 14096 11883 14148 11892
rect 14096 11849 14105 11883
rect 14105 11849 14139 11883
rect 14139 11849 14148 11883
rect 14096 11840 14148 11849
rect 7472 11704 7524 11756
rect 9956 11704 10008 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 17040 11840 17092 11892
rect 17132 11840 17184 11892
rect 19156 11883 19208 11892
rect 19156 11849 19165 11883
rect 19165 11849 19199 11883
rect 19199 11849 19208 11883
rect 19156 11840 19208 11849
rect 19708 11840 19760 11892
rect 19984 11772 20036 11824
rect 14648 11747 14700 11756
rect 14648 11713 14657 11747
rect 14657 11713 14691 11747
rect 14691 11713 14700 11747
rect 15660 11747 15712 11756
rect 14648 11704 14700 11713
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 16028 11704 16080 11756
rect 16764 11704 16816 11756
rect 18236 11704 18288 11756
rect 18604 11704 18656 11756
rect 19708 11747 19760 11756
rect 19708 11713 19717 11747
rect 19717 11713 19751 11747
rect 19751 11713 19760 11747
rect 19708 11704 19760 11713
rect 20444 11704 20496 11756
rect 2504 11636 2556 11688
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 2964 11500 3016 11552
rect 3700 11543 3752 11552
rect 3700 11509 3709 11543
rect 3709 11509 3743 11543
rect 3743 11509 3752 11543
rect 3700 11500 3752 11509
rect 4068 11500 4120 11552
rect 8208 11679 8260 11688
rect 4344 11568 4396 11620
rect 4804 11568 4856 11620
rect 5080 11568 5132 11620
rect 6736 11568 6788 11620
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 8760 11636 8812 11688
rect 10048 11636 10100 11688
rect 11796 11636 11848 11688
rect 12256 11636 12308 11688
rect 12348 11636 12400 11688
rect 15016 11636 15068 11688
rect 15200 11636 15252 11688
rect 19340 11636 19392 11688
rect 19524 11679 19576 11688
rect 19524 11645 19533 11679
rect 19533 11645 19567 11679
rect 19567 11645 19576 11679
rect 19524 11636 19576 11645
rect 11152 11568 11204 11620
rect 8668 11500 8720 11552
rect 9312 11500 9364 11552
rect 11520 11568 11572 11620
rect 11796 11543 11848 11552
rect 11796 11509 11805 11543
rect 11805 11509 11839 11543
rect 11839 11509 11848 11543
rect 11796 11500 11848 11509
rect 14188 11568 14240 11620
rect 12348 11500 12400 11552
rect 12624 11500 12676 11552
rect 14648 11568 14700 11620
rect 16948 11568 17000 11620
rect 17868 11568 17920 11620
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 16304 11500 16356 11552
rect 16488 11543 16540 11552
rect 16488 11509 16497 11543
rect 16497 11509 16531 11543
rect 16531 11509 16540 11543
rect 16488 11500 16540 11509
rect 18696 11500 18748 11552
rect 19524 11500 19576 11552
rect 19892 11500 19944 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2596 11296 2648 11348
rect 2964 11339 3016 11348
rect 2964 11305 2973 11339
rect 2973 11305 3007 11339
rect 3007 11305 3016 11339
rect 2964 11296 3016 11305
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 5632 11296 5684 11348
rect 10232 11296 10284 11348
rect 10600 11296 10652 11348
rect 10876 11296 10928 11348
rect 11796 11296 11848 11348
rect 2044 11228 2096 11280
rect 2412 11271 2464 11280
rect 2412 11237 2421 11271
rect 2421 11237 2455 11271
rect 2455 11237 2464 11271
rect 2412 11228 2464 11237
rect 16396 11296 16448 11348
rect 17132 11339 17184 11348
rect 17132 11305 17141 11339
rect 17141 11305 17175 11339
rect 17175 11305 17184 11339
rect 17132 11296 17184 11305
rect 18696 11339 18748 11348
rect 12348 11228 12400 11280
rect 12532 11228 12584 11280
rect 13636 11228 13688 11280
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 19156 11339 19208 11348
rect 19156 11305 19165 11339
rect 19165 11305 19199 11339
rect 19199 11305 19208 11339
rect 19156 11296 19208 11305
rect 19248 11296 19300 11348
rect 19984 11296 20036 11348
rect 4252 11160 4304 11212
rect 4712 11160 4764 11212
rect 5448 11203 5500 11212
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 6552 11203 6604 11212
rect 6552 11169 6561 11203
rect 6561 11169 6595 11203
rect 6595 11169 6604 11203
rect 6552 11160 6604 11169
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 8484 11160 8536 11212
rect 10048 11160 10100 11212
rect 10140 11203 10192 11212
rect 10140 11169 10149 11203
rect 10149 11169 10183 11203
rect 10183 11169 10192 11203
rect 10140 11160 10192 11169
rect 10324 11160 10376 11212
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 4344 11092 4396 11144
rect 4988 11092 5040 11144
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 7472 11092 7524 11144
rect 6828 11024 6880 11076
rect 7656 11024 7708 11076
rect 6276 10956 6328 11008
rect 9312 11092 9364 11144
rect 10048 11024 10100 11076
rect 10692 11160 10744 11212
rect 12624 11160 12676 11212
rect 13912 11160 13964 11212
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 12440 11092 12492 11144
rect 15844 11160 15896 11212
rect 16028 11203 16080 11212
rect 16028 11169 16062 11203
rect 16062 11169 16080 11203
rect 16028 11160 16080 11169
rect 14096 11067 14148 11076
rect 10140 10956 10192 11008
rect 10508 10956 10560 11008
rect 14096 11033 14105 11067
rect 14105 11033 14139 11067
rect 14139 11033 14148 11067
rect 14096 11024 14148 11033
rect 18604 11160 18656 11212
rect 18696 11160 18748 11212
rect 19616 11160 19668 11212
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 19248 11135 19300 11144
rect 19248 11101 19257 11135
rect 19257 11101 19291 11135
rect 19291 11101 19300 11135
rect 19248 11092 19300 11101
rect 19708 11092 19760 11144
rect 12440 10956 12492 11008
rect 19064 11024 19116 11076
rect 17316 10956 17368 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 2688 10752 2740 10804
rect 3332 10752 3384 10804
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 6552 10752 6604 10804
rect 7564 10795 7616 10804
rect 7564 10761 7573 10795
rect 7573 10761 7607 10795
rect 7607 10761 7616 10795
rect 7564 10752 7616 10761
rect 12624 10795 12676 10804
rect 7012 10727 7064 10736
rect 1584 10548 1636 10600
rect 2504 10548 2556 10600
rect 3332 10480 3384 10532
rect 4988 10548 5040 10600
rect 7012 10693 7021 10727
rect 7021 10693 7055 10727
rect 7055 10693 7064 10727
rect 7012 10684 7064 10693
rect 6276 10659 6328 10668
rect 6276 10625 6285 10659
rect 6285 10625 6319 10659
rect 6319 10625 6328 10659
rect 6276 10616 6328 10625
rect 8484 10684 8536 10736
rect 9588 10684 9640 10736
rect 8300 10616 8352 10668
rect 9312 10616 9364 10668
rect 6368 10548 6420 10600
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 8484 10548 8536 10600
rect 9956 10548 10008 10600
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 12624 10761 12633 10795
rect 12633 10761 12667 10795
rect 12667 10761 12676 10795
rect 12624 10752 12676 10761
rect 13360 10752 13412 10804
rect 16028 10795 16080 10804
rect 16028 10761 16037 10795
rect 16037 10761 16071 10795
rect 16071 10761 16080 10795
rect 16028 10752 16080 10761
rect 16488 10752 16540 10804
rect 18604 10795 18656 10804
rect 18604 10761 18613 10795
rect 18613 10761 18647 10795
rect 18647 10761 18656 10795
rect 18604 10752 18656 10761
rect 19340 10752 19392 10804
rect 19708 10752 19760 10804
rect 20260 10752 20312 10804
rect 11704 10684 11756 10736
rect 12440 10684 12492 10736
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 14188 10659 14240 10668
rect 14188 10625 14197 10659
rect 14197 10625 14231 10659
rect 14231 10625 14240 10659
rect 14188 10616 14240 10625
rect 13176 10548 13228 10600
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 14556 10548 14608 10600
rect 3608 10480 3660 10532
rect 4068 10480 4120 10532
rect 10600 10480 10652 10532
rect 11152 10480 11204 10532
rect 7104 10412 7156 10464
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 9864 10412 9916 10464
rect 15016 10480 15068 10532
rect 17960 10616 18012 10668
rect 18604 10616 18656 10668
rect 19156 10659 19208 10668
rect 17040 10548 17092 10600
rect 18696 10548 18748 10600
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 19248 10548 19300 10600
rect 19616 10548 19668 10600
rect 20628 10591 20680 10600
rect 20628 10557 20637 10591
rect 20637 10557 20671 10591
rect 20671 10557 20680 10591
rect 20628 10548 20680 10557
rect 17500 10480 17552 10532
rect 11888 10455 11940 10464
rect 11888 10421 11897 10455
rect 11897 10421 11931 10455
rect 11931 10421 11940 10455
rect 11888 10412 11940 10421
rect 12348 10412 12400 10464
rect 14004 10412 14056 10464
rect 15108 10412 15160 10464
rect 19524 10480 19576 10532
rect 20168 10480 20220 10532
rect 20260 10480 20312 10532
rect 20996 10480 21048 10532
rect 18696 10412 18748 10464
rect 19340 10412 19392 10464
rect 20352 10412 20404 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 2136 10208 2188 10260
rect 3700 10208 3752 10260
rect 5448 10208 5500 10260
rect 6000 10208 6052 10260
rect 6184 10208 6236 10260
rect 6736 10208 6788 10260
rect 7472 10208 7524 10260
rect 9496 10208 9548 10260
rect 10140 10251 10192 10260
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 2780 10140 2832 10192
rect 4068 10140 4120 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 2872 9936 2924 9988
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 3700 10004 3752 10056
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 4160 9936 4212 9988
rect 6276 10072 6328 10124
rect 7012 10072 7064 10124
rect 8300 10140 8352 10192
rect 9956 10140 10008 10192
rect 11888 10140 11940 10192
rect 11704 10072 11756 10124
rect 12072 10208 12124 10260
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 17776 10208 17828 10260
rect 18512 10208 18564 10260
rect 19064 10208 19116 10260
rect 13728 10183 13780 10192
rect 13728 10149 13737 10183
rect 13737 10149 13771 10183
rect 13771 10149 13780 10183
rect 13728 10140 13780 10149
rect 15752 10140 15804 10192
rect 16580 10140 16632 10192
rect 16856 10140 16908 10192
rect 17316 10140 17368 10192
rect 7932 10047 7984 10056
rect 5172 9868 5224 9920
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 9404 10004 9456 10056
rect 10508 10004 10560 10056
rect 10876 10047 10928 10056
rect 10876 10013 10885 10047
rect 10885 10013 10919 10047
rect 10919 10013 10928 10047
rect 10876 10004 10928 10013
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 13268 10004 13320 10056
rect 14096 10004 14148 10056
rect 14556 10004 14608 10056
rect 15200 10004 15252 10056
rect 15844 10004 15896 10056
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 9588 9936 9640 9988
rect 7840 9868 7892 9920
rect 11888 9868 11940 9920
rect 12256 9911 12308 9920
rect 12256 9877 12265 9911
rect 12265 9877 12299 9911
rect 12299 9877 12308 9911
rect 12256 9868 12308 9877
rect 12440 9868 12492 9920
rect 13360 9911 13412 9920
rect 13360 9877 13369 9911
rect 13369 9877 13403 9911
rect 13403 9877 13412 9911
rect 13360 9868 13412 9877
rect 14004 9936 14056 9988
rect 14648 9936 14700 9988
rect 17960 9936 18012 9988
rect 18236 10072 18288 10124
rect 18144 10004 18196 10056
rect 19156 10140 19208 10192
rect 19800 10140 19852 10192
rect 19064 10072 19116 10124
rect 19340 10072 19392 10124
rect 19984 10072 20036 10124
rect 19708 10004 19760 10056
rect 19156 9936 19208 9988
rect 18788 9868 18840 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 2964 9664 3016 9716
rect 1768 9639 1820 9648
rect 1768 9605 1777 9639
rect 1777 9605 1811 9639
rect 1811 9605 1820 9639
rect 1768 9596 1820 9605
rect 2504 9528 2556 9580
rect 1492 9460 1544 9512
rect 7104 9664 7156 9716
rect 4712 9596 4764 9648
rect 4804 9596 4856 9648
rect 5448 9596 5500 9648
rect 5632 9639 5684 9648
rect 5632 9605 5641 9639
rect 5641 9605 5675 9639
rect 5675 9605 5684 9639
rect 5632 9596 5684 9605
rect 6276 9571 6328 9580
rect 6276 9537 6285 9571
rect 6285 9537 6319 9571
rect 6319 9537 6328 9571
rect 6276 9528 6328 9537
rect 1584 9392 1636 9444
rect 2872 9392 2924 9444
rect 4712 9392 4764 9444
rect 4804 9392 4856 9444
rect 5172 9324 5224 9376
rect 5540 9460 5592 9512
rect 6000 9460 6052 9512
rect 7840 9664 7892 9716
rect 8300 9664 8352 9716
rect 9404 9664 9456 9716
rect 7932 9460 7984 9512
rect 5448 9392 5500 9444
rect 7104 9324 7156 9376
rect 7380 9367 7432 9376
rect 7380 9333 7389 9367
rect 7389 9333 7423 9367
rect 7423 9333 7432 9367
rect 7380 9324 7432 9333
rect 9312 9460 9364 9512
rect 8208 9324 8260 9376
rect 12164 9664 12216 9716
rect 10876 9596 10928 9648
rect 12532 9596 12584 9648
rect 16396 9664 16448 9716
rect 18512 9664 18564 9716
rect 20536 9664 20588 9716
rect 21088 9664 21140 9716
rect 16580 9639 16632 9648
rect 9496 9528 9548 9580
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 12348 9528 12400 9580
rect 16580 9605 16589 9639
rect 16589 9605 16623 9639
rect 16623 9605 16632 9639
rect 16580 9596 16632 9605
rect 14648 9528 14700 9580
rect 10232 9503 10284 9512
rect 10232 9469 10241 9503
rect 10241 9469 10275 9503
rect 10275 9469 10284 9503
rect 10232 9460 10284 9469
rect 9496 9392 9548 9444
rect 11888 9392 11940 9444
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 12716 9460 12768 9512
rect 13360 9460 13412 9512
rect 15200 9503 15252 9512
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 16212 9528 16264 9580
rect 17040 9528 17092 9580
rect 20628 9596 20680 9648
rect 16396 9460 16448 9512
rect 16856 9460 16908 9512
rect 19248 9460 19300 9512
rect 19616 9460 19668 9512
rect 13820 9435 13872 9444
rect 13820 9401 13854 9435
rect 13854 9401 13872 9435
rect 13820 9392 13872 9401
rect 13912 9324 13964 9376
rect 15016 9392 15068 9444
rect 15844 9392 15896 9444
rect 16028 9392 16080 9444
rect 20076 9392 20128 9444
rect 20536 9392 20588 9444
rect 20628 9392 20680 9444
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 17224 9367 17276 9376
rect 16856 9324 16908 9333
rect 17224 9333 17233 9367
rect 17233 9333 17267 9367
rect 17267 9333 17276 9367
rect 17224 9324 17276 9333
rect 19524 9324 19576 9376
rect 19892 9367 19944 9376
rect 19892 9333 19901 9367
rect 19901 9333 19935 9367
rect 19935 9333 19944 9367
rect 19892 9324 19944 9333
rect 20168 9324 20220 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 1124 9120 1176 9172
rect 3608 9120 3660 9172
rect 4252 9163 4304 9172
rect 4252 9129 4261 9163
rect 4261 9129 4295 9163
rect 4295 9129 4304 9163
rect 4252 9120 4304 9129
rect 4988 9120 5040 9172
rect 5724 9120 5776 9172
rect 6092 9120 6144 9172
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 9864 9120 9916 9172
rect 1400 9052 1452 9104
rect 3148 9052 3200 9104
rect 1860 8984 1912 9036
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3608 8916 3660 8968
rect 5264 9052 5316 9104
rect 5448 9052 5500 9104
rect 7380 9052 7432 9104
rect 8576 9052 8628 9104
rect 9496 9052 9548 9104
rect 11796 9052 11848 9104
rect 12256 9052 12308 9104
rect 5080 8984 5132 9036
rect 6736 8984 6788 9036
rect 5540 8916 5592 8968
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 6920 8916 6972 8968
rect 4068 8848 4120 8900
rect 8300 8984 8352 9036
rect 10876 8984 10928 9036
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 12348 9027 12400 9036
rect 12348 8993 12382 9027
rect 12382 8993 12400 9027
rect 12348 8984 12400 8993
rect 12532 9120 12584 9172
rect 13728 9120 13780 9172
rect 16028 9120 16080 9172
rect 16764 9163 16816 9172
rect 16764 9129 16773 9163
rect 16773 9129 16807 9163
rect 16807 9129 16816 9163
rect 16764 9120 16816 9129
rect 16856 9120 16908 9172
rect 17224 9120 17276 9172
rect 20076 9120 20128 9172
rect 20352 9120 20404 9172
rect 12716 9052 12768 9104
rect 19616 9052 19668 9104
rect 14464 8984 14516 9036
rect 15292 8984 15344 9036
rect 8024 8959 8076 8968
rect 8024 8925 8033 8959
rect 8033 8925 8067 8959
rect 8067 8925 8076 8959
rect 8024 8916 8076 8925
rect 8208 8916 8260 8968
rect 14096 8916 14148 8968
rect 15016 8916 15068 8968
rect 5540 8780 5592 8832
rect 9956 8848 10008 8900
rect 13452 8891 13504 8900
rect 11612 8780 11664 8832
rect 13452 8857 13461 8891
rect 13461 8857 13495 8891
rect 13495 8857 13504 8891
rect 13452 8848 13504 8857
rect 13820 8848 13872 8900
rect 14280 8848 14332 8900
rect 15752 9027 15804 9036
rect 15752 8993 15761 9027
rect 15761 8993 15795 9027
rect 15795 8993 15804 9027
rect 15752 8984 15804 8993
rect 19340 8984 19392 9036
rect 15660 8848 15712 8900
rect 17868 8916 17920 8968
rect 17500 8848 17552 8900
rect 14188 8780 14240 8832
rect 15752 8780 15804 8832
rect 16304 8823 16356 8832
rect 16304 8789 16313 8823
rect 16313 8789 16347 8823
rect 16347 8789 16356 8823
rect 16304 8780 16356 8789
rect 16396 8780 16448 8832
rect 19800 8780 19852 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2872 8576 2924 8628
rect 4160 8576 4212 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 6000 8576 6052 8628
rect 12440 8576 12492 8628
rect 12624 8576 12676 8628
rect 14096 8619 14148 8628
rect 4344 8508 4396 8560
rect 2688 8440 2740 8492
rect 3976 8440 4028 8492
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 5632 8440 5684 8492
rect 1584 8372 1636 8424
rect 4436 8372 4488 8424
rect 5448 8372 5500 8424
rect 2320 8304 2372 8356
rect 2504 8304 2556 8356
rect 3700 8304 3752 8356
rect 4160 8304 4212 8356
rect 4344 8304 4396 8356
rect 8024 8508 8076 8560
rect 8576 8508 8628 8560
rect 2780 8236 2832 8288
rect 3792 8236 3844 8288
rect 4620 8236 4672 8288
rect 4712 8236 4764 8288
rect 5724 8236 5776 8288
rect 8208 8372 8260 8424
rect 9956 8440 10008 8492
rect 11060 8508 11112 8560
rect 14096 8585 14105 8619
rect 14105 8585 14139 8619
rect 14139 8585 14148 8619
rect 14096 8576 14148 8585
rect 14188 8576 14240 8628
rect 15476 8576 15528 8628
rect 15568 8576 15620 8628
rect 16672 8576 16724 8628
rect 17408 8576 17460 8628
rect 17500 8576 17552 8628
rect 11612 8440 11664 8492
rect 13452 8440 13504 8492
rect 15660 8440 15712 8492
rect 18052 8508 18104 8560
rect 19340 8576 19392 8628
rect 20076 8508 20128 8560
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 20628 8440 20680 8492
rect 11704 8415 11756 8424
rect 7196 8304 7248 8356
rect 7564 8304 7616 8356
rect 8116 8304 8168 8356
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 12072 8372 12124 8424
rect 16948 8415 17000 8424
rect 10968 8304 11020 8356
rect 11152 8304 11204 8356
rect 12256 8304 12308 8356
rect 12716 8347 12768 8356
rect 12716 8313 12750 8347
rect 12750 8313 12768 8347
rect 12716 8304 12768 8313
rect 7012 8279 7064 8288
rect 7012 8245 7021 8279
rect 7021 8245 7055 8279
rect 7055 8245 7064 8279
rect 7012 8236 7064 8245
rect 7104 8236 7156 8288
rect 8852 8236 8904 8288
rect 9956 8279 10008 8288
rect 9956 8245 9965 8279
rect 9965 8245 9999 8279
rect 9999 8245 10008 8279
rect 9956 8236 10008 8245
rect 10232 8279 10284 8288
rect 10232 8245 10241 8279
rect 10241 8245 10275 8279
rect 10275 8245 10284 8279
rect 10232 8236 10284 8245
rect 10324 8236 10376 8288
rect 13268 8236 13320 8288
rect 13912 8236 13964 8288
rect 16948 8381 16957 8415
rect 16957 8381 16991 8415
rect 16991 8381 17000 8415
rect 16948 8372 17000 8381
rect 17132 8372 17184 8424
rect 17868 8372 17920 8424
rect 19984 8372 20036 8424
rect 18604 8304 18656 8356
rect 19156 8304 19208 8356
rect 15016 8236 15068 8288
rect 15292 8279 15344 8288
rect 15292 8245 15301 8279
rect 15301 8245 15335 8279
rect 15335 8245 15344 8279
rect 15292 8236 15344 8245
rect 15568 8236 15620 8288
rect 16396 8236 16448 8288
rect 19616 8236 19668 8288
rect 20352 8304 20404 8356
rect 20720 8236 20772 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 1860 8032 1912 8084
rect 3884 8032 3936 8084
rect 4436 8032 4488 8084
rect 2780 7896 2832 7948
rect 2872 7896 2924 7948
rect 3608 7964 3660 8016
rect 6000 7964 6052 8016
rect 7012 8032 7064 8084
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 9128 8032 9180 8084
rect 9588 8032 9640 8084
rect 10232 8032 10284 8084
rect 15016 8032 15068 8084
rect 16304 8032 16356 8084
rect 18052 8032 18104 8084
rect 20352 8032 20404 8084
rect 4160 7896 4212 7948
rect 4804 7896 4856 7948
rect 5724 7896 5776 7948
rect 6276 7896 6328 7948
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 3332 7828 3384 7880
rect 4344 7828 4396 7880
rect 4712 7828 4764 7880
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 9956 7964 10008 8016
rect 10324 7964 10376 8016
rect 12532 7964 12584 8016
rect 15384 7964 15436 8016
rect 15752 8007 15804 8016
rect 15752 7973 15761 8007
rect 15761 7973 15795 8007
rect 15795 7973 15804 8007
rect 15752 7964 15804 7973
rect 17224 7964 17276 8016
rect 20260 8007 20312 8016
rect 20260 7973 20269 8007
rect 20269 7973 20303 8007
rect 20303 7973 20312 8007
rect 20260 7964 20312 7973
rect 8852 7871 8904 7880
rect 8852 7837 8861 7871
rect 8861 7837 8895 7871
rect 8895 7837 8904 7871
rect 8852 7828 8904 7837
rect 9956 7828 10008 7880
rect 10968 7896 11020 7948
rect 11980 7896 12032 7948
rect 12992 7939 13044 7948
rect 12992 7905 13001 7939
rect 13001 7905 13035 7939
rect 13035 7905 13044 7939
rect 12992 7896 13044 7905
rect 18972 7896 19024 7948
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 4068 7760 4120 7812
rect 5448 7692 5500 7744
rect 6920 7760 6972 7812
rect 7196 7760 7248 7812
rect 8208 7760 8260 7812
rect 11704 7828 11756 7880
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 17040 7871 17092 7880
rect 17040 7837 17049 7871
rect 17049 7837 17083 7871
rect 17083 7837 17092 7871
rect 17040 7828 17092 7837
rect 12348 7760 12400 7812
rect 16856 7760 16908 7812
rect 18604 7760 18656 7812
rect 20628 7828 20680 7880
rect 12532 7692 12584 7744
rect 13912 7692 13964 7744
rect 15936 7692 15988 7744
rect 17960 7692 18012 7744
rect 19708 7692 19760 7744
rect 20628 7692 20680 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 1584 7284 1636 7336
rect 3332 7284 3384 7336
rect 3976 7463 4028 7472
rect 3976 7429 3985 7463
rect 3985 7429 4019 7463
rect 4019 7429 4028 7463
rect 3976 7420 4028 7429
rect 2320 7148 2372 7200
rect 5632 7488 5684 7540
rect 4252 7284 4304 7336
rect 17684 7488 17736 7540
rect 18972 7488 19024 7540
rect 19248 7531 19300 7540
rect 19248 7497 19257 7531
rect 19257 7497 19291 7531
rect 19291 7497 19300 7531
rect 19248 7488 19300 7497
rect 19524 7488 19576 7540
rect 4068 7216 4120 7268
rect 5264 7259 5316 7268
rect 5264 7225 5298 7259
rect 5298 7225 5316 7259
rect 5264 7216 5316 7225
rect 6920 7284 6972 7336
rect 8576 7284 8628 7336
rect 12992 7420 13044 7472
rect 19064 7420 19116 7472
rect 19340 7420 19392 7472
rect 17224 7352 17276 7404
rect 19708 7395 19760 7404
rect 19708 7361 19717 7395
rect 19717 7361 19751 7395
rect 19751 7361 19760 7395
rect 19708 7352 19760 7361
rect 19892 7352 19944 7404
rect 18512 7284 18564 7336
rect 18972 7284 19024 7336
rect 19616 7327 19668 7336
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 20628 7327 20680 7336
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 20628 7284 20680 7293
rect 7564 7216 7616 7268
rect 5540 7148 5592 7200
rect 5724 7148 5776 7200
rect 8852 7216 8904 7268
rect 18696 7148 18748 7200
rect 18880 7148 18932 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 2780 6987 2832 6996
rect 2780 6953 2789 6987
rect 2789 6953 2823 6987
rect 2823 6953 2832 6987
rect 2780 6944 2832 6953
rect 17224 6944 17276 6996
rect 5264 6876 5316 6928
rect 3148 6851 3200 6860
rect 3148 6817 3157 6851
rect 3157 6817 3191 6851
rect 3191 6817 3200 6851
rect 3148 6808 3200 6817
rect 3884 6808 3936 6860
rect 4988 6808 5040 6860
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 5172 6740 5224 6792
rect 6000 6851 6052 6860
rect 6000 6817 6009 6851
rect 6009 6817 6043 6851
rect 6043 6817 6052 6851
rect 6000 6808 6052 6817
rect 17040 6876 17092 6928
rect 4804 6672 4856 6724
rect 14280 6672 14332 6724
rect 5540 6604 5592 6656
rect 8944 6604 8996 6656
rect 17960 6604 18012 6656
rect 19432 6808 19484 6860
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 20076 6604 20128 6656
rect 20352 6604 20404 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 3056 6400 3108 6452
rect 5080 6443 5132 6452
rect 5080 6409 5089 6443
rect 5089 6409 5123 6443
rect 5123 6409 5132 6443
rect 5080 6400 5132 6409
rect 12256 6400 12308 6452
rect 18512 6400 18564 6452
rect 20076 6400 20128 6452
rect 20444 6443 20496 6452
rect 20444 6409 20453 6443
rect 20453 6409 20487 6443
rect 20487 6409 20496 6443
rect 20444 6400 20496 6409
rect 4068 6332 4120 6384
rect 12164 6332 12216 6384
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 3148 6264 3200 6316
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 13636 6264 13688 6316
rect 18788 6264 18840 6316
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 2228 6128 2280 6180
rect 19800 6196 19852 6248
rect 20076 6196 20128 6248
rect 20352 6128 20404 6180
rect 19708 6060 19760 6112
rect 20536 6060 20588 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 4068 5584 4120 5636
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 19800 5559 19852 5568
rect 19800 5525 19809 5559
rect 19809 5525 19843 5559
rect 19843 5525 19852 5559
rect 19800 5516 19852 5525
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 5908 5312 5960 5364
rect 17960 5312 18012 5364
rect 19708 5312 19760 5364
rect 3976 5244 4028 5296
rect 5356 5244 5408 5296
rect 19800 5176 19852 5228
rect 20444 5219 20496 5228
rect 20444 5185 20453 5219
rect 20453 5185 20487 5219
rect 20487 5185 20496 5219
rect 20444 5176 20496 5185
rect 20536 5108 20588 5160
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 6736 4088 6788 4140
rect 7472 4088 7524 4140
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 20444 3000 20496 3052
rect 11152 2932 11204 2984
rect 15844 2932 15896 2984
rect 6092 2864 6144 2916
rect 9772 2864 9824 2916
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 2964 1164 3016 1216
rect 6276 1164 6328 1216
<< metal2 >>
rect 202 22000 258 22800
rect 570 22000 626 22800
rect 1030 22000 1086 22800
rect 1398 22000 1454 22800
rect 1858 22000 1914 22800
rect 2226 22000 2282 22800
rect 2686 22000 2742 22800
rect 3054 22536 3110 22545
rect 3054 22471 3110 22480
rect 2778 22128 2834 22137
rect 2778 22063 2834 22072
rect 216 19310 244 22000
rect 204 19304 256 19310
rect 204 19246 256 19252
rect 584 16726 612 22000
rect 1044 18902 1072 22000
rect 1032 18896 1084 18902
rect 1032 18838 1084 18844
rect 1412 18086 1440 22000
rect 1872 18290 1900 22000
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1964 18970 1992 19751
rect 2042 19272 2098 19281
rect 2042 19207 2098 19216
rect 2056 19174 2084 19207
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 2044 18828 2096 18834
rect 1964 18426 1992 18799
rect 2044 18770 2096 18776
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 572 16720 624 16726
rect 572 16662 624 16668
rect 1688 14618 1716 17682
rect 1780 17542 1808 18158
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 1780 14929 1808 16594
rect 1872 15026 1900 17070
rect 1952 16992 2004 16998
rect 1950 16960 1952 16969
rect 2004 16960 2006 16969
rect 1950 16895 2006 16904
rect 1950 16552 2006 16561
rect 1950 16487 1952 16496
rect 2004 16487 2006 16496
rect 1952 16458 2004 16464
rect 2056 16454 2084 18770
rect 2136 18760 2188 18766
rect 2134 18728 2136 18737
rect 2188 18728 2190 18737
rect 2134 18663 2190 18672
rect 2240 18358 2268 22000
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2608 18873 2636 19654
rect 2700 18902 2728 22000
rect 2792 20058 2820 22063
rect 2962 21584 3018 21593
rect 2962 21519 3018 21528
rect 2870 20632 2926 20641
rect 2870 20567 2926 20576
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2884 19242 2912 20567
rect 2872 19236 2924 19242
rect 2872 19178 2924 19184
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2688 18896 2740 18902
rect 2594 18864 2650 18873
rect 2688 18838 2740 18844
rect 2594 18799 2650 18808
rect 2792 18426 2820 19071
rect 2976 18970 3004 21519
rect 3068 18970 3096 22471
rect 3146 22000 3202 22800
rect 3514 22000 3570 22800
rect 3974 22000 4030 22800
rect 4342 22000 4398 22800
rect 4802 22000 4858 22800
rect 5262 22000 5318 22800
rect 5630 22000 5686 22800
rect 6090 22000 6146 22800
rect 6458 22000 6514 22800
rect 6918 22000 6974 22800
rect 7378 22000 7434 22800
rect 7746 22000 7802 22800
rect 8206 22000 8262 22800
rect 8574 22000 8630 22800
rect 9034 22000 9090 22800
rect 9494 22000 9550 22800
rect 9862 22000 9918 22800
rect 10322 22000 10378 22800
rect 10690 22000 10746 22800
rect 11150 22000 11206 22800
rect 11610 22000 11666 22800
rect 11978 22000 12034 22800
rect 12438 22000 12494 22800
rect 12806 22000 12862 22800
rect 13266 22000 13322 22800
rect 13634 22000 13690 22800
rect 14094 22000 14150 22800
rect 14554 22000 14610 22800
rect 14922 22000 14978 22800
rect 15382 22000 15438 22800
rect 15750 22000 15806 22800
rect 16210 22000 16266 22800
rect 16670 22000 16726 22800
rect 17038 22000 17094 22800
rect 17498 22000 17554 22800
rect 17774 22536 17830 22545
rect 17774 22471 17830 22480
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3160 18630 3188 22000
rect 3528 20346 3556 22000
rect 3528 20318 3648 20346
rect 3514 20224 3570 20233
rect 3514 20159 3570 20168
rect 3528 19514 3556 20159
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 3620 18970 3648 20318
rect 3700 19916 3752 19922
rect 3700 19858 3752 19864
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2228 18352 2280 18358
rect 2228 18294 2280 18300
rect 3146 18320 3202 18329
rect 3146 18255 3202 18264
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2332 17814 2360 18158
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 2136 17672 2188 17678
rect 2134 17640 2136 17649
rect 2188 17640 2190 17649
rect 2134 17575 2190 17584
rect 2778 17368 2834 17377
rect 2778 17303 2780 17312
rect 2832 17303 2834 17312
rect 2780 17274 2832 17280
rect 2884 17270 2912 18022
rect 2872 17264 2924 17270
rect 2872 17206 2924 17212
rect 2412 17060 2464 17066
rect 2412 17002 2464 17008
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1964 15609 1992 15846
rect 1950 15600 2006 15609
rect 1950 15535 2006 15544
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1964 15065 1992 15302
rect 1950 15056 2006 15065
rect 1860 15020 1912 15026
rect 1950 14991 2006 15000
rect 1860 14962 1912 14968
rect 1766 14920 1822 14929
rect 1766 14855 1822 14864
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1688 14074 1716 14418
rect 1858 14104 1914 14113
rect 1676 14068 1728 14074
rect 1858 14039 1914 14048
rect 1676 14010 1728 14016
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1504 11898 1532 13330
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 12306 1624 12786
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1492 11892 1544 11898
rect 1492 11834 1544 11840
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1124 9172 1176 9178
rect 1124 9114 1176 9120
rect 1136 4321 1164 9114
rect 1412 9110 1440 10066
rect 1504 9518 1532 11494
rect 1596 10606 1624 12242
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1596 9450 1624 10542
rect 1780 9654 1808 13670
rect 1872 12986 1900 14039
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 2056 11286 2084 16390
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2332 15366 2360 15982
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 2148 10266 2176 13806
rect 2240 13530 2268 14350
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2332 13190 2360 13874
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2424 11286 2452 17002
rect 2884 16658 2912 17206
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2502 16008 2558 16017
rect 2502 15943 2558 15952
rect 2516 15910 2544 15943
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2870 14648 2926 14657
rect 2870 14583 2926 14592
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2700 13462 2728 13806
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2516 11150 2544 11630
rect 2608 11354 2636 13330
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12374 2728 13126
rect 2792 12782 2820 14350
rect 2884 14074 2912 14583
rect 2976 14464 3004 18158
rect 3054 17912 3110 17921
rect 3054 17847 3110 17856
rect 3068 17338 3096 17847
rect 3160 17338 3188 18255
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3252 16969 3280 18770
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3528 17882 3556 18362
rect 3606 18184 3662 18193
rect 3606 18119 3662 18128
rect 3620 18086 3648 18119
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3344 17542 3372 17682
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3436 17134 3464 17478
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3238 16960 3294 16969
rect 3238 16895 3294 16904
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3068 14958 3096 15982
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2976 14436 3096 14464
rect 2964 14340 3016 14346
rect 2964 14282 3016 14288
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2870 13696 2926 13705
rect 2870 13631 2926 13640
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2792 12442 2820 12718
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2516 10606 2544 11086
rect 2700 10810 2728 12310
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2516 10062 2544 10542
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 2516 9586 2544 9998
rect 2792 9874 2820 10134
rect 2884 9994 2912 13631
rect 2976 13394 3004 14282
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 3068 13297 3096 14436
rect 3160 13462 3188 15914
rect 3252 15706 3280 16730
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3240 14884 3292 14890
rect 3344 14872 3372 16526
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3436 15502 3464 15914
rect 3528 15638 3556 17818
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3620 16046 3648 16526
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3516 15632 3568 15638
rect 3516 15574 3568 15580
rect 3608 15564 3660 15570
rect 3608 15506 3660 15512
rect 3424 15496 3476 15502
rect 3620 15450 3648 15506
rect 3424 15438 3476 15444
rect 3436 15094 3464 15438
rect 3528 15422 3648 15450
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3292 14844 3372 14872
rect 3240 14826 3292 14832
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 3054 13288 3110 13297
rect 3054 13223 3110 13232
rect 3252 13172 3280 14826
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3344 13716 3372 14486
rect 3436 14414 3464 15030
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3528 14278 3556 15422
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 3344 13688 3464 13716
rect 3068 13144 3280 13172
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 11354 3004 11494
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2792 9846 3004 9874
rect 2976 9722 3004 9846
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 1400 9104 1452 9110
rect 1400 9046 1452 9052
rect 1596 8430 1624 9386
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 7342 1624 8366
rect 1872 8090 1900 8978
rect 2884 8974 2912 9386
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2700 8498 2728 8910
rect 2884 8634 2912 8910
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 2332 7886 2360 8298
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 6322 1624 7278
rect 2332 7206 2360 7822
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 1122 4312 1178 4321
rect 1122 4247 1178 4256
rect 2240 800 2268 6122
rect 2226 0 2282 800
rect 2516 649 2544 8298
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 8106 2820 8230
rect 2700 8078 2820 8106
rect 2700 7585 2728 8078
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2686 7576 2742 7585
rect 2686 7511 2742 7520
rect 2792 7002 2820 7890
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2884 2553 2912 7890
rect 2870 2544 2926 2553
rect 2870 2479 2926 2488
rect 2976 1306 3004 9658
rect 3068 6458 3096 13144
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3160 9110 3188 12650
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3344 10810 3372 11766
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3344 10538 3372 10746
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3344 7342 3372 7822
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3160 6322 3188 6802
rect 3344 6798 3372 7278
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3252 3505 3280 6734
rect 3436 5817 3464 13688
rect 3528 12986 3556 13738
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3620 10826 3648 14418
rect 3712 12458 3740 19858
rect 3988 19310 4016 22000
rect 4066 21176 4122 21185
rect 4066 21111 4122 21120
rect 4080 21010 4108 21111
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4356 19700 4384 22000
rect 4172 19672 4384 19700
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3792 18828 3844 18834
rect 3792 18770 3844 18776
rect 3804 12628 3832 18770
rect 3976 18352 4028 18358
rect 3974 18320 3976 18329
rect 4028 18320 4030 18329
rect 3974 18255 4030 18264
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3896 12730 3924 18158
rect 3976 15972 4028 15978
rect 3976 15914 4028 15920
rect 3988 15366 4016 15914
rect 4172 15722 4200 19672
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4816 18154 4844 22000
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4724 16726 4752 17138
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4724 16182 4752 16662
rect 4816 16250 4844 16934
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4172 15694 4844 15722
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4816 15314 4844 15694
rect 4908 15434 4936 16934
rect 5000 15745 5028 19790
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5092 17338 5120 17682
rect 5184 17513 5212 19246
rect 5170 17504 5226 17513
rect 5170 17439 5226 17448
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5276 16250 5304 22000
rect 5354 18728 5410 18737
rect 5354 18663 5356 18672
rect 5408 18663 5410 18672
rect 5356 18634 5408 18640
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5172 16176 5224 16182
rect 5172 16118 5224 16124
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 4986 15736 5042 15745
rect 4986 15671 5042 15680
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 4896 15428 4948 15434
rect 4896 15370 4948 15376
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3988 14482 4016 14894
rect 4172 14618 4200 15302
rect 4816 15286 4936 15314
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4252 14884 4304 14890
rect 4252 14826 4304 14832
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3988 13870 4016 14418
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4172 12850 4200 13330
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 3896 12702 4016 12730
rect 3804 12600 3924 12628
rect 3712 12430 3832 12458
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3528 10798 3648 10826
rect 3528 9908 3556 10798
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3620 10062 3648 10474
rect 3712 10266 3740 11494
rect 3804 11393 3832 12430
rect 3790 11384 3846 11393
rect 3790 11319 3846 11328
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3528 9880 3648 9908
rect 3620 9178 3648 9880
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3620 8022 3648 8910
rect 3712 8362 3740 9998
rect 3896 9160 3924 12600
rect 3988 9489 4016 12702
rect 4264 12442 4292 14826
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4632 14618 4660 14758
rect 4724 14618 4752 14758
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4816 14006 4844 14350
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4068 12368 4120 12374
rect 4066 12336 4068 12345
rect 4120 12336 4122 12345
rect 4632 12306 4660 12582
rect 4724 12442 4752 13126
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4066 12271 4122 12280
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4816 12238 4844 13942
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11801 4108 12038
rect 4172 11830 4200 12106
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4160 11824 4212 11830
rect 4066 11792 4122 11801
rect 4160 11766 4212 11772
rect 4066 11727 4122 11736
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4264 11642 4292 11698
rect 4264 11626 4384 11642
rect 4264 11620 4396 11626
rect 4264 11614 4344 11620
rect 4344 11562 4396 11568
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 11354 4108 11494
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4066 10840 4122 10849
rect 4066 10775 4122 10784
rect 4080 10538 4108 10775
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4080 10198 4108 10367
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 3974 9480 4030 9489
rect 3974 9415 4030 9424
rect 3804 9132 3924 9160
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3804 8294 3832 9132
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4080 8537 4108 8842
rect 4172 8634 4200 9930
rect 4264 9178 4292 11154
rect 4356 11150 4384 11562
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4724 9654 4752 11154
rect 4816 10810 4844 11562
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4816 9450 4844 9590
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4344 8560 4396 8566
rect 4066 8528 4122 8537
rect 3976 8492 4028 8498
rect 4264 8508 4344 8514
rect 4264 8502 4396 8508
rect 4066 8463 4122 8472
rect 4160 8492 4212 8498
rect 3976 8434 4028 8440
rect 4160 8434 4212 8440
rect 4264 8486 4384 8502
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3896 6866 3924 8026
rect 3988 7478 4016 8434
rect 4172 8362 4200 8434
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 4080 7818 4108 8055
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4080 7177 4108 7210
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 4066 6760 4122 6769
rect 4066 6695 4122 6704
rect 4080 6390 4108 6695
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3422 5808 3478 5817
rect 3422 5743 3478 5752
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3976 5296 4028 5302
rect 3974 5264 3976 5273
rect 4028 5264 4030 5273
rect 3974 5199 4030 5208
rect 4080 4865 4108 5578
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 4066 1592 4122 1601
rect 4172 1578 4200 7890
rect 4264 7342 4292 8486
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4618 8392 4674 8401
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4356 7886 4384 8298
rect 4448 8090 4476 8366
rect 4618 8327 4674 8336
rect 4632 8294 4660 8327
rect 4724 8294 4752 9386
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4724 7886 4752 8230
rect 4816 7954 4844 9386
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4724 3913 4752 7822
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4816 6225 4844 6666
rect 4802 6216 4858 6225
rect 4802 6151 4858 6160
rect 4710 3904 4766 3913
rect 4710 3839 4766 3848
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4908 3058 4936 15286
rect 5000 15026 5028 15506
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5000 12442 5028 13330
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5092 11801 5120 15846
rect 5184 15570 5212 16118
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5276 15502 5304 16050
rect 5264 15496 5316 15502
rect 5170 15464 5226 15473
rect 5264 15438 5316 15444
rect 5170 15399 5226 15408
rect 5184 13394 5212 15399
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 5184 12986 5212 13194
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5184 12850 5212 12922
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5078 11792 5134 11801
rect 5078 11727 5134 11736
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5000 10606 5028 11086
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 5092 10146 5120 11562
rect 5000 10118 5120 10146
rect 5000 9178 5028 10118
rect 5080 10056 5132 10062
rect 5184 10044 5212 12650
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5132 10016 5212 10044
rect 5080 9998 5132 10004
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5184 9382 5212 9862
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5000 6866 5028 9114
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 5000 2961 5028 6802
rect 5092 6458 5120 8978
rect 5184 6798 5212 9318
rect 5276 9110 5304 12378
rect 5368 11529 5396 18090
rect 5460 16697 5488 18566
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5446 16688 5502 16697
rect 5446 16623 5502 16632
rect 5460 16046 5488 16623
rect 5552 16590 5580 16730
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5538 16008 5594 16017
rect 5538 15943 5594 15952
rect 5552 15706 5580 15943
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5552 15076 5580 15642
rect 5644 15144 5672 22000
rect 5724 21004 5776 21010
rect 5724 20946 5776 20952
rect 5736 19514 5764 20946
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 6104 19394 6132 22000
rect 6104 19366 6224 19394
rect 6196 19310 6224 19366
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 6184 19304 6236 19310
rect 6184 19246 6236 19252
rect 6104 18290 6132 19246
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6380 18465 6408 19110
rect 6366 18456 6422 18465
rect 6366 18391 6422 18400
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5816 17604 5868 17610
rect 5816 17546 5868 17552
rect 5828 17338 5856 17546
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5736 15586 5764 16186
rect 5828 15706 5856 16934
rect 5920 16590 5948 18022
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6012 16726 6040 17138
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5920 16250 5948 16526
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5736 15558 5856 15586
rect 5644 15116 5764 15144
rect 5552 15048 5672 15076
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5460 14482 5488 14894
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5460 14056 5488 14418
rect 5540 14068 5592 14074
rect 5460 14028 5540 14056
rect 5540 14010 5592 14016
rect 5644 13954 5672 15048
rect 5460 13926 5672 13954
rect 5354 11520 5410 11529
rect 5354 11455 5410 11464
rect 5460 11370 5488 13926
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5552 12646 5580 13330
rect 5736 13190 5764 15116
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5736 11898 5764 12242
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5828 11778 5856 15558
rect 6288 15366 6316 17070
rect 6380 16538 6408 18391
rect 6472 17105 6500 22000
rect 6932 19938 6960 22000
rect 6932 19910 7144 19938
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6564 18290 6592 18702
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6458 17096 6514 17105
rect 6458 17031 6514 17040
rect 6550 16960 6606 16969
rect 6550 16895 6606 16904
rect 6380 16510 6500 16538
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6288 14958 6316 15302
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6366 14920 6422 14929
rect 6366 14855 6422 14864
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 6104 13530 6132 14486
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5368 11342 5488 11370
rect 5736 11750 5856 11778
rect 5906 11792 5962 11801
rect 5632 11348 5684 11354
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5276 7274 5304 7822
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5276 6934 5304 7210
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 4986 2952 5042 2961
rect 4986 2887 5042 2896
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 5184 2009 5212 6734
rect 5368 5302 5396 11342
rect 5632 11290 5684 11296
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10266 5488 11154
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5644 9654 5672 11290
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5460 9450 5488 9590
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5460 8430 5488 9046
rect 5552 8974 5580 9454
rect 5736 9178 5764 11750
rect 5906 11727 5962 11736
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5540 8968 5592 8974
rect 5724 8968 5776 8974
rect 5592 8916 5672 8922
rect 5540 8910 5672 8916
rect 5724 8910 5776 8916
rect 5552 8894 5672 8910
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 6254 5488 7686
rect 5552 7206 5580 8774
rect 5644 8498 5672 8894
rect 5736 8634 5764 8910
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 7954 5764 8230
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5644 7546 5672 7822
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5736 7206 5764 7890
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6322 5580 6598
rect 5736 6322 5764 7142
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5920 5370 5948 11727
rect 6012 10266 6040 12718
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6288 10674 6316 10950
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 5998 9616 6054 9625
rect 5998 9551 6054 9560
rect 6012 9518 6040 9551
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6196 9466 6224 10202
rect 6288 10130 6316 10610
rect 6380 10606 6408 14855
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6288 9586 6316 10066
rect 6472 10033 6500 16510
rect 6564 12850 6592 16895
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6656 15638 6684 15914
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6748 15314 6776 18158
rect 6840 17785 6868 19246
rect 6932 18902 6960 19722
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 6932 18086 6960 18838
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 7024 17882 7052 19246
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6826 17776 6882 17785
rect 6826 17711 6882 17720
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 17202 6960 17478
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6840 16794 6868 16934
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6748 15286 6868 15314
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6656 13326 6684 14962
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 10810 6592 11154
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6656 10146 6684 13126
rect 6748 11626 6776 13262
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10266 6776 11086
rect 6840 11082 6868 15286
rect 6932 14618 6960 15982
rect 7024 15162 7052 17614
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7024 14414 7052 14962
rect 7116 14550 7144 19910
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17134 7236 17478
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7300 16946 7328 19110
rect 7208 16918 7328 16946
rect 7208 16658 7236 16918
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7208 15910 7236 16594
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7300 15978 7328 16390
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15026 7236 15846
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 7024 13870 7052 14350
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6932 13297 6960 13330
rect 6918 13288 6974 13297
rect 6918 13223 6974 13232
rect 7024 12306 7052 13806
rect 7116 13462 7144 14486
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7208 11898 7236 14418
rect 7392 12442 7420 22000
rect 7760 20074 7788 22000
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7668 20046 7788 20074
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7484 17882 7512 19654
rect 7576 19514 7604 19790
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7576 18766 7604 19178
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7576 17202 7604 18566
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7484 16726 7512 17138
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7484 16250 7512 16662
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7484 15484 7512 16186
rect 7564 15496 7616 15502
rect 7484 15456 7564 15484
rect 7564 15438 7616 15444
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7576 13870 7604 14214
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 13462 7604 13806
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6656 10118 6776 10146
rect 7024 10130 7052 10678
rect 7208 10606 7236 11834
rect 7484 11762 7512 13330
rect 7576 12850 7604 13398
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7668 11830 7696 20046
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7760 19446 7788 19858
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 7944 19224 7972 19450
rect 8116 19236 8168 19242
rect 7944 19196 8116 19224
rect 8116 19178 8168 19184
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18630 7788 19110
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8220 18970 8248 22000
rect 8484 19984 8536 19990
rect 8484 19926 8536 19932
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 7760 17678 7788 18566
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17882 8248 18566
rect 8312 18086 8340 18702
rect 8404 18698 8432 18770
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8312 17728 8340 18022
rect 8404 17882 8432 18634
rect 8496 18290 8524 19926
rect 8588 18358 8616 22000
rect 9048 19938 9076 22000
rect 9048 19910 9260 19938
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8680 18426 8708 18702
rect 8864 18601 8892 18770
rect 8850 18592 8906 18601
rect 8850 18527 8906 18536
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8484 17740 8536 17746
rect 8312 17700 8484 17728
rect 8484 17682 8536 17688
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8036 17241 8064 17274
rect 8022 17232 8078 17241
rect 8022 17167 8078 17176
rect 8680 17134 8708 18362
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8312 16658 8340 17002
rect 8680 16998 8708 17070
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8588 16794 8616 16934
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15162 8340 15506
rect 8404 15434 8432 16594
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8496 15910 8524 16050
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8680 14890 8708 15574
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8668 14884 8720 14890
rect 8588 14844 8668 14872
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7760 12986 7788 14758
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8128 14074 8156 14418
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8312 13530 8340 14758
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7852 12782 7880 13330
rect 8036 12986 8064 13398
rect 8404 13326 8432 14010
rect 8392 13320 8444 13326
rect 8114 13288 8170 13297
rect 8392 13262 8444 13268
rect 8114 13223 8116 13232
rect 8168 13223 8170 13232
rect 8116 13194 8168 13200
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8312 12782 8340 13126
rect 8404 12850 8432 13262
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 6458 10024 6514 10033
rect 6458 9959 6514 9968
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6196 9438 6316 9466
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 5998 9072 6054 9081
rect 5998 9007 6054 9016
rect 6012 8634 6040 9007
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6000 8016 6052 8022
rect 6000 7958 6052 7964
rect 6012 6866 6040 7958
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 6104 2922 6132 9114
rect 6288 7954 6316 9438
rect 6472 8401 6500 9959
rect 6748 9042 6776 10118
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7116 9722 7144 10406
rect 7484 10266 7512 11086
rect 7576 10810 7604 11154
rect 7668 11082 7696 11766
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6458 8392 6514 8401
rect 6458 8327 6514 8336
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6092 2916 6144 2922
rect 6092 2858 6144 2864
rect 5170 2000 5226 2009
rect 5170 1935 5226 1944
rect 4122 1550 4200 1578
rect 4066 1527 4122 1536
rect 2884 1278 3004 1306
rect 2502 640 2558 649
rect 2502 575 2558 584
rect 2884 241 2912 1278
rect 6288 1222 6316 7890
rect 6932 7818 6960 8910
rect 7116 8294 7144 9318
rect 7392 9110 7420 9318
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7024 8090 7052 8230
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7208 7818 7236 8298
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 6932 7342 6960 7754
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 7484 4146 7512 10202
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9722 7880 9862
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7944 9518 7972 9998
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 8220 9382 8248 11630
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8496 10742 8524 11154
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8312 10198 8340 10610
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8312 9722 8340 10134
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8220 8974 8248 9318
rect 8496 9178 8524 10542
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8588 9110 8616 14844
rect 8668 14826 8720 14832
rect 8772 14278 8800 14962
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8680 12170 8708 12786
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8680 11558 8708 12106
rect 8772 11694 8800 14214
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8864 9625 8892 18527
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8956 17202 8984 17614
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8956 15978 8984 17138
rect 9048 17082 9076 18906
rect 9140 18426 9168 19790
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9232 18154 9260 19910
rect 9312 19236 9364 19242
rect 9364 19196 9444 19224
rect 9312 19178 9364 19184
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9140 17202 9168 17682
rect 9324 17610 9352 18022
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9048 17054 9168 17082
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9048 16046 9076 16526
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8944 15972 8996 15978
rect 8944 15914 8996 15920
rect 8956 15502 8984 15914
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8956 15026 8984 15438
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 9034 14920 9090 14929
rect 8944 14884 8996 14890
rect 9034 14855 9090 14864
rect 8944 14826 8996 14832
rect 8850 9616 8906 9625
rect 8850 9551 8906 9560
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8036 8566 8064 8910
rect 8024 8560 8076 8566
rect 8220 8514 8248 8910
rect 8024 8502 8076 8508
rect 8128 8486 8248 8514
rect 8128 8362 8156 8486
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 7576 7274 7604 8298
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8220 7818 8248 8366
rect 8312 8090 8340 8978
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8588 7342 8616 8502
rect 8864 8294 8892 9551
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8864 7274 8892 7822
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8956 6662 8984 14826
rect 9048 14822 9076 14855
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 13530 9076 13670
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9140 8090 9168 17054
rect 9416 16250 9444 19196
rect 9404 16244 9456 16250
rect 9232 16204 9404 16232
rect 9232 10169 9260 16204
rect 9404 16186 9456 16192
rect 9310 16008 9366 16017
rect 9310 15943 9312 15952
rect 9364 15943 9366 15952
rect 9312 15914 9364 15920
rect 9508 13818 9536 22000
rect 9772 20732 9824 20738
rect 9772 20674 9824 20680
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 19310 9628 19654
rect 9784 19310 9812 20674
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9692 18834 9720 19178
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9876 18714 9904 22000
rect 10336 20738 10364 22000
rect 10324 20732 10376 20738
rect 10324 20674 10376 20680
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10244 20058 10272 20334
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9692 18686 9904 18714
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9600 18426 9628 18566
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9588 17808 9640 17814
rect 9588 17750 9640 17756
rect 9600 17649 9628 17750
rect 9586 17640 9642 17649
rect 9586 17575 9642 17584
rect 9692 17218 9720 18686
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9770 18456 9826 18465
rect 9770 18391 9826 18400
rect 9784 18086 9812 18391
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9876 17882 9904 18566
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9692 17190 9812 17218
rect 9680 17128 9732 17134
rect 9586 17096 9642 17105
rect 9680 17070 9732 17076
rect 9586 17031 9642 17040
rect 9600 14074 9628 17031
rect 9692 16522 9720 17070
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9680 15088 9732 15094
rect 9678 15056 9680 15065
rect 9732 15056 9734 15065
rect 9678 14991 9734 15000
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9416 13802 9536 13818
rect 9404 13796 9536 13802
rect 9456 13790 9536 13796
rect 9404 13738 9456 13744
rect 9692 13394 9720 14894
rect 9784 14618 9812 17190
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9784 13258 9812 14554
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9600 12753 9628 12786
rect 9586 12744 9642 12753
rect 9586 12679 9642 12688
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12442 9720 12582
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 11150 9352 11494
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9324 10674 9352 11086
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9218 10160 9274 10169
rect 9218 10095 9274 10104
rect 9324 9518 9352 10610
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10266 9536 10406
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 9722 9444 9998
rect 9600 9994 9628 10678
rect 9876 10470 9904 17138
rect 9968 12442 9996 19246
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10060 18902 10088 19110
rect 10048 18896 10100 18902
rect 10048 18838 10100 18844
rect 10060 18290 10088 18838
rect 10152 18290 10180 19858
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10244 19378 10272 19790
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 17678 10088 18022
rect 10138 17776 10194 17785
rect 10244 17746 10272 19110
rect 10336 18902 10364 19790
rect 10416 19236 10468 19242
rect 10416 19178 10468 19184
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10428 18834 10456 19178
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10138 17711 10194 17720
rect 10232 17740 10284 17746
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 13462 10088 13670
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9956 12436 10008 12442
rect 10008 12396 10088 12424
rect 9956 12378 10008 12384
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9968 11762 9996 12174
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 10060 11694 10088 12396
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10152 11218 10180 17711
rect 10232 17682 10284 17688
rect 10324 17672 10376 17678
rect 10230 17640 10286 17649
rect 10324 17614 10376 17620
rect 10230 17575 10232 17584
rect 10284 17575 10286 17584
rect 10232 17546 10284 17552
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10244 16726 10272 16934
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10336 16658 10364 17614
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10230 16552 10286 16561
rect 10230 16487 10286 16496
rect 10244 15978 10272 16487
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10336 16153 10364 16186
rect 10322 16144 10378 16153
rect 10322 16079 10378 16088
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10244 13938 10272 14486
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10428 12714 10456 18362
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10520 13734 10548 16730
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10244 12345 10272 12650
rect 10230 12336 10286 12345
rect 10230 12271 10286 12280
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10060 11082 10088 11154
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9968 10198 9996 10542
rect 10152 10266 10180 10950
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9494 9616 9550 9625
rect 9494 9551 9496 9560
rect 9548 9551 9550 9560
rect 9496 9522 9548 9528
rect 10244 9518 10272 11290
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10336 9586 10364 11154
rect 10520 11014 10548 12174
rect 10612 11354 10640 18090
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10704 11218 10732 22000
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10784 19236 10836 19242
rect 10784 19178 10836 19184
rect 10796 18970 10824 19178
rect 10980 18970 11008 19246
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10796 16998 10824 17274
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10796 15978 10824 16934
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10888 15892 10916 18294
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 10980 17270 11008 17682
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 11072 17202 11100 19246
rect 11164 18426 11192 22000
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11532 18970 11560 19110
rect 11520 18964 11572 18970
rect 11520 18906 11572 18912
rect 11532 18766 11560 18906
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11164 17338 11192 18090
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11440 17882 11468 18022
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11242 17232 11298 17241
rect 11060 17196 11112 17202
rect 11242 17167 11298 17176
rect 11060 17138 11112 17144
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10980 16046 11008 17002
rect 11256 16998 11284 17167
rect 11428 17060 11480 17066
rect 11428 17002 11480 17008
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11242 16688 11298 16697
rect 11440 16674 11468 17002
rect 11298 16646 11468 16674
rect 11242 16623 11244 16632
rect 11296 16623 11298 16632
rect 11244 16594 11296 16600
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 11072 16114 11100 16458
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10968 16040 11020 16046
rect 10966 16008 10968 16017
rect 11020 16008 11022 16017
rect 10966 15943 11022 15952
rect 10888 15864 11008 15892
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10888 15162 10916 15506
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10796 14006 10824 14350
rect 10888 14074 10916 14350
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10796 11762 10824 12242
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10888 11354 10916 11766
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10606 10548 10950
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10598 10568 10654 10577
rect 10520 10062 10548 10542
rect 10598 10503 10600 10512
rect 10652 10503 10654 10512
rect 10600 10474 10652 10480
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9654 10916 9998
rect 10876 9648 10928 9654
rect 10506 9616 10562 9625
rect 10324 9580 10376 9586
rect 10876 9590 10928 9596
rect 10506 9551 10508 9560
rect 10324 9522 10376 9528
rect 10560 9551 10562 9560
rect 10508 9522 10560 9528
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9110 9536 9386
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 9178 9904 9318
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 10888 9042 10916 9590
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9586 8528 9642 8537
rect 9968 8498 9996 8842
rect 9586 8463 9642 8472
rect 9956 8492 10008 8498
rect 9600 8090 9628 8463
rect 9956 8434 10008 8440
rect 10980 8362 11008 15864
rect 11348 15638 11376 16118
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11520 14816 11572 14822
rect 11518 14784 11520 14793
rect 11572 14784 11574 14793
rect 11518 14719 11574 14728
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11072 8786 11100 14418
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11440 13530 11468 13874
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11532 13394 11560 13738
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 11626 11192 12582
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11518 11656 11574 11665
rect 11152 11620 11204 11626
rect 11518 11591 11520 11600
rect 11152 11562 11204 11568
rect 11572 11591 11574 11600
rect 11520 11562 11572 11568
rect 11336 11144 11388 11150
rect 11334 11112 11336 11121
rect 11388 11112 11390 11121
rect 11164 11070 11334 11098
rect 11164 10538 11192 11070
rect 11334 11047 11390 11056
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11624 9500 11652 22000
rect 11992 19310 12020 22000
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11992 18902 12020 19110
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11716 17490 11744 18362
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11808 17610 11836 18158
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11716 17462 11836 17490
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11716 15026 11744 16050
rect 11808 15042 11836 17462
rect 11900 17202 11928 17682
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 15994 11928 16934
rect 11992 16114 12020 18158
rect 12176 17610 12204 19858
rect 12268 19718 12296 20538
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12268 17542 12296 19246
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12176 16250 12204 16526
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11900 15966 12020 15994
rect 11886 15736 11942 15745
rect 11992 15722 12020 15966
rect 11992 15694 12112 15722
rect 11886 15671 11888 15680
rect 11940 15671 11942 15680
rect 11888 15642 11940 15648
rect 11886 15192 11942 15201
rect 11886 15127 11888 15136
rect 11940 15127 11942 15136
rect 11888 15098 11940 15104
rect 11704 15020 11756 15026
rect 11808 15014 11928 15042
rect 11704 14962 11756 14968
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11716 14618 11744 14826
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11716 13394 11744 13874
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11808 11694 11836 14758
rect 11900 13308 11928 15014
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 13462 12020 14214
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11900 13280 12020 13308
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11900 11898 11928 12174
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11808 11354 11836 11494
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11900 11200 11928 11698
rect 11808 11172 11928 11200
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11716 10130 11744 10678
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11624 9472 11744 9500
rect 11612 8832 11664 8838
rect 11072 8758 11192 8786
rect 11612 8774 11664 8780
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9968 8022 9996 8230
rect 10244 8090 10272 8230
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10336 8022 10364 8230
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 9968 7886 9996 7958
rect 10980 7954 11008 8298
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 9956 7880 10008 7886
rect 11072 7868 11100 8502
rect 11164 8362 11192 8758
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8498 11652 8774
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11716 8430 11744 9472
rect 11808 9110 11836 11172
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11900 10198 11928 10406
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11900 9761 11928 9862
rect 11886 9752 11942 9761
rect 11886 9687 11942 9696
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11716 7886 11744 8366
rect 11152 7880 11204 7886
rect 11072 7840 11152 7868
rect 9956 7822 10008 7828
rect 11152 7822 11204 7828
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11900 6225 11928 9386
rect 11992 8673 12020 13280
rect 12084 10266 12112 15694
rect 12268 15201 12296 16526
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12360 16250 12388 16390
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12360 15706 12388 15982
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12254 15192 12310 15201
rect 12254 15127 12310 15136
rect 12452 14482 12480 22000
rect 12820 19394 12848 22000
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 12544 19366 12848 19394
rect 12544 15065 12572 19366
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12728 18766 12756 18906
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12728 17746 12756 18294
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12636 17338 12664 17614
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12820 17202 12848 19178
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 19009 12940 19110
rect 12898 19000 12954 19009
rect 12898 18935 12954 18944
rect 13004 18426 13032 19858
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13096 19514 13124 19790
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12912 16182 12940 18294
rect 13096 18154 13124 19110
rect 13188 18970 13216 19790
rect 13280 19530 13308 22000
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13280 19502 13400 19530
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18426 13216 18702
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13280 18290 13308 19314
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 12992 18080 13044 18086
rect 12990 18048 12992 18057
rect 13044 18048 13046 18057
rect 12990 17983 13046 17992
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16658 13124 16934
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 12912 15910 12940 16118
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12530 15056 12586 15065
rect 12530 14991 12586 15000
rect 12544 14618 12572 14991
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12636 14362 12664 15302
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 13004 14793 13032 14826
rect 12990 14784 13046 14793
rect 13046 14742 13124 14770
rect 12990 14719 13046 14728
rect 13004 14659 13032 14719
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12544 14334 12664 14362
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12544 13870 12572 14334
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12544 13190 12572 13806
rect 12636 13530 12664 14214
rect 12728 14074 12756 14350
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12728 13870 12756 14010
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12912 13530 12940 14214
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12636 13410 12664 13466
rect 12636 13382 12756 13410
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12636 12714 12664 13262
rect 12728 13190 12756 13382
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11898 12480 12038
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12348 11688 12400 11694
rect 12400 11648 12480 11676
rect 12348 11630 12400 11636
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12268 10169 12296 11630
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 11286 12388 11494
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12452 11150 12480 11648
rect 12636 11558 12664 12650
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12360 10470 12388 11086
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10742 12480 10950
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12254 10160 12310 10169
rect 12084 10118 12254 10146
rect 12084 9160 12112 10118
rect 12254 10095 12310 10104
rect 12256 9920 12308 9926
rect 12162 9888 12218 9897
rect 12256 9862 12308 9868
rect 12162 9823 12218 9832
rect 12176 9722 12204 9823
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12084 9132 12204 9160
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11978 8664 12034 8673
rect 11978 8599 12034 8608
rect 11992 7954 12020 8599
rect 12084 8430 12112 8978
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 12176 6390 12204 9132
rect 12268 9110 12296 9862
rect 12360 9586 12388 10406
rect 12440 9920 12492 9926
rect 12438 9888 12440 9897
rect 12492 9888 12494 9897
rect 12438 9823 12494 9832
rect 12544 9654 12572 11222
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12636 10810 12664 11154
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12728 9518 12756 9998
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 12268 6458 12296 8298
rect 12360 7818 12388 8978
rect 12544 8650 12572 9114
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12452 8634 12572 8650
rect 12440 8628 12572 8634
rect 12492 8622 12572 8628
rect 12624 8628 12676 8634
rect 12440 8570 12492 8576
rect 12624 8570 12676 8576
rect 12636 8537 12664 8570
rect 12622 8528 12678 8537
rect 12622 8463 12678 8472
rect 12728 8362 12756 9046
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12544 7750 12572 7958
rect 13004 7954 13032 14418
rect 13096 14074 13124 14742
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 13096 12442 13124 12650
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13188 10606 13216 18090
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13280 12617 13308 17818
rect 13372 13326 13400 19502
rect 13450 17640 13506 17649
rect 13450 17575 13506 17584
rect 13464 17542 13492 17575
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17134 13492 17478
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13360 12640 13412 12646
rect 13266 12608 13322 12617
rect 13360 12582 13412 12588
rect 13266 12543 13322 12552
rect 13266 11112 13322 11121
rect 13266 11047 13322 11056
rect 13280 10674 13308 11047
rect 13372 10810 13400 12582
rect 13464 12442 13492 12786
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13556 10690 13584 19858
rect 13648 18154 13676 22000
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13832 19310 13860 19654
rect 13924 19514 13952 19654
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 14016 19394 14044 19858
rect 13924 19366 14044 19394
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13636 18148 13688 18154
rect 13636 18090 13688 18096
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13648 16998 13676 17614
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13636 16584 13688 16590
rect 13740 16572 13768 17138
rect 13924 17066 13952 19366
rect 14108 19242 14136 22000
rect 14372 20664 14424 20670
rect 14372 20606 14424 20612
rect 14384 20058 14412 20606
rect 14568 20482 14596 22000
rect 14476 20454 14596 20482
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14200 17270 14228 18770
rect 14476 18630 14504 20454
rect 14936 20346 14964 22000
rect 14556 20324 14608 20330
rect 14936 20318 15056 20346
rect 14556 20266 14608 20272
rect 14568 19786 14596 20266
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14844 19446 14872 19858
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14752 18222 14780 18634
rect 15028 18426 15056 20318
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15120 20058 15148 20198
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15108 19304 15160 19310
rect 15292 19304 15344 19310
rect 15160 19252 15240 19258
rect 15108 19246 15240 19252
rect 15292 19246 15344 19252
rect 15120 19230 15240 19246
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 15016 18148 15068 18154
rect 15016 18090 15068 18096
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14568 17270 14596 17818
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14936 17066 14964 17682
rect 15028 17678 15056 18090
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15212 17066 15240 19230
rect 15304 17882 15332 19246
rect 15396 19174 15424 22000
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15672 20058 15700 20402
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15488 19242 15516 19858
rect 15476 19236 15528 19242
rect 15476 19178 15528 19184
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15580 18902 15608 19926
rect 15764 19174 15792 22000
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15672 17882 15700 18566
rect 15764 18222 15792 18770
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 13912 17060 13964 17066
rect 13912 17002 13964 17008
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14924 17060 14976 17066
rect 14924 17002 14976 17008
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 13924 16726 13952 17002
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13688 16544 13768 16572
rect 13636 16526 13688 16532
rect 13648 16046 13676 16526
rect 14016 16522 14044 17002
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 14004 16516 14056 16522
rect 14004 16458 14056 16464
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13648 15366 13676 15982
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13818 15192 13874 15201
rect 13818 15127 13874 15136
rect 13832 15026 13860 15127
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13924 14890 13952 15914
rect 14016 15745 14044 16050
rect 14002 15736 14058 15745
rect 14002 15671 14058 15680
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13924 14618 13952 14826
rect 14016 14770 14044 15671
rect 14108 15094 14136 16934
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 15706 14320 16390
rect 14568 15978 14596 16526
rect 14660 16454 14688 16662
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14292 15162 14320 15506
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14384 15026 14412 15846
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 15028 14958 15056 16730
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14016 14742 14504 14770
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13648 11898 13676 12786
rect 13740 12714 13768 13670
rect 13832 13258 13860 14350
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 14108 12986 14136 14418
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13726 12608 13782 12617
rect 13726 12543 13782 12552
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13648 11286 13676 11834
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13268 10668 13320 10674
rect 13556 10662 13676 10690
rect 13268 10610 13320 10616
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13280 10062 13308 10610
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13372 9518 13400 9862
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13464 8498 13492 8842
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 13004 7478 13032 7890
rect 13280 7886 13308 8230
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 13648 6322 13676 10662
rect 13740 10198 13768 12543
rect 14108 12306 14136 12922
rect 14200 12782 14228 13806
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14384 13326 14412 13738
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 13924 12186 13952 12242
rect 14188 12232 14240 12238
rect 13924 12158 14136 12186
rect 14188 12174 14240 12180
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13924 11218 13952 12038
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13740 9178 13768 10134
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13832 8906 13860 9386
rect 13924 9382 13952 11154
rect 14016 10606 14044 12038
rect 14108 11898 14136 12158
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14200 11626 14228 12174
rect 14384 12102 14412 12854
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14476 11744 14504 14742
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 15120 14618 15148 16594
rect 15580 16250 15608 16934
rect 15764 16658 15792 18158
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15856 17678 15884 18090
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15198 16144 15254 16153
rect 15198 16079 15254 16088
rect 15212 15978 15240 16079
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15292 13728 15344 13734
rect 15290 13696 15292 13705
rect 15344 13696 15346 13705
rect 14684 13628 14980 13648
rect 15290 13631 15346 13640
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14660 11762 14688 12106
rect 14292 11716 14504 11744
rect 14648 11756 14700 11762
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14016 9994 14044 10406
rect 14108 10062 14136 11018
rect 14200 10674 14228 11562
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 14108 8634 14136 8910
rect 14292 8906 14320 11716
rect 14648 11698 14700 11704
rect 15016 11688 15068 11694
rect 14476 11626 14688 11642
rect 15200 11688 15252 11694
rect 15016 11630 15068 11636
rect 15198 11656 15200 11665
rect 15252 11656 15254 11665
rect 14476 11620 14700 11626
rect 14476 11614 14648 11620
rect 14476 9042 14504 11614
rect 14648 11562 14700 11568
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15028 10713 15056 11630
rect 15198 11591 15254 11600
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15014 10704 15070 10713
rect 15014 10639 15070 10648
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14568 10062 14596 10542
rect 15016 10532 15068 10538
rect 15016 10474 15068 10480
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14648 9988 14700 9994
rect 14648 9930 14700 9936
rect 14660 9586 14688 9930
rect 15028 9625 15056 10474
rect 15120 10470 15148 11494
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15014 9616 15070 9625
rect 14648 9580 14700 9586
rect 15014 9551 15070 9560
rect 14648 9522 14700 9528
rect 15212 9518 15240 9998
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 15028 8974 15056 9386
rect 15304 9194 15332 13398
rect 15396 12374 15424 13806
rect 15488 13734 15516 14282
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 12782 15516 13670
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15474 12608 15530 12617
rect 15474 12543 15530 12552
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15488 11558 15516 12543
rect 15580 11801 15608 16186
rect 15752 15360 15804 15366
rect 15856 15314 15884 16526
rect 15948 15570 15976 16594
rect 16040 16250 16068 17138
rect 16224 16250 16252 22000
rect 16684 20602 16712 22000
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 17052 20330 17080 22000
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 17512 20058 17540 22000
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 16856 19984 16908 19990
rect 16856 19926 16908 19932
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16040 15638 16068 16186
rect 16316 16130 16344 18158
rect 16592 17202 16620 19246
rect 16684 19242 16712 19858
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16776 17882 16804 19178
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16868 17218 16896 19926
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 16960 18902 16988 19110
rect 16948 18896 17000 18902
rect 16948 18838 17000 18844
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 17052 18426 17080 18770
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16776 17190 16896 17218
rect 16224 16102 16344 16130
rect 16028 15632 16080 15638
rect 16028 15574 16080 15580
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15804 15308 15884 15314
rect 15752 15302 15884 15308
rect 15764 15286 15884 15302
rect 15856 15026 15884 15286
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15844 14816 15896 14822
rect 15948 14804 15976 15506
rect 16028 14816 16080 14822
rect 15948 14776 16028 14804
rect 15844 14758 15896 14764
rect 16028 14758 16080 14764
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 13258 15700 14418
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15764 13326 15792 13670
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15566 11792 15622 11801
rect 15672 11762 15700 12922
rect 15856 12918 15884 14758
rect 16040 14414 16068 14758
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16040 14074 16068 14350
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15566 11727 15622 11736
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15382 10432 15438 10441
rect 15382 10367 15438 10376
rect 15396 10033 15424 10367
rect 15382 10024 15438 10033
rect 15382 9959 15438 9968
rect 15304 9166 15424 9194
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8634 14228 8774
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7750 13952 8230
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 14292 6730 14320 8842
rect 15304 8294 15332 8978
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15028 8090 15056 8230
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 15396 8022 15424 9166
rect 15488 8634 15516 11494
rect 15764 11234 15792 12174
rect 15764 11218 15884 11234
rect 15764 11212 15896 11218
rect 15764 11206 15844 11212
rect 15844 11154 15896 11160
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15764 9042 15792 10134
rect 15856 10062 15884 11154
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15580 8294 15608 8570
rect 15672 8498 15700 8842
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15764 8022 15792 8774
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15856 7886 15884 9386
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15948 7750 15976 14010
rect 16132 13870 16160 14486
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 12850 16068 13670
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16132 12986 16160 13126
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16224 12442 16252 16102
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16592 14958 16620 15370
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16316 13938 16344 14214
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16316 13326 16344 13874
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16408 13530 16436 13738
rect 16500 13530 16528 14010
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16500 13326 16528 13466
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16316 12238 16344 12718
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16040 11218 16068 11698
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 11257 16344 11494
rect 16408 11354 16436 12854
rect 16592 12850 16620 13398
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16488 11552 16540 11558
rect 16684 11529 16712 13330
rect 16776 11762 16804 17190
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16868 16250 16896 17070
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16960 16130 16988 17818
rect 17052 17678 17080 18362
rect 17236 17882 17264 19110
rect 17420 18970 17448 19246
rect 17512 18970 17540 19314
rect 17696 19258 17724 20334
rect 17604 19242 17724 19258
rect 17604 19236 17736 19242
rect 17604 19230 17684 19236
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 16868 16102 16988 16130
rect 16868 12345 16896 16102
rect 17052 15978 17080 16186
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 17052 13938 17080 15302
rect 17144 14006 17172 17682
rect 17224 17060 17276 17066
rect 17224 17002 17276 17008
rect 17236 16046 17264 17002
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17236 13954 17264 15302
rect 17328 14074 17356 15846
rect 17420 14113 17448 18906
rect 17512 18154 17540 18906
rect 17500 18148 17552 18154
rect 17500 18090 17552 18096
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 17512 16794 17540 17206
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17498 16008 17554 16017
rect 17498 15943 17554 15952
rect 17512 15638 17540 15943
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17604 15366 17632 19230
rect 17684 19178 17736 19184
rect 17682 19136 17738 19145
rect 17682 19071 17738 19080
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17406 14104 17462 14113
rect 17316 14068 17368 14074
rect 17406 14039 17462 14048
rect 17316 14010 17368 14016
rect 17040 13932 17092 13938
rect 17236 13926 17356 13954
rect 17040 13874 17092 13880
rect 17222 13832 17278 13841
rect 17222 13767 17278 13776
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16960 12714 16988 13466
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16854 12336 16910 12345
rect 16854 12271 16910 12280
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16960 11626 16988 12650
rect 17236 12374 17264 13767
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17052 11898 17080 12310
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17144 11898 17172 12242
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 16488 11494 16540 11500
rect 16670 11520 16726 11529
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16302 11248 16358 11257
rect 16028 11212 16080 11218
rect 16302 11183 16358 11192
rect 16028 11154 16080 11160
rect 16040 11121 16068 11154
rect 16026 11112 16082 11121
rect 16026 11047 16082 11056
rect 16040 10810 16068 11047
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16120 10056 16172 10062
rect 16172 10016 16252 10044
rect 16120 9998 16172 10004
rect 16224 9586 16252 10016
rect 16408 9722 16436 11290
rect 16500 10810 16528 11494
rect 16670 11455 16726 11464
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16592 9654 16620 10134
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 16040 9178 16068 9386
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16408 8838 16436 9454
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16316 8090 16344 8774
rect 16408 8294 16436 8774
rect 16684 8634 16712 11455
rect 17144 11354 17172 11834
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17328 11014 17356 13926
rect 17512 13682 17540 14826
rect 17604 14482 17632 15030
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 13977 17632 14418
rect 17696 14278 17724 19071
rect 17788 18426 17816 22471
rect 17866 22000 17922 22800
rect 18326 22000 18382 22800
rect 18510 22128 18566 22137
rect 18510 22063 18566 22072
rect 17880 20466 17908 22000
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 18340 19786 18368 22000
rect 18524 20058 18552 22063
rect 18786 22000 18842 22800
rect 19154 22000 19210 22800
rect 19614 22000 19670 22800
rect 19982 22000 20038 22800
rect 20442 22000 20498 22800
rect 20902 22000 20958 22800
rect 21270 22000 21326 22800
rect 21730 22000 21786 22800
rect 22098 22000 22154 22800
rect 22558 22000 22614 22800
rect 18602 21584 18658 21593
rect 18602 21519 18658 21528
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17972 18902 18000 19654
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17972 18057 18000 18158
rect 17958 18048 18014 18057
rect 17958 17983 18014 17992
rect 18524 17746 18552 19858
rect 18616 19174 18644 21519
rect 18800 19854 18828 22000
rect 19062 21176 19118 21185
rect 19062 21111 19118 21120
rect 19076 20058 19104 21111
rect 19168 20262 19196 22000
rect 19628 20670 19656 22000
rect 19616 20664 19668 20670
rect 19246 20632 19302 20641
rect 19616 20606 19668 20612
rect 19246 20567 19302 20576
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19260 20058 19288 20567
rect 19614 20224 19670 20233
rect 19614 20159 19670 20168
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18616 17678 18644 18158
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18602 17368 18658 17377
rect 17868 17332 17920 17338
rect 18602 17303 18658 17312
rect 17868 17274 17920 17280
rect 17880 16794 17908 17274
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17866 16552 17922 16561
rect 17866 16487 17922 16496
rect 17880 16454 17908 16487
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17788 15434 17816 16390
rect 17972 15706 18000 17002
rect 18340 16726 18368 17138
rect 18616 16794 18644 17303
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17776 15428 17828 15434
rect 18064 15416 18092 16050
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18510 16008 18566 16017
rect 18432 15722 18460 15982
rect 18510 15943 18566 15952
rect 18604 15972 18656 15978
rect 18524 15910 18552 15943
rect 18604 15914 18656 15920
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18432 15694 18552 15722
rect 17776 15370 17828 15376
rect 17972 15388 18092 15416
rect 17972 14890 18000 15388
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17880 14618 17908 14758
rect 17972 14618 18000 14826
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17776 14544 17828 14550
rect 17776 14486 17828 14492
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17590 13968 17646 13977
rect 17590 13903 17592 13912
rect 17644 13903 17646 13912
rect 17592 13874 17644 13880
rect 17512 13654 17632 13682
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 12442 17540 12786
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 16856 10192 16908 10198
rect 16776 10140 16856 10146
rect 16776 10134 16908 10140
rect 16776 10118 16896 10134
rect 16776 9178 16804 10118
rect 17052 9761 17080 10542
rect 17328 10198 17356 10950
rect 17500 10532 17552 10538
rect 17500 10474 17552 10480
rect 17512 10266 17540 10474
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17038 9752 17094 9761
rect 17038 9687 17094 9696
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16868 9382 16896 9454
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16868 7818 16896 9114
rect 16946 8664 17002 8673
rect 16946 8599 17002 8608
rect 16960 8430 16988 8599
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 17052 8378 17080 9522
rect 17604 9489 17632 13654
rect 17682 12608 17738 12617
rect 17682 12543 17738 12552
rect 17590 9480 17646 9489
rect 17590 9415 17646 9424
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17236 9178 17264 9318
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17512 8634 17540 8842
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17132 8424 17184 8430
rect 17052 8372 17132 8378
rect 17052 8366 17184 8372
rect 17052 8350 17172 8366
rect 17052 7886 17080 8350
rect 17236 8022 17264 8434
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 17052 6934 17080 7822
rect 17236 7410 17264 7958
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17236 7002 17264 7346
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17040 6928 17092 6934
rect 17040 6870 17092 6876
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 9494 6216 9550 6225
rect 9494 6151 9550 6160
rect 11886 6216 11942 6225
rect 11886 6151 11942 6160
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 2964 1216 3016 1222
rect 2964 1158 3016 1164
rect 6276 1216 6328 1222
rect 6276 1158 6328 1164
rect 2976 1057 3004 1158
rect 2962 1048 3018 1057
rect 2962 983 3018 992
rect 6748 800 6776 4082
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 9508 2836 9536 6151
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9508 2808 9720 2836
rect 9692 2802 9720 2808
rect 9784 2802 9812 2858
rect 9692 2774 9812 2802
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 11164 1442 11192 2926
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11164 1414 11376 1442
rect 11348 800 11376 1414
rect 15856 800 15884 2926
rect 17420 2553 17448 8570
rect 17696 7546 17724 12543
rect 17788 12442 17816 14486
rect 18064 14328 18092 15030
rect 17972 14300 18092 14328
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17880 12374 17908 12922
rect 17972 12918 18000 14300
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18524 13394 18552 15694
rect 18616 14074 18644 15914
rect 18708 15706 18736 18838
rect 18800 18698 18828 19246
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18788 18692 18840 18698
rect 18788 18634 18840 18640
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18800 18057 18828 18158
rect 18786 18048 18842 18057
rect 18786 17983 18842 17992
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18800 16590 18828 17478
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18892 16794 18920 17138
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18800 16046 18828 16526
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18708 14482 18736 14758
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18696 14340 18748 14346
rect 18696 14282 18748 14288
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18602 13968 18658 13977
rect 18602 13903 18604 13912
rect 18656 13903 18658 13912
rect 18604 13874 18656 13880
rect 18708 13802 18736 14282
rect 18800 13818 18828 14894
rect 18892 14804 18920 15302
rect 18984 14906 19012 18770
rect 19340 18760 19392 18766
rect 19260 18708 19340 18714
rect 19260 18702 19392 18708
rect 19260 18686 19380 18702
rect 19260 18290 19288 18686
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19260 18086 19288 18226
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19260 17814 19288 18022
rect 19248 17808 19300 17814
rect 19248 17750 19300 17756
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 19168 17105 19196 17206
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19154 17096 19210 17105
rect 19154 17031 19210 17040
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 19076 15026 19104 16594
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 18984 14878 19104 14906
rect 18892 14776 19012 14804
rect 18878 14648 18934 14657
rect 18878 14583 18880 14592
rect 18932 14583 18934 14592
rect 18880 14554 18932 14560
rect 18696 13796 18748 13802
rect 18800 13790 18920 13818
rect 18696 13738 18748 13744
rect 18788 13728 18840 13734
rect 18788 13670 18840 13676
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18708 13394 18736 13466
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 17960 12912 18012 12918
rect 17960 12854 18012 12860
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17868 11620 17920 11626
rect 17868 11562 17920 11568
rect 17774 10568 17830 10577
rect 17774 10503 17830 10512
rect 17788 10266 17816 10503
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17880 9874 17908 11562
rect 17972 10674 18000 12242
rect 18432 12209 18460 12650
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18418 12200 18474 12209
rect 18418 12135 18474 12144
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18248 11150 18276 11698
rect 18236 11144 18288 11150
rect 18234 11112 18236 11121
rect 18288 11112 18290 11121
rect 18234 11047 18290 11056
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 18234 10568 18290 10577
rect 18234 10503 18290 10512
rect 18142 10160 18198 10169
rect 18248 10130 18276 10503
rect 18524 10266 18552 12310
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18616 11762 18644 12174
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 11354 18736 11494
rect 18800 11393 18828 13670
rect 18786 11384 18842 11393
rect 18696 11348 18748 11354
rect 18786 11319 18842 11328
rect 18696 11290 18748 11296
rect 18694 11248 18750 11257
rect 18604 11212 18656 11218
rect 18694 11183 18696 11192
rect 18604 11154 18656 11160
rect 18748 11183 18750 11192
rect 18696 11154 18748 11160
rect 18616 10810 18644 11154
rect 18694 10840 18750 10849
rect 18604 10804 18656 10810
rect 18694 10775 18750 10784
rect 18604 10746 18656 10752
rect 18602 10704 18658 10713
rect 18602 10639 18604 10648
rect 18656 10639 18658 10648
rect 18604 10610 18656 10616
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18142 10095 18198 10104
rect 18236 10124 18288 10130
rect 18156 10062 18184 10095
rect 18236 10066 18288 10072
rect 18144 10056 18196 10062
rect 17958 10024 18014 10033
rect 18144 9998 18196 10004
rect 17958 9959 17960 9968
rect 18012 9959 18014 9968
rect 17960 9930 18012 9936
rect 17880 9846 18000 9874
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8430 17908 8910
rect 17972 8537 18000 9846
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18524 8945 18552 9658
rect 18510 8936 18566 8945
rect 18510 8871 18566 8880
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18052 8560 18104 8566
rect 17958 8528 18014 8537
rect 18616 8514 18644 10610
rect 18708 10606 18736 10775
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18052 8502 18104 8508
rect 17958 8463 18014 8472
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 18064 8090 18092 8502
rect 18524 8486 18644 8514
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17972 6769 18000 7686
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18524 7342 18552 8486
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18616 7818 18644 8298
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18708 7206 18736 10406
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18800 9081 18828 9862
rect 18786 9072 18842 9081
rect 18786 9007 18842 9016
rect 18786 8936 18842 8945
rect 18786 8871 18842 8880
rect 18696 7200 18748 7206
rect 18800 7177 18828 8871
rect 18892 7585 18920 13790
rect 18984 8129 19012 14776
rect 19076 13705 19104 14878
rect 19062 13696 19118 13705
rect 19062 13631 19118 13640
rect 19076 12753 19104 13631
rect 19168 13297 19196 16934
rect 19260 16658 19288 17138
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16250 19288 16594
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19260 15502 19288 16186
rect 19444 15722 19472 19722
rect 19536 18426 19564 19858
rect 19628 19514 19656 20159
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19628 17320 19656 19246
rect 19996 18850 20024 22000
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20166 19816 20222 19825
rect 20166 19751 20168 19760
rect 20220 19751 20222 19760
rect 20168 19722 20220 19728
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19904 18822 20024 18850
rect 19720 18426 19748 18770
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19904 18329 19932 18822
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19890 18320 19946 18329
rect 19890 18255 19946 18264
rect 19996 17542 20024 18702
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19536 17292 19656 17320
rect 19536 17134 19564 17292
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19352 15694 19472 15722
rect 19536 15706 19564 16934
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 19524 15700 19576 15706
rect 19352 15570 19380 15694
rect 19524 15642 19576 15648
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19352 15314 19380 15506
rect 19628 15502 19656 15914
rect 19720 15638 19748 16934
rect 19708 15632 19760 15638
rect 19708 15574 19760 15580
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19260 15286 19380 15314
rect 19154 13288 19210 13297
rect 19154 13223 19210 13232
rect 19260 12889 19288 15286
rect 19628 15162 19656 15438
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 19812 15008 19840 17478
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19996 16046 20024 16390
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 20088 15722 20116 19246
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20180 18873 20208 19110
rect 20166 18864 20222 18873
rect 20166 18799 20222 18808
rect 20272 17864 20300 19858
rect 20456 19009 20484 22000
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20442 19000 20498 19009
rect 20442 18935 20498 18944
rect 20548 17921 20576 19110
rect 20640 18329 20668 19654
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20626 18320 20682 18329
rect 20626 18255 20682 18264
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20180 17836 20300 17864
rect 20534 17912 20590 17921
rect 20534 17847 20590 17856
rect 20180 15978 20208 17836
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 19996 15694 20116 15722
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19536 14980 19840 15008
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19352 14074 19380 14350
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19444 13462 19472 13874
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19444 12986 19472 13398
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19246 12880 19302 12889
rect 19536 12866 19564 14980
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19616 13796 19668 13802
rect 19616 13738 19668 13744
rect 19246 12815 19302 12824
rect 19352 12838 19564 12866
rect 19062 12744 19118 12753
rect 19062 12679 19118 12688
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19154 12200 19210 12209
rect 19154 12135 19210 12144
rect 19168 11898 19196 12135
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19154 11520 19210 11529
rect 19154 11455 19210 11464
rect 19168 11354 19196 11455
rect 19260 11354 19288 12582
rect 19352 12322 19380 12838
rect 19628 12442 19656 13738
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19352 12294 19472 12322
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19248 11144 19300 11150
rect 19168 11104 19248 11132
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 19076 10266 19104 11018
rect 19168 10674 19196 11104
rect 19248 11086 19300 11092
rect 19352 10810 19380 11630
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19168 10198 19196 10610
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 18970 8120 19026 8129
rect 18970 8055 19026 8064
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18878 7576 18934 7585
rect 18984 7546 19012 7890
rect 18878 7511 18934 7520
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 19076 7478 19104 10066
rect 19168 9994 19196 10134
rect 19156 9988 19208 9994
rect 19156 9930 19208 9936
rect 19260 9874 19288 10542
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19352 10130 19380 10406
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19168 9846 19288 9874
rect 19168 8362 19196 9846
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 18880 7200 18932 7206
rect 18696 7142 18748 7148
rect 18786 7168 18842 7177
rect 18880 7142 18932 7148
rect 18786 7103 18842 7112
rect 18788 6792 18840 6798
rect 17958 6760 18014 6769
rect 18788 6734 18840 6740
rect 17958 6695 18014 6704
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 5817 18000 6598
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 17958 5808 18014 5817
rect 17958 5743 18014 5752
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17972 4865 18000 5306
rect 18524 5273 18552 6394
rect 18800 6322 18828 6734
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 17958 4856 18014 4865
rect 17958 4791 18014 4800
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 17406 2544 17462 2553
rect 17406 2479 17462 2488
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 2870 232 2926 241
rect 2870 167 2926 176
rect 6734 0 6790 800
rect 11334 0 11390 800
rect 15842 0 15898 800
rect 18892 241 18920 7142
rect 18984 1057 19012 7278
rect 18970 1048 19026 1057
rect 18970 983 19026 992
rect 19076 649 19104 7414
rect 19168 2961 19196 8298
rect 19260 7546 19288 9454
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8634 19380 8978
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19352 7478 19380 8570
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19444 6866 19472 12294
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19536 11694 19564 12038
rect 19720 11898 19748 13670
rect 19812 13530 19840 14350
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19904 13394 19932 15506
rect 19996 14074 20024 15694
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20088 14618 20116 15506
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19996 12986 20024 13670
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19536 10538 19564 11494
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19628 10606 19656 11154
rect 19720 11150 19748 11698
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 19720 10062 19748 10746
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19536 7546 19564 9318
rect 19628 9110 19656 9454
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19812 8838 19840 10134
rect 19904 10112 19932 11494
rect 19996 11354 20024 11766
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19984 10124 20036 10130
rect 19904 10084 19984 10112
rect 19984 10066 20036 10072
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19628 7342 19656 8230
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 7410 19748 7686
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19812 6254 19840 8774
rect 19904 7410 19932 9318
rect 19996 8430 20024 10066
rect 20088 9450 20116 14418
rect 20180 14074 20208 14486
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20180 10538 20208 12174
rect 20272 10810 20300 17682
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20364 15609 20392 16934
rect 20456 16561 20484 17478
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20442 16552 20498 16561
rect 20442 16487 20498 16496
rect 20548 15638 20576 17070
rect 20640 16969 20668 18022
rect 20732 17882 20760 18702
rect 20916 18193 20944 22000
rect 21284 18737 21312 22000
rect 21270 18728 21326 18737
rect 21270 18663 21326 18672
rect 20996 18216 21048 18222
rect 20902 18184 20958 18193
rect 20812 18148 20864 18154
rect 20996 18158 21048 18164
rect 20902 18119 20958 18128
rect 20812 18090 20864 18096
rect 20824 17882 20852 18090
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 21008 17270 21036 18158
rect 21744 17814 21772 22000
rect 21822 19272 21878 19281
rect 22112 19242 22140 22000
rect 21822 19207 21878 19216
rect 22100 19236 22152 19242
rect 21836 19122 21864 19207
rect 22100 19178 22152 19184
rect 22572 19122 22600 22000
rect 21836 19094 22600 19122
rect 21732 17808 21784 17814
rect 21732 17750 21784 17756
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20626 16960 20682 16969
rect 20626 16895 20682 16904
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20536 15632 20588 15638
rect 20350 15600 20406 15609
rect 20536 15574 20588 15580
rect 20350 15535 20406 15544
rect 20640 15065 20668 15846
rect 20626 15056 20682 15065
rect 20626 14991 20682 15000
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20456 14113 20484 14214
rect 20442 14104 20498 14113
rect 20442 14039 20498 14048
rect 20442 13696 20498 13705
rect 20442 13631 20498 13640
rect 20456 13530 20484 13631
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20364 12186 20392 12786
rect 20718 12608 20774 12617
rect 20718 12543 20774 12552
rect 20732 12442 20760 12543
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20444 12232 20496 12238
rect 20364 12180 20444 12186
rect 20364 12174 20496 12180
rect 20364 12158 20484 12174
rect 20456 11762 20484 12158
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 20824 10674 20852 13330
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20916 12442 20944 12650
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 20260 10532 20312 10538
rect 20260 10474 20312 10480
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 20180 9382 20208 10474
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 20088 8566 20116 9114
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 20088 8242 20116 8502
rect 19996 8214 20116 8242
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19720 5370 19748 6054
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19812 5234 19840 5510
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19996 3505 20024 8214
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20088 6458 20116 6598
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20076 6248 20128 6254
rect 20076 6190 20128 6196
rect 19982 3496 20038 3505
rect 19982 3431 20038 3440
rect 19154 2952 19210 2961
rect 19154 2887 19210 2896
rect 20088 1601 20116 6190
rect 20180 3913 20208 9318
rect 20272 8022 20300 10474
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 9178 20392 10406
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20548 9450 20576 9658
rect 20640 9654 20668 10542
rect 21008 10538 21036 15914
rect 20996 10532 21048 10538
rect 20996 10474 21048 10480
rect 21100 9722 21128 15982
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20640 8498 20668 9386
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20352 8356 20404 8362
rect 20352 8298 20404 8304
rect 20364 8090 20392 8298
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20640 7886 20668 8434
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20640 7342 20668 7686
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20364 6186 20392 6598
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20352 6180 20404 6186
rect 20352 6122 20404 6128
rect 20364 5710 20392 6122
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20272 4321 20300 5646
rect 20456 5234 20484 6394
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20548 5166 20576 6054
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20258 4312 20314 4321
rect 20258 4247 20314 4256
rect 20166 3904 20222 3913
rect 20166 3839 20222 3848
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20074 1592 20130 1601
rect 20074 1527 20130 1536
rect 20456 800 20484 2994
rect 20732 2009 20760 8230
rect 20718 2000 20774 2009
rect 20718 1935 20774 1944
rect 19062 640 19118 649
rect 19062 575 19118 584
rect 18878 232 18934 241
rect 18878 167 18934 176
rect 20442 0 20498 800
<< via2 >>
rect 3054 22480 3110 22536
rect 2778 22072 2834 22128
rect 1950 19760 2006 19816
rect 2042 19216 2098 19272
rect 1950 18808 2006 18864
rect 1950 16940 1952 16960
rect 1952 16940 2004 16960
rect 2004 16940 2006 16960
rect 1950 16904 2006 16940
rect 1950 16516 2006 16552
rect 1950 16496 1952 16516
rect 1952 16496 2004 16516
rect 2004 16496 2006 16516
rect 2134 18708 2136 18728
rect 2136 18708 2188 18728
rect 2188 18708 2190 18728
rect 2134 18672 2190 18708
rect 2962 21528 3018 21584
rect 2870 20576 2926 20632
rect 2778 19080 2834 19136
rect 2594 18808 2650 18864
rect 17774 22480 17830 22536
rect 3514 20168 3570 20224
rect 3146 18264 3202 18320
rect 2134 17620 2136 17640
rect 2136 17620 2188 17640
rect 2188 17620 2190 17640
rect 2134 17584 2190 17620
rect 2778 17332 2834 17368
rect 2778 17312 2780 17332
rect 2780 17312 2832 17332
rect 2832 17312 2834 17332
rect 1950 15544 2006 15600
rect 1950 15000 2006 15056
rect 1766 14864 1822 14920
rect 1858 14048 1914 14104
rect 2502 15952 2558 16008
rect 2870 14592 2926 14648
rect 3054 17856 3110 17912
rect 3606 18128 3662 18184
rect 3238 16904 3294 16960
rect 2870 13640 2926 13696
rect 3054 13232 3110 13288
rect 1122 4256 1178 4312
rect 2686 7520 2742 7576
rect 2870 2488 2926 2544
rect 4066 21120 4122 21176
rect 3974 18300 3976 18320
rect 3976 18300 4028 18320
rect 4028 18300 4030 18320
rect 3974 18264 4030 18300
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 5170 17448 5226 17504
rect 5354 18692 5410 18728
rect 5354 18672 5356 18692
rect 5356 18672 5408 18692
rect 5408 18672 5410 18692
rect 4986 15680 5042 15736
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 3790 11328 3846 11384
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4066 12316 4068 12336
rect 4068 12316 4120 12336
rect 4120 12316 4122 12336
rect 4066 12280 4122 12316
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4066 11736 4122 11792
rect 4066 10784 4122 10840
rect 4066 10376 4122 10432
rect 3974 9424 4030 9480
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4066 8472 4122 8528
rect 4066 8064 4122 8120
rect 4066 7112 4122 7168
rect 4066 6704 4122 6760
rect 3422 5752 3478 5808
rect 3974 5244 3976 5264
rect 3976 5244 4028 5264
rect 4028 5244 4030 5264
rect 3974 5208 4030 5244
rect 4066 4800 4122 4856
rect 3238 3440 3294 3496
rect 4066 1536 4122 1592
rect 4618 8336 4674 8392
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4802 6160 4858 6216
rect 4710 3848 4766 3904
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 5170 15408 5226 15464
rect 5078 11736 5134 11792
rect 5446 16632 5502 16688
rect 5538 15952 5594 16008
rect 6366 18400 6422 18456
rect 5354 11464 5410 11520
rect 6458 17040 6514 17096
rect 6550 16904 6606 16960
rect 6366 14864 6422 14920
rect 4986 2896 5042 2952
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5906 11736 5962 11792
rect 5998 9560 6054 9616
rect 6826 17720 6882 17776
rect 6918 13232 6974 13288
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 8850 18536 8906 18592
rect 8022 17176 8078 17232
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 8114 13252 8170 13288
rect 8114 13232 8116 13252
rect 8116 13232 8168 13252
rect 8168 13232 8170 13252
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 6458 9968 6514 10024
rect 5998 9016 6054 9072
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 6458 8336 6514 8392
rect 5170 1944 5226 2000
rect 2502 584 2558 640
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 9034 14864 9090 14920
rect 8850 9560 8906 9616
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 9310 15972 9366 16008
rect 9310 15952 9312 15972
rect 9312 15952 9364 15972
rect 9364 15952 9366 15972
rect 9586 17584 9642 17640
rect 9770 18400 9826 18456
rect 9586 17040 9642 17096
rect 9678 15036 9680 15056
rect 9680 15036 9732 15056
rect 9732 15036 9734 15056
rect 9678 15000 9734 15036
rect 9586 12688 9642 12744
rect 9218 10104 9274 10160
rect 10138 17720 10194 17776
rect 10230 17604 10286 17640
rect 10230 17584 10232 17604
rect 10232 17584 10284 17604
rect 10284 17584 10286 17604
rect 10230 16496 10286 16552
rect 10322 16088 10378 16144
rect 10230 12280 10286 12336
rect 9494 9580 9550 9616
rect 9494 9560 9496 9580
rect 9496 9560 9548 9580
rect 9548 9560 9550 9580
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11242 17176 11298 17232
rect 11242 16652 11298 16688
rect 11242 16632 11244 16652
rect 11244 16632 11296 16652
rect 11296 16632 11298 16652
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 10966 15988 10968 16008
rect 10968 15988 11020 16008
rect 11020 15988 11022 16008
rect 10966 15952 11022 15988
rect 10598 10532 10654 10568
rect 10598 10512 10600 10532
rect 10600 10512 10652 10532
rect 10652 10512 10654 10532
rect 10506 9580 10562 9616
rect 10506 9560 10508 9580
rect 10508 9560 10560 9580
rect 10560 9560 10562 9580
rect 9586 8472 9642 8528
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11518 14764 11520 14784
rect 11520 14764 11572 14784
rect 11572 14764 11574 14784
rect 11518 14728 11574 14764
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11518 11620 11574 11656
rect 11518 11600 11520 11620
rect 11520 11600 11572 11620
rect 11572 11600 11574 11620
rect 11334 11092 11336 11112
rect 11336 11092 11388 11112
rect 11388 11092 11390 11112
rect 11334 11056 11390 11092
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11886 15700 11942 15736
rect 11886 15680 11888 15700
rect 11888 15680 11940 15700
rect 11940 15680 11942 15700
rect 11886 15156 11942 15192
rect 11886 15136 11888 15156
rect 11888 15136 11940 15156
rect 11940 15136 11942 15156
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11886 9696 11942 9752
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 12254 15136 12310 15192
rect 12898 18944 12954 19000
rect 12990 18028 12992 18048
rect 12992 18028 13044 18048
rect 13044 18028 13046 18048
rect 12990 17992 13046 18028
rect 12530 15000 12586 15056
rect 12990 14728 13046 14784
rect 12254 10104 12310 10160
rect 12162 9832 12218 9888
rect 11978 8608 12034 8664
rect 12438 9868 12440 9888
rect 12440 9868 12492 9888
rect 12492 9868 12494 9888
rect 12438 9832 12494 9868
rect 12622 8472 12678 8528
rect 13450 17584 13506 17640
rect 13266 12552 13322 12608
rect 13266 11056 13322 11112
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 13818 15136 13874 15192
rect 14002 15680 14058 15736
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 13726 12552 13782 12608
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 15198 16088 15254 16144
rect 15290 13676 15292 13696
rect 15292 13676 15344 13696
rect 15344 13676 15346 13696
rect 15290 13640 15346 13676
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 15198 11636 15200 11656
rect 15200 11636 15252 11656
rect 15252 11636 15254 11656
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 15198 11600 15254 11636
rect 15014 10648 15070 10704
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 15014 9560 15070 9616
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 15474 12552 15530 12608
rect 15566 11736 15622 11792
rect 15382 10376 15438 10432
rect 15382 9968 15438 10024
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 17498 15952 17554 16008
rect 17682 19080 17738 19136
rect 17406 14048 17462 14104
rect 17222 13776 17278 13832
rect 16854 12280 16910 12336
rect 16302 11192 16358 11248
rect 16026 11056 16082 11112
rect 16670 11464 16726 11520
rect 18510 22072 18566 22128
rect 18602 21528 18658 21584
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 17958 17992 18014 18048
rect 19062 21120 19118 21176
rect 19246 20576 19302 20632
rect 19614 20168 19670 20224
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18602 17312 18658 17368
rect 17866 16496 17922 16552
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18510 15952 18566 16008
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 17590 13932 17646 13968
rect 17590 13912 17592 13932
rect 17592 13912 17644 13932
rect 17644 13912 17646 13932
rect 17038 9696 17094 9752
rect 16946 8608 17002 8664
rect 17682 12552 17738 12608
rect 17590 9424 17646 9480
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 9494 6160 9550 6216
rect 11886 6160 11942 6216
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 2962 992 3018 1048
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18786 17992 18842 18048
rect 18602 13932 18658 13968
rect 18602 13912 18604 13932
rect 18604 13912 18656 13932
rect 18656 13912 18658 13932
rect 19154 17040 19210 17096
rect 18878 14612 18934 14648
rect 18878 14592 18880 14612
rect 18880 14592 18932 14612
rect 18932 14592 18934 14612
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 17774 10512 17830 10568
rect 18418 12144 18474 12200
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18234 11092 18236 11112
rect 18236 11092 18288 11112
rect 18288 11092 18290 11112
rect 18234 11056 18290 11092
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18234 10512 18290 10568
rect 18142 10104 18198 10160
rect 18786 11328 18842 11384
rect 18694 11212 18750 11248
rect 18694 11192 18696 11212
rect 18696 11192 18748 11212
rect 18748 11192 18750 11212
rect 18694 10784 18750 10840
rect 18602 10668 18658 10704
rect 18602 10648 18604 10668
rect 18604 10648 18656 10668
rect 18656 10648 18658 10668
rect 17958 9988 18014 10024
rect 17958 9968 17960 9988
rect 17960 9968 18012 9988
rect 18012 9968 18014 9988
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18510 8880 18566 8936
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 17958 8472 18014 8528
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18786 9016 18842 9072
rect 18786 8880 18842 8936
rect 19062 13640 19118 13696
rect 20166 19780 20222 19816
rect 20166 19760 20168 19780
rect 20168 19760 20220 19780
rect 20220 19760 20222 19780
rect 19890 18264 19946 18320
rect 19154 13232 19210 13288
rect 20166 18808 20222 18864
rect 20442 18944 20498 19000
rect 20626 18264 20682 18320
rect 20534 17856 20590 17912
rect 19246 12824 19302 12880
rect 19062 12688 19118 12744
rect 19154 12144 19210 12200
rect 19154 11464 19210 11520
rect 18970 8064 19026 8120
rect 18878 7520 18934 7576
rect 18786 7112 18842 7168
rect 17958 6704 18014 6760
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17958 5752 18014 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18510 5208 18566 5264
rect 17958 4800 18014 4856
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 17406 2488 17462 2544
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 2870 176 2926 232
rect 18970 992 19026 1048
rect 20442 16496 20498 16552
rect 21270 18672 21326 18728
rect 20902 18128 20958 18184
rect 21822 19216 21878 19272
rect 20626 16904 20682 16960
rect 20350 15544 20406 15600
rect 20626 15000 20682 15056
rect 20442 14048 20498 14104
rect 20442 13640 20498 13696
rect 20718 12552 20774 12608
rect 19982 3440 20038 3496
rect 19154 2896 19210 2952
rect 20258 4256 20314 4312
rect 20166 3848 20222 3904
rect 20074 1536 20130 1592
rect 20718 1944 20774 2000
rect 19062 584 19118 640
rect 18878 176 18934 232
<< metal3 >>
rect 0 22538 800 22568
rect 3049 22538 3115 22541
rect 0 22536 3115 22538
rect 0 22480 3054 22536
rect 3110 22480 3115 22536
rect 0 22478 3115 22480
rect 0 22448 800 22478
rect 3049 22475 3115 22478
rect 17769 22538 17835 22541
rect 22000 22538 22800 22568
rect 17769 22536 22800 22538
rect 17769 22480 17774 22536
rect 17830 22480 22800 22536
rect 17769 22478 22800 22480
rect 17769 22475 17835 22478
rect 22000 22448 22800 22478
rect 0 22130 800 22160
rect 2773 22130 2839 22133
rect 0 22128 2839 22130
rect 0 22072 2778 22128
rect 2834 22072 2839 22128
rect 0 22070 2839 22072
rect 0 22040 800 22070
rect 2773 22067 2839 22070
rect 18505 22130 18571 22133
rect 22000 22130 22800 22160
rect 18505 22128 22800 22130
rect 18505 22072 18510 22128
rect 18566 22072 22800 22128
rect 18505 22070 22800 22072
rect 18505 22067 18571 22070
rect 22000 22040 22800 22070
rect 0 21586 800 21616
rect 2957 21586 3023 21589
rect 0 21584 3023 21586
rect 0 21528 2962 21584
rect 3018 21528 3023 21584
rect 0 21526 3023 21528
rect 0 21496 800 21526
rect 2957 21523 3023 21526
rect 18597 21586 18663 21589
rect 22000 21586 22800 21616
rect 18597 21584 22800 21586
rect 18597 21528 18602 21584
rect 18658 21528 22800 21584
rect 18597 21526 22800 21528
rect 18597 21523 18663 21526
rect 22000 21496 22800 21526
rect 0 21178 800 21208
rect 4061 21178 4127 21181
rect 0 21176 4127 21178
rect 0 21120 4066 21176
rect 4122 21120 4127 21176
rect 0 21118 4127 21120
rect 0 21088 800 21118
rect 4061 21115 4127 21118
rect 19057 21178 19123 21181
rect 22000 21178 22800 21208
rect 19057 21176 22800 21178
rect 19057 21120 19062 21176
rect 19118 21120 22800 21176
rect 19057 21118 22800 21120
rect 19057 21115 19123 21118
rect 22000 21088 22800 21118
rect 0 20634 800 20664
rect 2865 20634 2931 20637
rect 0 20632 2931 20634
rect 0 20576 2870 20632
rect 2926 20576 2931 20632
rect 0 20574 2931 20576
rect 0 20544 800 20574
rect 2865 20571 2931 20574
rect 19241 20634 19307 20637
rect 22000 20634 22800 20664
rect 19241 20632 22800 20634
rect 19241 20576 19246 20632
rect 19302 20576 22800 20632
rect 19241 20574 22800 20576
rect 19241 20571 19307 20574
rect 22000 20544 22800 20574
rect 0 20226 800 20256
rect 3509 20226 3575 20229
rect 0 20224 3575 20226
rect 0 20168 3514 20224
rect 3570 20168 3575 20224
rect 0 20166 3575 20168
rect 0 20136 800 20166
rect 3509 20163 3575 20166
rect 19609 20226 19675 20229
rect 22000 20226 22800 20256
rect 19609 20224 22800 20226
rect 19609 20168 19614 20224
rect 19670 20168 22800 20224
rect 19609 20166 22800 20168
rect 19609 20163 19675 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22000 20136 22800 20166
rect 14672 20095 14992 20096
rect 0 19818 800 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 800 19758
rect 1945 19755 2011 19758
rect 20161 19818 20227 19821
rect 22000 19818 22800 19848
rect 20161 19816 22800 19818
rect 20161 19760 20166 19816
rect 20222 19760 22800 19816
rect 20161 19758 22800 19760
rect 20161 19755 20227 19758
rect 22000 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 800 19304
rect 2037 19274 2103 19277
rect 21817 19274 21883 19277
rect 22000 19274 22800 19304
rect 0 19214 1962 19274
rect 0 19184 800 19214
rect 1902 19138 1962 19214
rect 2037 19272 21883 19274
rect 2037 19216 2042 19272
rect 2098 19216 21822 19272
rect 21878 19216 21883 19272
rect 2037 19214 21883 19216
rect 2037 19211 2103 19214
rect 21817 19211 21883 19214
rect 21958 19184 22800 19274
rect 2773 19138 2839 19141
rect 1902 19136 2839 19138
rect 1902 19080 2778 19136
rect 2834 19080 2839 19136
rect 1902 19078 2839 19080
rect 2773 19075 2839 19078
rect 17677 19138 17743 19141
rect 21958 19138 22018 19184
rect 17677 19136 22018 19138
rect 17677 19080 17682 19136
rect 17738 19080 22018 19136
rect 17677 19078 22018 19080
rect 17677 19075 17743 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 8334 18940 8340 19004
rect 8404 19002 8410 19004
rect 12893 19002 12959 19005
rect 20437 19002 20503 19005
rect 8404 19000 12959 19002
rect 8404 18944 12898 19000
rect 12954 18944 12959 19000
rect 8404 18942 12959 18944
rect 8404 18940 8410 18942
rect 12893 18939 12959 18942
rect 16438 19000 20503 19002
rect 16438 18944 20442 19000
rect 20498 18944 20503 19000
rect 16438 18942 20503 18944
rect 0 18866 800 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 800 18806
rect 1945 18803 2011 18806
rect 2589 18866 2655 18869
rect 16438 18866 16498 18942
rect 20437 18939 20503 18942
rect 2589 18864 16498 18866
rect 2589 18808 2594 18864
rect 2650 18808 16498 18864
rect 2589 18806 16498 18808
rect 20161 18866 20227 18869
rect 22000 18866 22800 18896
rect 20161 18864 22800 18866
rect 20161 18808 20166 18864
rect 20222 18808 22800 18864
rect 20161 18806 22800 18808
rect 2589 18803 2655 18806
rect 20161 18803 20227 18806
rect 22000 18776 22800 18806
rect 2129 18730 2195 18733
rect 5349 18730 5415 18733
rect 21265 18730 21331 18733
rect 2129 18728 4906 18730
rect 2129 18672 2134 18728
rect 2190 18672 4906 18728
rect 2129 18670 4906 18672
rect 2129 18667 2195 18670
rect 4846 18594 4906 18670
rect 5349 18728 21331 18730
rect 5349 18672 5354 18728
rect 5410 18672 21270 18728
rect 21326 18672 21331 18728
rect 5349 18670 21331 18672
rect 5349 18667 5415 18670
rect 21265 18667 21331 18670
rect 8845 18594 8911 18597
rect 4846 18592 8911 18594
rect 4846 18536 8850 18592
rect 8906 18536 8911 18592
rect 4846 18534 8911 18536
rect 8845 18531 8911 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 6361 18458 6427 18461
rect 9765 18458 9831 18461
rect 6361 18456 9831 18458
rect 6361 18400 6366 18456
rect 6422 18400 9770 18456
rect 9826 18400 9831 18456
rect 6361 18398 9831 18400
rect 6361 18395 6427 18398
rect 9765 18395 9831 18398
rect 0 18322 800 18352
rect 3141 18322 3207 18325
rect 0 18320 3207 18322
rect 0 18264 3146 18320
rect 3202 18264 3207 18320
rect 0 18262 3207 18264
rect 0 18232 800 18262
rect 3141 18259 3207 18262
rect 3969 18322 4035 18325
rect 19885 18322 19951 18325
rect 3969 18320 19951 18322
rect 3969 18264 3974 18320
rect 4030 18264 19890 18320
rect 19946 18264 19951 18320
rect 3969 18262 19951 18264
rect 3969 18259 4035 18262
rect 19885 18259 19951 18262
rect 20621 18322 20687 18325
rect 22000 18322 22800 18352
rect 20621 18320 22800 18322
rect 20621 18264 20626 18320
rect 20682 18264 22800 18320
rect 20621 18262 22800 18264
rect 20621 18259 20687 18262
rect 22000 18232 22800 18262
rect 3601 18186 3667 18189
rect 20897 18186 20963 18189
rect 3601 18184 20963 18186
rect 3601 18128 3606 18184
rect 3662 18128 20902 18184
rect 20958 18128 20963 18184
rect 3601 18126 20963 18128
rect 3601 18123 3667 18126
rect 20897 18123 20963 18126
rect 12985 18052 13051 18053
rect 12934 17988 12940 18052
rect 13004 18050 13051 18052
rect 17953 18050 18019 18053
rect 18781 18050 18847 18053
rect 13004 18048 13096 18050
rect 13046 17992 13096 18048
rect 13004 17990 13096 17992
rect 17953 18048 18847 18050
rect 17953 17992 17958 18048
rect 18014 17992 18786 18048
rect 18842 17992 18847 18048
rect 17953 17990 18847 17992
rect 13004 17988 13051 17990
rect 12985 17987 13051 17988
rect 17953 17987 18019 17990
rect 18781 17987 18847 17990
rect 7808 17984 8128 17985
rect 0 17914 800 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 3049 17914 3115 17917
rect 0 17912 3115 17914
rect 0 17856 3054 17912
rect 3110 17856 3115 17912
rect 0 17854 3115 17856
rect 0 17824 800 17854
rect 3049 17851 3115 17854
rect 20529 17914 20595 17917
rect 22000 17914 22800 17944
rect 20529 17912 22800 17914
rect 20529 17856 20534 17912
rect 20590 17856 22800 17912
rect 20529 17854 22800 17856
rect 20529 17851 20595 17854
rect 22000 17824 22800 17854
rect 6821 17778 6887 17781
rect 10133 17778 10199 17781
rect 6821 17776 10199 17778
rect 6821 17720 6826 17776
rect 6882 17720 10138 17776
rect 10194 17720 10199 17776
rect 6821 17718 10199 17720
rect 6821 17715 6887 17718
rect 10133 17715 10199 17718
rect 2129 17642 2195 17645
rect 9581 17642 9647 17645
rect 2129 17640 9647 17642
rect 2129 17584 2134 17640
rect 2190 17584 9586 17640
rect 9642 17584 9647 17640
rect 2129 17582 9647 17584
rect 2129 17579 2195 17582
rect 9581 17579 9647 17582
rect 10225 17642 10291 17645
rect 13445 17642 13511 17645
rect 10225 17640 13511 17642
rect 10225 17584 10230 17640
rect 10286 17584 13450 17640
rect 13506 17584 13511 17640
rect 10225 17582 13511 17584
rect 10225 17579 10291 17582
rect 13445 17579 13511 17582
rect 5165 17506 5231 17509
rect 8334 17506 8340 17508
rect 5165 17504 8340 17506
rect 5165 17448 5170 17504
rect 5226 17448 8340 17504
rect 5165 17446 8340 17448
rect 5165 17443 5231 17446
rect 8334 17444 8340 17446
rect 8404 17444 8410 17508
rect 4376 17440 4696 17441
rect 0 17370 800 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 2773 17370 2839 17373
rect 0 17368 2839 17370
rect 0 17312 2778 17368
rect 2834 17312 2839 17368
rect 0 17310 2839 17312
rect 0 17280 800 17310
rect 2773 17307 2839 17310
rect 18597 17370 18663 17373
rect 22000 17370 22800 17400
rect 18597 17368 22800 17370
rect 18597 17312 18602 17368
rect 18658 17312 22800 17368
rect 18597 17310 22800 17312
rect 18597 17307 18663 17310
rect 22000 17280 22800 17310
rect 8017 17234 8083 17237
rect 11237 17234 11303 17237
rect 8017 17232 11303 17234
rect 8017 17176 8022 17232
rect 8078 17176 11242 17232
rect 11298 17176 11303 17232
rect 8017 17174 11303 17176
rect 8017 17171 8083 17174
rect 11237 17171 11303 17174
rect 6453 17098 6519 17101
rect 9581 17098 9647 17101
rect 6453 17096 9647 17098
rect 6453 17040 6458 17096
rect 6514 17040 9586 17096
rect 9642 17040 9647 17096
rect 6453 17038 9647 17040
rect 6453 17035 6519 17038
rect 9581 17035 9647 17038
rect 19149 17100 19215 17101
rect 19149 17096 19196 17100
rect 19260 17098 19266 17100
rect 19149 17040 19154 17096
rect 19149 17036 19196 17040
rect 19260 17038 19306 17098
rect 19260 17036 19266 17038
rect 19149 17035 19215 17036
rect 0 16962 800 16992
rect 1945 16962 2011 16965
rect 0 16960 2011 16962
rect 0 16904 1950 16960
rect 2006 16904 2011 16960
rect 0 16902 2011 16904
rect 0 16872 800 16902
rect 1945 16899 2011 16902
rect 3233 16962 3299 16965
rect 6545 16962 6611 16965
rect 3233 16960 6611 16962
rect 3233 16904 3238 16960
rect 3294 16904 6550 16960
rect 6606 16904 6611 16960
rect 3233 16902 6611 16904
rect 3233 16899 3299 16902
rect 6545 16899 6611 16902
rect 20621 16962 20687 16965
rect 22000 16962 22800 16992
rect 20621 16960 22800 16962
rect 20621 16904 20626 16960
rect 20682 16904 22800 16960
rect 20621 16902 22800 16904
rect 20621 16899 20687 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22000 16872 22800 16902
rect 14672 16831 14992 16832
rect 5441 16690 5507 16693
rect 11237 16690 11303 16693
rect 5441 16688 11303 16690
rect 5441 16632 5446 16688
rect 5502 16632 11242 16688
rect 11298 16632 11303 16688
rect 5441 16630 11303 16632
rect 5441 16627 5507 16630
rect 11237 16627 11303 16630
rect 0 16554 800 16584
rect 1945 16554 2011 16557
rect 0 16552 2011 16554
rect 0 16496 1950 16552
rect 2006 16496 2011 16552
rect 0 16494 2011 16496
rect 0 16464 800 16494
rect 1945 16491 2011 16494
rect 10225 16554 10291 16557
rect 17861 16554 17927 16557
rect 10225 16552 17927 16554
rect 10225 16496 10230 16552
rect 10286 16496 17866 16552
rect 17922 16496 17927 16552
rect 10225 16494 17927 16496
rect 10225 16491 10291 16494
rect 17861 16491 17927 16494
rect 20437 16554 20503 16557
rect 22000 16554 22800 16584
rect 20437 16552 22800 16554
rect 20437 16496 20442 16552
rect 20498 16496 22800 16552
rect 20437 16494 22800 16496
rect 20437 16491 20503 16494
rect 22000 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 10317 16146 10383 16149
rect 15193 16146 15259 16149
rect 10317 16144 15259 16146
rect 10317 16088 10322 16144
rect 10378 16088 15198 16144
rect 15254 16088 15259 16144
rect 10317 16086 15259 16088
rect 10317 16083 10383 16086
rect 15193 16083 15259 16086
rect 0 16010 800 16040
rect 2497 16010 2563 16013
rect 0 16008 2563 16010
rect 0 15952 2502 16008
rect 2558 15952 2563 16008
rect 0 15950 2563 15952
rect 0 15920 800 15950
rect 2497 15947 2563 15950
rect 5533 16010 5599 16013
rect 9305 16010 9371 16013
rect 5533 16008 9371 16010
rect 5533 15952 5538 16008
rect 5594 15952 9310 16008
rect 9366 15952 9371 16008
rect 5533 15950 9371 15952
rect 5533 15947 5599 15950
rect 9305 15947 9371 15950
rect 10961 16010 11027 16013
rect 17493 16010 17559 16013
rect 10961 16008 17559 16010
rect 10961 15952 10966 16008
rect 11022 15952 17498 16008
rect 17554 15952 17559 16008
rect 10961 15950 17559 15952
rect 10961 15947 11027 15950
rect 17493 15947 17559 15950
rect 18505 16010 18571 16013
rect 22000 16010 22800 16040
rect 18505 16008 22800 16010
rect 18505 15952 18510 16008
rect 18566 15952 22800 16008
rect 18505 15950 22800 15952
rect 18505 15947 18571 15950
rect 22000 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 4981 15738 5047 15741
rect 11881 15738 11947 15741
rect 13997 15738 14063 15741
rect 4981 15736 5090 15738
rect 4981 15680 4986 15736
rect 5042 15680 5090 15736
rect 4981 15675 5090 15680
rect 11881 15736 14063 15738
rect 11881 15680 11886 15736
rect 11942 15680 14002 15736
rect 14058 15680 14063 15736
rect 11881 15678 14063 15680
rect 11881 15675 11947 15678
rect 13997 15675 14063 15678
rect 0 15602 800 15632
rect 1945 15602 2011 15605
rect 0 15600 2011 15602
rect 0 15544 1950 15600
rect 2006 15544 2011 15600
rect 0 15542 2011 15544
rect 0 15512 800 15542
rect 1945 15539 2011 15542
rect 5030 15466 5090 15675
rect 20345 15602 20411 15605
rect 22000 15602 22800 15632
rect 20345 15600 22800 15602
rect 20345 15544 20350 15600
rect 20406 15544 22800 15600
rect 20345 15542 22800 15544
rect 20345 15539 20411 15542
rect 22000 15512 22800 15542
rect 5165 15466 5231 15469
rect 5030 15464 5231 15466
rect 5030 15408 5170 15464
rect 5226 15408 5231 15464
rect 5030 15406 5231 15408
rect 5165 15403 5231 15406
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 11881 15194 11947 15197
rect 12249 15194 12315 15197
rect 13813 15194 13879 15197
rect 11881 15192 13879 15194
rect 11881 15136 11886 15192
rect 11942 15136 12254 15192
rect 12310 15136 13818 15192
rect 13874 15136 13879 15192
rect 11881 15134 13879 15136
rect 11881 15131 11947 15134
rect 12249 15131 12315 15134
rect 13813 15131 13879 15134
rect 0 15058 800 15088
rect 1945 15058 2011 15061
rect 0 15056 2011 15058
rect 0 15000 1950 15056
rect 2006 15000 2011 15056
rect 0 14998 2011 15000
rect 0 14968 800 14998
rect 1945 14995 2011 14998
rect 9673 15058 9739 15061
rect 12525 15058 12591 15061
rect 9673 15056 12591 15058
rect 9673 15000 9678 15056
rect 9734 15000 12530 15056
rect 12586 15000 12591 15056
rect 9673 14998 12591 15000
rect 9673 14995 9739 14998
rect 12525 14995 12591 14998
rect 20621 15058 20687 15061
rect 22000 15058 22800 15088
rect 20621 15056 22800 15058
rect 20621 15000 20626 15056
rect 20682 15000 22800 15056
rect 20621 14998 22800 15000
rect 20621 14995 20687 14998
rect 22000 14968 22800 14998
rect 1761 14922 1827 14925
rect 6361 14922 6427 14925
rect 9029 14922 9095 14925
rect 1761 14920 9095 14922
rect 1761 14864 1766 14920
rect 1822 14864 6366 14920
rect 6422 14864 9034 14920
rect 9090 14864 9095 14920
rect 1761 14862 9095 14864
rect 1761 14859 1827 14862
rect 6361 14859 6427 14862
rect 9029 14859 9095 14862
rect 11513 14786 11579 14789
rect 12985 14786 13051 14789
rect 11513 14784 13051 14786
rect 11513 14728 11518 14784
rect 11574 14728 12990 14784
rect 13046 14728 13051 14784
rect 11513 14726 13051 14728
rect 11513 14723 11579 14726
rect 12985 14723 13051 14726
rect 7808 14720 8128 14721
rect 0 14650 800 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 2865 14650 2931 14653
rect 0 14648 2931 14650
rect 0 14592 2870 14648
rect 2926 14592 2931 14648
rect 0 14590 2931 14592
rect 0 14560 800 14590
rect 2865 14587 2931 14590
rect 18873 14650 18939 14653
rect 22000 14650 22800 14680
rect 18873 14648 22800 14650
rect 18873 14592 18878 14648
rect 18934 14592 22800 14648
rect 18873 14590 22800 14592
rect 18873 14587 18939 14590
rect 22000 14560 22800 14590
rect 4376 14176 4696 14177
rect 0 14106 800 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1853 14106 1919 14109
rect 17401 14106 17467 14109
rect 0 14104 1919 14106
rect 0 14048 1858 14104
rect 1914 14048 1919 14104
rect 0 14046 1919 14048
rect 0 14016 800 14046
rect 1853 14043 1919 14046
rect 17358 14104 17467 14106
rect 17358 14048 17406 14104
rect 17462 14048 17467 14104
rect 17358 14043 17467 14048
rect 20437 14106 20503 14109
rect 22000 14106 22800 14136
rect 20437 14104 22800 14106
rect 20437 14048 20442 14104
rect 20498 14048 22800 14104
rect 20437 14046 22800 14048
rect 20437 14043 20503 14046
rect 17217 13834 17283 13837
rect 17358 13834 17418 14043
rect 22000 14016 22800 14046
rect 17585 13970 17651 13973
rect 18597 13970 18663 13973
rect 17585 13968 18663 13970
rect 17585 13912 17590 13968
rect 17646 13912 18602 13968
rect 18658 13912 18663 13968
rect 17585 13910 18663 13912
rect 17585 13907 17651 13910
rect 18597 13907 18663 13910
rect 17217 13832 17418 13834
rect 17217 13776 17222 13832
rect 17278 13776 17418 13832
rect 17217 13774 17418 13776
rect 17217 13771 17283 13774
rect 0 13698 800 13728
rect 2865 13698 2931 13701
rect 0 13696 2931 13698
rect 0 13640 2870 13696
rect 2926 13640 2931 13696
rect 0 13638 2931 13640
rect 0 13608 800 13638
rect 2865 13635 2931 13638
rect 15285 13698 15351 13701
rect 19057 13698 19123 13701
rect 15285 13696 19123 13698
rect 15285 13640 15290 13696
rect 15346 13640 19062 13696
rect 19118 13640 19123 13696
rect 15285 13638 19123 13640
rect 15285 13635 15351 13638
rect 19057 13635 19123 13638
rect 20437 13698 20503 13701
rect 22000 13698 22800 13728
rect 20437 13696 22800 13698
rect 20437 13640 20442 13696
rect 20498 13640 22800 13696
rect 20437 13638 22800 13640
rect 20437 13635 20503 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22000 13608 22800 13638
rect 14672 13567 14992 13568
rect 0 13290 800 13320
rect 3049 13290 3115 13293
rect 0 13288 3115 13290
rect 0 13232 3054 13288
rect 3110 13232 3115 13288
rect 0 13230 3115 13232
rect 0 13200 800 13230
rect 3049 13227 3115 13230
rect 6913 13290 6979 13293
rect 8109 13290 8175 13293
rect 6913 13288 8175 13290
rect 6913 13232 6918 13288
rect 6974 13232 8114 13288
rect 8170 13232 8175 13288
rect 6913 13230 8175 13232
rect 6913 13227 6979 13230
rect 8109 13227 8175 13230
rect 19149 13290 19215 13293
rect 22000 13290 22800 13320
rect 19149 13288 22800 13290
rect 19149 13232 19154 13288
rect 19210 13232 22800 13288
rect 19149 13230 22800 13232
rect 19149 13227 19215 13230
rect 22000 13200 22800 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 19241 12882 19307 12885
rect 16070 12880 19307 12882
rect 16070 12824 19246 12880
rect 19302 12824 19307 12880
rect 16070 12822 19307 12824
rect 0 12746 800 12776
rect 9581 12746 9647 12749
rect 0 12744 9647 12746
rect 0 12688 9586 12744
rect 9642 12688 9647 12744
rect 0 12686 9647 12688
rect 0 12656 800 12686
rect 9581 12683 9647 12686
rect 13261 12610 13327 12613
rect 13721 12610 13787 12613
rect 13261 12608 13787 12610
rect 13261 12552 13266 12608
rect 13322 12552 13726 12608
rect 13782 12552 13787 12608
rect 13261 12550 13787 12552
rect 13261 12547 13327 12550
rect 13721 12547 13787 12550
rect 15469 12610 15535 12613
rect 16070 12610 16130 12822
rect 19241 12819 19307 12822
rect 19057 12746 19123 12749
rect 22000 12746 22800 12776
rect 19057 12744 22800 12746
rect 19057 12688 19062 12744
rect 19118 12688 22800 12744
rect 19057 12686 22800 12688
rect 19057 12683 19123 12686
rect 22000 12656 22800 12686
rect 15469 12608 16130 12610
rect 15469 12552 15474 12608
rect 15530 12552 16130 12608
rect 15469 12550 16130 12552
rect 17677 12610 17743 12613
rect 19190 12610 19196 12612
rect 17677 12608 19196 12610
rect 17677 12552 17682 12608
rect 17738 12552 19196 12608
rect 17677 12550 19196 12552
rect 15469 12547 15535 12550
rect 17677 12547 17743 12550
rect 19190 12548 19196 12550
rect 19260 12610 19266 12612
rect 20713 12610 20779 12613
rect 19260 12608 20779 12610
rect 19260 12552 20718 12608
rect 20774 12552 20779 12608
rect 19260 12550 20779 12552
rect 19260 12548 19266 12550
rect 20713 12547 20779 12550
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 800 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 800 12278
rect 4061 12275 4127 12278
rect 10225 12338 10291 12341
rect 16849 12338 16915 12341
rect 22000 12338 22800 12368
rect 10225 12336 22800 12338
rect 10225 12280 10230 12336
rect 10286 12280 16854 12336
rect 16910 12280 22800 12336
rect 10225 12278 22800 12280
rect 10225 12275 10291 12278
rect 16849 12275 16915 12278
rect 22000 12248 22800 12278
rect 18413 12202 18479 12205
rect 19149 12202 19215 12205
rect 18413 12200 19215 12202
rect 18413 12144 18418 12200
rect 18474 12144 19154 12200
rect 19210 12144 19215 12200
rect 18413 12142 19215 12144
rect 18413 12139 18479 12142
rect 19149 12139 19215 12142
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 800 11824
rect 4061 11794 4127 11797
rect 0 11792 4127 11794
rect 0 11736 4066 11792
rect 4122 11736 4127 11792
rect 0 11734 4127 11736
rect 0 11704 800 11734
rect 4061 11731 4127 11734
rect 5073 11794 5139 11797
rect 5901 11794 5967 11797
rect 5073 11792 5967 11794
rect 5073 11736 5078 11792
rect 5134 11736 5906 11792
rect 5962 11736 5967 11792
rect 5073 11734 5967 11736
rect 5073 11731 5139 11734
rect 5901 11731 5967 11734
rect 15561 11794 15627 11797
rect 22000 11794 22800 11824
rect 15561 11792 22800 11794
rect 15561 11736 15566 11792
rect 15622 11736 22800 11792
rect 15561 11734 22800 11736
rect 15561 11731 15627 11734
rect 22000 11704 22800 11734
rect 11513 11658 11579 11661
rect 15193 11658 15259 11661
rect 11513 11656 15259 11658
rect 11513 11600 11518 11656
rect 11574 11600 15198 11656
rect 15254 11600 15259 11656
rect 11513 11598 15259 11600
rect 11513 11595 11579 11598
rect 15193 11595 15259 11598
rect 5206 11460 5212 11524
rect 5276 11522 5282 11524
rect 5349 11522 5415 11525
rect 5276 11520 5415 11522
rect 5276 11464 5354 11520
rect 5410 11464 5415 11520
rect 5276 11462 5415 11464
rect 5276 11460 5282 11462
rect 5349 11459 5415 11462
rect 16665 11522 16731 11525
rect 19149 11522 19215 11525
rect 16665 11520 19215 11522
rect 16665 11464 16670 11520
rect 16726 11464 19154 11520
rect 19210 11464 19215 11520
rect 16665 11462 19215 11464
rect 16665 11459 16731 11462
rect 19149 11459 19215 11462
rect 7808 11456 8128 11457
rect 0 11386 800 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 3785 11386 3851 11389
rect 0 11384 3851 11386
rect 0 11328 3790 11384
rect 3846 11328 3851 11384
rect 0 11326 3851 11328
rect 0 11296 800 11326
rect 3785 11323 3851 11326
rect 18781 11386 18847 11389
rect 22000 11386 22800 11416
rect 18781 11384 22800 11386
rect 18781 11328 18786 11384
rect 18842 11328 22800 11384
rect 18781 11326 22800 11328
rect 18781 11323 18847 11326
rect 22000 11296 22800 11326
rect 16297 11250 16363 11253
rect 18689 11250 18755 11253
rect 16297 11248 18755 11250
rect 16297 11192 16302 11248
rect 16358 11192 18694 11248
rect 18750 11192 18755 11248
rect 16297 11190 18755 11192
rect 16297 11187 16363 11190
rect 18689 11187 18755 11190
rect 11329 11114 11395 11117
rect 13261 11114 13327 11117
rect 11329 11112 13327 11114
rect 11329 11056 11334 11112
rect 11390 11056 13266 11112
rect 13322 11056 13327 11112
rect 11329 11054 13327 11056
rect 11329 11051 11395 11054
rect 13261 11051 13327 11054
rect 16021 11114 16087 11117
rect 18229 11114 18295 11117
rect 16021 11112 18295 11114
rect 16021 11056 16026 11112
rect 16082 11056 18234 11112
rect 18290 11056 18295 11112
rect 16021 11054 18295 11056
rect 16021 11051 16087 11054
rect 18229 11051 18295 11054
rect 4376 10912 4696 10913
rect 0 10842 800 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 0 10752 800 10782
rect 4061 10779 4127 10782
rect 18689 10842 18755 10845
rect 22000 10842 22800 10872
rect 18689 10840 22800 10842
rect 18689 10784 18694 10840
rect 18750 10784 22800 10840
rect 18689 10782 22800 10784
rect 18689 10779 18755 10782
rect 22000 10752 22800 10782
rect 15009 10706 15075 10709
rect 18597 10706 18663 10709
rect 15009 10704 18663 10706
rect 15009 10648 15014 10704
rect 15070 10648 18602 10704
rect 18658 10648 18663 10704
rect 15009 10646 18663 10648
rect 15009 10643 15075 10646
rect 18597 10643 18663 10646
rect 10593 10570 10659 10573
rect 12934 10570 12940 10572
rect 10593 10568 12940 10570
rect 10593 10512 10598 10568
rect 10654 10512 12940 10568
rect 10593 10510 12940 10512
rect 10593 10507 10659 10510
rect 12934 10508 12940 10510
rect 13004 10570 13010 10572
rect 17769 10570 17835 10573
rect 18229 10570 18295 10573
rect 13004 10568 18295 10570
rect 13004 10512 17774 10568
rect 17830 10512 18234 10568
rect 18290 10512 18295 10568
rect 13004 10510 18295 10512
rect 13004 10508 13010 10510
rect 17769 10507 17835 10510
rect 18229 10507 18295 10510
rect 0 10434 800 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 800 10374
rect 4061 10371 4127 10374
rect 15377 10434 15443 10437
rect 22000 10434 22800 10464
rect 15377 10432 22800 10434
rect 15377 10376 15382 10432
rect 15438 10376 22800 10432
rect 15377 10374 22800 10376
rect 15377 10371 15443 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22000 10344 22800 10374
rect 14672 10303 14992 10304
rect 9213 10162 9279 10165
rect 6318 10160 9279 10162
rect 6318 10104 9218 10160
rect 9274 10104 9279 10160
rect 6318 10102 9279 10104
rect 0 10026 800 10056
rect 6318 10026 6378 10102
rect 9213 10099 9279 10102
rect 12249 10162 12315 10165
rect 18137 10162 18203 10165
rect 12249 10160 18203 10162
rect 12249 10104 12254 10160
rect 12310 10104 18142 10160
rect 18198 10104 18203 10160
rect 12249 10102 18203 10104
rect 12249 10099 12315 10102
rect 18137 10099 18203 10102
rect 0 9966 6378 10026
rect 6453 10026 6519 10029
rect 15377 10026 15443 10029
rect 6453 10024 15443 10026
rect 6453 9968 6458 10024
rect 6514 9968 15382 10024
rect 15438 9968 15443 10024
rect 6453 9966 15443 9968
rect 0 9936 800 9966
rect 6453 9963 6519 9966
rect 15377 9963 15443 9966
rect 17953 10026 18019 10029
rect 22000 10026 22800 10056
rect 17953 10024 22800 10026
rect 17953 9968 17958 10024
rect 18014 9968 22800 10024
rect 17953 9966 22800 9968
rect 17953 9963 18019 9966
rect 22000 9936 22800 9966
rect 12157 9890 12223 9893
rect 12433 9890 12499 9893
rect 12157 9888 12499 9890
rect 12157 9832 12162 9888
rect 12218 9832 12438 9888
rect 12494 9832 12499 9888
rect 12157 9830 12499 9832
rect 12157 9827 12223 9830
rect 12433 9827 12499 9830
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 8334 9754 8340 9756
rect 5950 9694 8340 9754
rect 5950 9621 6010 9694
rect 8334 9692 8340 9694
rect 8404 9692 8410 9756
rect 11881 9754 11947 9757
rect 17033 9754 17099 9757
rect 11881 9752 17099 9754
rect 11881 9696 11886 9752
rect 11942 9696 17038 9752
rect 17094 9696 17099 9752
rect 11881 9694 17099 9696
rect 11881 9691 11947 9694
rect 17033 9691 17099 9694
rect 5950 9616 6059 9621
rect 5950 9560 5998 9616
rect 6054 9560 6059 9616
rect 5950 9558 6059 9560
rect 5993 9555 6059 9558
rect 8845 9618 8911 9621
rect 9489 9618 9555 9621
rect 8845 9616 9555 9618
rect 8845 9560 8850 9616
rect 8906 9560 9494 9616
rect 9550 9560 9555 9616
rect 8845 9558 9555 9560
rect 8845 9555 8911 9558
rect 9489 9555 9555 9558
rect 10501 9618 10567 9621
rect 15009 9618 15075 9621
rect 10501 9616 15075 9618
rect 10501 9560 10506 9616
rect 10562 9560 15014 9616
rect 15070 9560 15075 9616
rect 10501 9558 15075 9560
rect 10501 9555 10567 9558
rect 15009 9555 15075 9558
rect 0 9482 800 9512
rect 3969 9482 4035 9485
rect 0 9480 4035 9482
rect 0 9424 3974 9480
rect 4030 9424 4035 9480
rect 0 9422 4035 9424
rect 0 9392 800 9422
rect 3969 9419 4035 9422
rect 17585 9482 17651 9485
rect 22000 9482 22800 9512
rect 17585 9480 22800 9482
rect 17585 9424 17590 9480
rect 17646 9424 22800 9480
rect 17585 9422 22800 9424
rect 17585 9419 17651 9422
rect 22000 9392 22800 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 800 9104
rect 5993 9074 6059 9077
rect 0 9072 6059 9074
rect 0 9016 5998 9072
rect 6054 9016 6059 9072
rect 0 9014 6059 9016
rect 0 8984 800 9014
rect 5993 9011 6059 9014
rect 18781 9074 18847 9077
rect 22000 9074 22800 9104
rect 18781 9072 22800 9074
rect 18781 9016 18786 9072
rect 18842 9016 22800 9072
rect 18781 9014 22800 9016
rect 18781 9011 18847 9014
rect 22000 8984 22800 9014
rect 18505 8938 18571 8941
rect 18781 8938 18847 8941
rect 18505 8936 18847 8938
rect 18505 8880 18510 8936
rect 18566 8880 18786 8936
rect 18842 8880 18847 8936
rect 18505 8878 18847 8880
rect 18505 8875 18571 8878
rect 18781 8875 18847 8878
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 11973 8666 12039 8669
rect 16941 8666 17007 8669
rect 11973 8664 17007 8666
rect 11973 8608 11978 8664
rect 12034 8608 16946 8664
rect 17002 8608 17007 8664
rect 11973 8606 17007 8608
rect 11973 8603 12039 8606
rect 16941 8603 17007 8606
rect 0 8530 800 8560
rect 4061 8530 4127 8533
rect 0 8528 4127 8530
rect 0 8472 4066 8528
rect 4122 8472 4127 8528
rect 0 8470 4127 8472
rect 0 8440 800 8470
rect 4061 8467 4127 8470
rect 9581 8530 9647 8533
rect 12617 8530 12683 8533
rect 9581 8528 12683 8530
rect 9581 8472 9586 8528
rect 9642 8472 12622 8528
rect 12678 8472 12683 8528
rect 9581 8470 12683 8472
rect 9581 8467 9647 8470
rect 12617 8467 12683 8470
rect 17953 8530 18019 8533
rect 22000 8530 22800 8560
rect 17953 8528 22800 8530
rect 17953 8472 17958 8528
rect 18014 8472 22800 8528
rect 17953 8470 22800 8472
rect 17953 8467 18019 8470
rect 22000 8440 22800 8470
rect 4613 8394 4679 8397
rect 6453 8394 6519 8397
rect 4613 8392 6519 8394
rect 4613 8336 4618 8392
rect 4674 8336 6458 8392
rect 6514 8336 6519 8392
rect 4613 8334 6519 8336
rect 4613 8331 4679 8334
rect 6453 8331 6519 8334
rect 7808 8192 8128 8193
rect 0 8122 800 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 800 8062
rect 4061 8059 4127 8062
rect 18965 8122 19031 8125
rect 22000 8122 22800 8152
rect 18965 8120 22800 8122
rect 18965 8064 18970 8120
rect 19026 8064 22800 8120
rect 18965 8062 22800 8064
rect 18965 8059 19031 8062
rect 22000 8032 22800 8062
rect 4376 7648 4696 7649
rect 0 7578 800 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 2681 7578 2747 7581
rect 0 7576 2747 7578
rect 0 7520 2686 7576
rect 2742 7520 2747 7576
rect 0 7518 2747 7520
rect 0 7488 800 7518
rect 2681 7515 2747 7518
rect 18873 7578 18939 7581
rect 22000 7578 22800 7608
rect 18873 7576 22800 7578
rect 18873 7520 18878 7576
rect 18934 7520 22800 7576
rect 18873 7518 22800 7520
rect 18873 7515 18939 7518
rect 22000 7488 22800 7518
rect 0 7170 800 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 800 7110
rect 4061 7107 4127 7110
rect 18781 7170 18847 7173
rect 22000 7170 22800 7200
rect 18781 7168 22800 7170
rect 18781 7112 18786 7168
rect 18842 7112 22800 7168
rect 18781 7110 22800 7112
rect 18781 7107 18847 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22000 7080 22800 7110
rect 14672 7039 14992 7040
rect 0 6762 800 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 800 6702
rect 4061 6699 4127 6702
rect 17953 6762 18019 6765
rect 22000 6762 22800 6792
rect 17953 6760 22800 6762
rect 17953 6704 17958 6760
rect 18014 6704 22800 6760
rect 17953 6702 22800 6704
rect 17953 6699 18019 6702
rect 22000 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6218 800 6248
rect 4797 6218 4863 6221
rect 0 6216 4863 6218
rect 0 6160 4802 6216
rect 4858 6160 4863 6216
rect 0 6158 4863 6160
rect 0 6128 800 6158
rect 4797 6155 4863 6158
rect 5206 6156 5212 6220
rect 5276 6218 5282 6220
rect 9489 6218 9555 6221
rect 5276 6216 9555 6218
rect 5276 6160 9494 6216
rect 9550 6160 9555 6216
rect 5276 6158 9555 6160
rect 5276 6156 5282 6158
rect 9489 6155 9555 6158
rect 11881 6218 11947 6221
rect 22000 6218 22800 6248
rect 11881 6216 22800 6218
rect 11881 6160 11886 6216
rect 11942 6160 22800 6216
rect 11881 6158 22800 6160
rect 11881 6155 11947 6158
rect 22000 6128 22800 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 800 5840
rect 3417 5810 3483 5813
rect 0 5808 3483 5810
rect 0 5752 3422 5808
rect 3478 5752 3483 5808
rect 0 5750 3483 5752
rect 0 5720 800 5750
rect 3417 5747 3483 5750
rect 17953 5810 18019 5813
rect 22000 5810 22800 5840
rect 17953 5808 22800 5810
rect 17953 5752 17958 5808
rect 18014 5752 22800 5808
rect 17953 5750 22800 5752
rect 17953 5747 18019 5750
rect 22000 5720 22800 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 800 5296
rect 3969 5266 4035 5269
rect 0 5264 4035 5266
rect 0 5208 3974 5264
rect 4030 5208 4035 5264
rect 0 5206 4035 5208
rect 0 5176 800 5206
rect 3969 5203 4035 5206
rect 18505 5266 18571 5269
rect 22000 5266 22800 5296
rect 18505 5264 22800 5266
rect 18505 5208 18510 5264
rect 18566 5208 22800 5264
rect 18505 5206 22800 5208
rect 18505 5203 18571 5206
rect 22000 5176 22800 5206
rect 7808 4928 8128 4929
rect 0 4858 800 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 800 4798
rect 4061 4795 4127 4798
rect 17953 4858 18019 4861
rect 22000 4858 22800 4888
rect 17953 4856 22800 4858
rect 17953 4800 17958 4856
rect 18014 4800 22800 4856
rect 17953 4798 22800 4800
rect 17953 4795 18019 4798
rect 22000 4768 22800 4798
rect 4376 4384 4696 4385
rect 0 4314 800 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 1117 4314 1183 4317
rect 0 4312 1183 4314
rect 0 4256 1122 4312
rect 1178 4256 1183 4312
rect 0 4254 1183 4256
rect 0 4224 800 4254
rect 1117 4251 1183 4254
rect 20253 4314 20319 4317
rect 22000 4314 22800 4344
rect 20253 4312 22800 4314
rect 20253 4256 20258 4312
rect 20314 4256 22800 4312
rect 20253 4254 22800 4256
rect 20253 4251 20319 4254
rect 22000 4224 22800 4254
rect 0 3906 800 3936
rect 4705 3906 4771 3909
rect 0 3904 4771 3906
rect 0 3848 4710 3904
rect 4766 3848 4771 3904
rect 0 3846 4771 3848
rect 0 3816 800 3846
rect 4705 3843 4771 3846
rect 20161 3906 20227 3909
rect 22000 3906 22800 3936
rect 20161 3904 22800 3906
rect 20161 3848 20166 3904
rect 20222 3848 22800 3904
rect 20161 3846 22800 3848
rect 20161 3843 20227 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22000 3816 22800 3846
rect 14672 3775 14992 3776
rect 0 3498 800 3528
rect 3233 3498 3299 3501
rect 0 3496 3299 3498
rect 0 3440 3238 3496
rect 3294 3440 3299 3496
rect 0 3438 3299 3440
rect 0 3408 800 3438
rect 3233 3435 3299 3438
rect 19977 3498 20043 3501
rect 22000 3498 22800 3528
rect 19977 3496 22800 3498
rect 19977 3440 19982 3496
rect 20038 3440 22800 3496
rect 19977 3438 22800 3440
rect 19977 3435 20043 3438
rect 22000 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 800 2984
rect 4981 2954 5047 2957
rect 0 2952 5047 2954
rect 0 2896 4986 2952
rect 5042 2896 5047 2952
rect 0 2894 5047 2896
rect 0 2864 800 2894
rect 4981 2891 5047 2894
rect 19149 2954 19215 2957
rect 22000 2954 22800 2984
rect 19149 2952 22800 2954
rect 19149 2896 19154 2952
rect 19210 2896 22800 2952
rect 19149 2894 22800 2896
rect 19149 2891 19215 2894
rect 22000 2864 22800 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 800 2576
rect 2865 2546 2931 2549
rect 0 2544 2931 2546
rect 0 2488 2870 2544
rect 2926 2488 2931 2544
rect 0 2486 2931 2488
rect 0 2456 800 2486
rect 2865 2483 2931 2486
rect 17401 2546 17467 2549
rect 22000 2546 22800 2576
rect 17401 2544 22800 2546
rect 17401 2488 17406 2544
rect 17462 2488 22800 2544
rect 17401 2486 22800 2488
rect 17401 2483 17467 2486
rect 22000 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 800 2032
rect 5165 2002 5231 2005
rect 0 2000 5231 2002
rect 0 1944 5170 2000
rect 5226 1944 5231 2000
rect 0 1942 5231 1944
rect 0 1912 800 1942
rect 5165 1939 5231 1942
rect 20713 2002 20779 2005
rect 22000 2002 22800 2032
rect 20713 2000 22800 2002
rect 20713 1944 20718 2000
rect 20774 1944 22800 2000
rect 20713 1942 22800 1944
rect 20713 1939 20779 1942
rect 22000 1912 22800 1942
rect 0 1594 800 1624
rect 4061 1594 4127 1597
rect 0 1592 4127 1594
rect 0 1536 4066 1592
rect 4122 1536 4127 1592
rect 0 1534 4127 1536
rect 0 1504 800 1534
rect 4061 1531 4127 1534
rect 20069 1594 20135 1597
rect 22000 1594 22800 1624
rect 20069 1592 22800 1594
rect 20069 1536 20074 1592
rect 20130 1536 22800 1592
rect 20069 1534 22800 1536
rect 20069 1531 20135 1534
rect 22000 1504 22800 1534
rect 0 1050 800 1080
rect 2957 1050 3023 1053
rect 0 1048 3023 1050
rect 0 992 2962 1048
rect 3018 992 3023 1048
rect 0 990 3023 992
rect 0 960 800 990
rect 2957 987 3023 990
rect 18965 1050 19031 1053
rect 22000 1050 22800 1080
rect 18965 1048 22800 1050
rect 18965 992 18970 1048
rect 19026 992 22800 1048
rect 18965 990 22800 992
rect 18965 987 19031 990
rect 22000 960 22800 990
rect 0 642 800 672
rect 2497 642 2563 645
rect 0 640 2563 642
rect 0 584 2502 640
rect 2558 584 2563 640
rect 0 582 2563 584
rect 0 552 800 582
rect 2497 579 2563 582
rect 19057 642 19123 645
rect 22000 642 22800 672
rect 19057 640 22800 642
rect 19057 584 19062 640
rect 19118 584 22800 640
rect 19057 582 22800 584
rect 19057 579 19123 582
rect 22000 552 22800 582
rect 0 234 800 264
rect 2865 234 2931 237
rect 0 232 2931 234
rect 0 176 2870 232
rect 2926 176 2931 232
rect 0 174 2931 176
rect 0 144 800 174
rect 2865 171 2931 174
rect 18873 234 18939 237
rect 22000 234 22800 264
rect 18873 232 22800 234
rect 18873 176 18878 232
rect 18934 176 22800 232
rect 18873 174 22800 176
rect 18873 171 18939 174
rect 22000 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 8340 18940 8404 19004
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 12940 18048 13004 18052
rect 12940 17992 12990 18048
rect 12990 17992 13004 18048
rect 12940 17988 13004 17992
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 8340 17444 8404 17508
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 19196 17096 19260 17100
rect 19196 17040 19210 17096
rect 19210 17040 19260 17096
rect 19196 17036 19260 17040
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 19196 12548 19260 12612
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 5212 11460 5276 11524
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 12940 10508 13004 10572
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 8340 9692 8404 9756
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 5212 6156 5276 6220
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 8339 19004 8405 19005
rect 8339 18940 8340 19004
rect 8404 18940 8405 19004
rect 8339 18939 8405 18940
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 8342 17509 8402 18939
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 8339 17508 8405 17509
rect 8339 17444 8340 17508
rect 8404 17444 8405 17508
rect 8339 17443 8405 17444
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 5211 11524 5277 11525
rect 5211 11460 5212 11524
rect 5276 11460 5277 11524
rect 5211 11459 5277 11460
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 5214 6221 5274 11459
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 8342 9757 8402 17443
rect 11240 17440 11560 18464
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 12939 18052 13005 18053
rect 12939 17988 12940 18052
rect 13004 17988 13005 18052
rect 12939 17987 13005 17988
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 12942 10573 13002 17987
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 12939 10572 13005 10573
rect 12939 10508 12940 10572
rect 13004 10508 13005 10572
rect 12939 10507 13005 10508
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 8339 9756 8405 9757
rect 8339 9692 8340 9756
rect 8404 9692 8405 9756
rect 8339 9691 8405 9692
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 5211 6220 5277 6221
rect 5211 6156 5212 6220
rect 5276 6156 5277 6220
rect 5211 6155 5277 6156
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 19195 17100 19261 17101
rect 19195 17036 19196 17100
rect 19260 17036 19261 17100
rect 19195 17035 19261 17036
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 19198 12613 19258 17035
rect 19195 12612 19261 12613
rect 19195 12548 19196 12612
rect 19260 12548 19261 12612
rect 19195 12547 19261 12548
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608762278
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608762278
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608762278
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1608762278
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1608762278
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1608762278
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608762278
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608762278
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608762278
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1608762278
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1608762278
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1608762278
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608762278
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608762278
transform 1 0 16560 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608762278
transform 1 0 17296 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608762278
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1608762278
transform 1 0 16928 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1608762278
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608762278
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608762278
transform 1 0 16008 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608762278
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608762278
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_147
timestamp 1608762278
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1608762278
transform 1 0 15180 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1608762278
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_166
timestamp 1608762278
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608762278
transform 1 0 14260 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608762278
transform 1 0 13708 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_134
timestamp 1608762278
transform 1 0 13432 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1608762278
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608762278
transform 1 0 11960 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1608762278
transform 1 0 12604 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608762278
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_115
timestamp 1608762278
transform 1 0 11684 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1608762278
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1608762278
transform 1 0 9752 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608762278
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1608762278
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_103
timestamp 1608762278
transform 1 0 10580 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608762278
transform 1 0 8096 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1608762278
transform 1 0 7084 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608762278
transform 1 0 8648 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp 1608762278
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_74
timestamp 1608762278
transform 1 0 7912 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_80
timestamp 1608762278
transform 1 0 8464 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608762278
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608762278
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1608762278
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608762278
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1608762278
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608762278
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608762278
transform 1 0 1840 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608762278
transform 1 0 2392 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608762278
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1608762278
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1608762278
transform 1 0 1748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1608762278
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_18
timestamp 1608762278
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608762278
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608762278
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1608762278
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1608762278
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1608762278
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608762278
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608762278
transform 1 0 19412 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 18676 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_189
timestamp 1608762278
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1608762278
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1608762278
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608762278
transform 1 0 18124 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1608762278
transform 1 0 16836 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608762278
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_170
timestamp 1608762278
transform 1 0 16744 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1608762278
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1608762278
transform 1 0 18032 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608762278
transform 1 0 14720 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608762278
transform 1 0 16008 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 15272 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1608762278
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_152
timestamp 1608762278
transform 1 0 15088 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_160
timestamp 1608762278
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_166
timestamp 1608762278
transform 1 0 16376 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608762278
transform 1 0 13524 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 13984 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_133
timestamp 1608762278
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_138
timestamp 1608762278
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1608762278
transform 1 0 12512 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608762278
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_116
timestamp 1608762278
transform 1 0 11776 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_123
timestamp 1608762278
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 10304 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 9568 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_88
timestamp 1608762278
transform 1 0 9200 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_98
timestamp 1608762278
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 7728 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 6992 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1608762278
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608762278
transform 1 0 5520 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608762278
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_42
timestamp 1608762278
transform 1 0 4968 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_52
timestamp 1608762278
transform 1 0 5888 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1608762278
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1608762278
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608762278
transform 1 0 3312 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608762278
transform 1 0 3864 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_28
timestamp 1608762278
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1608762278
transform 1 0 1840 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608762278
transform 1 0 2392 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608762278
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1608762278
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1608762278
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_12
timestamp 1608762278
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_18
timestamp 1608762278
transform 1 0 2760 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608762278
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608762278
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608762278
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1608762278
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_218
timestamp 1608762278
transform 1 0 21160 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608762278
transform 1 0 18768 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608762278
transform 1 0 19780 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1608762278
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1608762278
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 18032 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1608762278
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 16376 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1608762278
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608762278
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1608762278
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_163
timestamp 1608762278
transform 1 0 16100 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 13340 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_131
timestamp 1608762278
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 11684 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_30_109
timestamp 1608762278
transform 1 0 11132 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608762278
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_86
timestamp 1608762278
transform 1 0 9016 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1608762278
transform 1 0 8188 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_75
timestamp 1608762278
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 6532 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_48
timestamp 1608762278
transform 1 0 5520 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_56
timestamp 1608762278
transform 1 0 6256 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608762278
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608762278
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_24
timestamp 1608762278
transform 1 0 3312 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1608762278
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_36
timestamp 1608762278
transform 1 0 4416 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608762278
transform 1 0 1840 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608762278
transform 1 0 2392 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608762278
transform 1 0 2944 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608762278
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1608762278
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1608762278
transform 1 0 1748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1608762278
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1608762278
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608762278
transform 1 0 20700 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608762278
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_211
timestamp 1608762278
transform 1 0 20516 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_217
timestamp 1608762278
transform 1 0 21068 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1608762278
transform 1 0 19688 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_200
timestamp 1608762278
transform 1 0 19504 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608762278
transform 1 0 17388 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 18032 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608762278
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1608762278
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1608762278
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 15732 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_157
timestamp 1608762278
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608762278
transform 1 0 13524 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 14076 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_133
timestamp 1608762278
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1608762278
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1608762278
transform 1 0 11040 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1608762278
transform 1 0 12512 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608762278
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_105
timestamp 1608762278
transform 1 0 10764 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1608762278
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1608762278
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_123
timestamp 1608762278
transform 1 0 12420 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608762278
transform 1 0 10488 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608762278
transform 1 0 9476 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_100
timestamp 1608762278
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608762278
transform 1 0 8464 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1608762278
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_83
timestamp 1608762278
transform 1 0 8740 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 6808 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 5888 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608762278
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_49
timestamp 1608762278
transform 1 0 5612 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_58
timestamp 1608762278
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608762278
transform 1 0 3404 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1608762278
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_29
timestamp 1608762278
transform 1 0 3772 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_41
timestamp 1608762278
transform 1 0 4876 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608762278
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608762278
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608762278
transform 1 0 2852 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608762278
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1608762278
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1608762278
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1608762278
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608762278
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608762278
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608762278
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1608762278
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_218
timestamp 1608762278
transform 1 0 21160 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608762278
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 18584 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1608762278
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1608762278
transform 1 0 16468 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1608762278
transform 1 0 17480 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_176
timestamp 1608762278
transform 1 0 17296 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_187
timestamp 1608762278
transform 1 0 18308 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1608762278
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608762278
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1608762278
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1608762278
transform 1 0 16100 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 13064 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1608762278
transform 1 0 14168 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_128
timestamp 1608762278
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_136
timestamp 1608762278
transform 1 0 13616 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1608762278
transform 1 0 12052 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_117
timestamp 1608762278
transform 1 0 11868 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608762278
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 10396 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608762278
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1608762278
transform 1 0 8924 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1608762278
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_97
timestamp 1608762278
transform 1 0 10028 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1608762278
transform 1 0 7084 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1608762278
transform 1 0 8096 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1608762278
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_74
timestamp 1608762278
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608762278
transform 1 0 5796 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 5060 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_49
timestamp 1608762278
transform 1 0 5612 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_55
timestamp 1608762278
transform 1 0 6164 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608762278
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1608762278
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_32
timestamp 1608762278
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_40
timestamp 1608762278
transform 1 0 4784 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608762278
transform 1 0 1656 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 2208 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608762278
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1608762278
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1608762278
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_18
timestamp 1608762278
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608762278
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608762278
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1608762278
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1608762278
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608762278
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1608762278
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1608762278
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608762278
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1608762278
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1608762278
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1608762278
transform 1 0 20056 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608762278
transform 1 0 18400 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 18952 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1608762278
transform 1 0 19044 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_192
timestamp 1608762278
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1608762278
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_204
timestamp 1608762278
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 16468 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1608762278
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 17112 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608762278
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1608762278
transform 1 0 17940 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_187
timestamp 1608762278
transform 1 0 18308 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_171
timestamp 1608762278
transform 1 0 16836 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1608762278
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1608762278
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 15364 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 16284 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608762278
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1608762278
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1608762278
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_153
timestamp 1608762278
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_161
timestamp 1608762278
transform 1 0 15916 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1608762278
transform 1 0 12972 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1608762278
transform 1 0 13064 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1608762278
transform 1 0 13984 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1608762278
transform 1 0 14352 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_26_128
timestamp 1608762278
transform 1 0 12880 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1608762278
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_128
timestamp 1608762278
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1608762278
transform 1 0 13892 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_143
timestamp 1608762278
transform 1 0 14260 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608762278
transform 1 0 12604 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1608762278
transform 1 0 12512 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1608762278
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608762278
transform 1 0 11684 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608762278
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1608762278
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1608762278
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1608762278
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1608762278
transform 1 0 10856 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_113
timestamp 1608762278
transform 1 0 11500 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608762278
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 8832 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1608762278
transform 1 0 10672 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608762278
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_86
timestamp 1608762278
transform 1 0 9016 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1608762278
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_90
timestamp 1608762278
transform 1 0 9384 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_102
timestamp 1608762278
transform 1 0 10488 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 7544 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608762278
transform 1 0 7820 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_68
timestamp 1608762278
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1608762278
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_82
timestamp 1608762278
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 5888 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1608762278
transform 1 0 5428 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608762278
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608762278
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_50
timestamp 1608762278
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_45
timestamp 1608762278
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_56
timestamp 1608762278
transform 1 0 6256 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1608762278
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608762278
transform 1 0 3404 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762278
transform 1 0 4232 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608762278
transform 1 0 4416 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608762278
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_25
timestamp 1608762278
transform 1 0 3404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1608762278
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1608762278
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_29
timestamp 1608762278
transform 1 0 3772 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_35
timestamp 1608762278
transform 1 0 4324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1608762278
transform 1 0 2300 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608762278
transform 1 0 2852 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608762278
transform 1 0 2576 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1608762278
transform 1 0 2116 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1608762278
transform 1 0 2484 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1608762278
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1608762278
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1608762278
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1608762278
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608762278
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608762278
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1608762278
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1608762278
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608762278
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608762278
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1608762278
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1608762278
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1608762278
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 18860 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_191
timestamp 1608762278
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608762278
transform 1 0 18308 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1608762278
transform 1 0 16836 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608762278
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1608762278
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1608762278
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_184
timestamp 1608762278
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608762278
transform 1 0 16284 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 14628 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_163
timestamp 1608762278
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 12972 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_128
timestamp 1608762278
transform 1 0 12880 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1608762278
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 11592 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608762278
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 12604 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_111
timestamp 1608762278
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1608762278
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1608762278
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608762278
transform 1 0 10488 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_99
timestamp 1608762278
transform 1 0 10212 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 8740 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 8464 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1608762278
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608762278
transform 1 0 4968 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608762278
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 5980 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_51
timestamp 1608762278
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_56
timestamp 1608762278
transform 1 0 6256 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1608762278
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 3036 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_37
timestamp 1608762278
transform 1 0 4508 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_41
timestamp 1608762278
transform 1 0 4876 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1608762278
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1608762278
transform 1 0 2300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608762278
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1608762278
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1608762278
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_17
timestamp 1608762278
transform 1 0 2668 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608762278
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608762278
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1608762278
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1608762278
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608762278
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 20056 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1608762278
transform 1 0 19044 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1608762278
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_204
timestamp 1608762278
transform 1 0 19872 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1608762278
transform 1 0 18032 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608762278
transform 1 0 17020 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_171
timestamp 1608762278
transform 1 0 16836 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1608762278
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 15364 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608762278
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1608762278
transform 1 0 14720 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1608762278
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_154
timestamp 1608762278
transform 1 0 15272 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608762278
transform 1 0 13892 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_137
timestamp 1608762278
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 12236 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_119
timestamp 1608762278
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608762278
transform 1 0 9016 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 10580 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608762278
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1608762278
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1608762278
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_93
timestamp 1608762278
transform 1 0 9660 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1608762278
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1608762278
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608762278
transform 1 0 6992 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_73
timestamp 1608762278
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1608762278
transform 1 0 5612 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_47
timestamp 1608762278
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_58
timestamp 1608762278
transform 1 0 6440 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1608762278
transform 1 0 4600 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608762278
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1608762278
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_32
timestamp 1608762278
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1608762278
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608762278
transform 1 0 2760 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608762278
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1608762278
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_11
timestamp 1608762278
transform 1 0 2116 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_17
timestamp 1608762278
transform 1 0 2668 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 20516 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608762278
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1608762278
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_217
timestamp 1608762278
transform 1 0 21068 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 19780 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_200
timestamp 1608762278
transform 1 0 19504 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 18032 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608762278
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1608762278
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 16284 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1608762278
transform 1 0 14904 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 15916 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_159
timestamp 1608762278
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_164
timestamp 1608762278
transform 1 0 16192 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608762278
transform 1 0 13248 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1608762278
transform 1 0 14076 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1608762278
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1608762278
transform 1 0 11316 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608762278
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_109
timestamp 1608762278
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608762278
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 9660 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_88
timestamp 1608762278
transform 1 0 9200 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_92
timestamp 1608762278
transform 1 0 9568 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1608762278
transform 1 0 7360 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1608762278
transform 1 0 8372 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_77
timestamp 1608762278
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1608762278
transform 1 0 5152 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1608762278
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608762278
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1608762278
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 1608762278
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1608762278
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_62
timestamp 1608762278
transform 1 0 6808 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1608762278
transform 1 0 4140 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_29
timestamp 1608762278
transform 1 0 3772 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 2300 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 1564 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608762278
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1608762278
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1608762278
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608762278
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608762278
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608762278
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1608762278
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1608762278
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608762278
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608762278
transform 1 0 18676 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1608762278
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_189
timestamp 1608762278
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_195
timestamp 1608762278
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1608762278
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608762278
transform 1 0 16468 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 17020 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1608762278
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608762278
transform 1 0 14720 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1608762278
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608762278
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1608762278
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1608762278
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1608762278
transform 1 0 12880 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 13892 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_127
timestamp 1608762278
transform 1 0 12788 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_137
timestamp 1608762278
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_142
timestamp 1608762278
transform 1 0 14168 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608762278
transform 1 0 12144 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608762278
transform 1 0 11316 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_22_105
timestamp 1608762278
transform 1 0 10764 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_123
timestamp 1608762278
transform 1 0 12420 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608762278
transform 1 0 9936 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608762278
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1608762278
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1608762278
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 7360 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 6992 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_67
timestamp 1608762278
transform 1 0 7268 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 5336 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_44
timestamp 1608762278
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_62
timestamp 1608762278
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608762278
transform 1 0 4324 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608762278
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608762278
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 1608762278
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1608762278
transform 1 0 1748 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1608762278
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608762278
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1608762278
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_16
timestamp 1608762278
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1608762278
transform 1 0 20332 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608762278
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_218
timestamp 1608762278
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1608762278
transform 1 0 19320 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_193
timestamp 1608762278
transform 1 0 18860 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_197
timestamp 1608762278
transform 1 0 19228 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_207
timestamp 1608762278
transform 1 0 20148 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608762278
transform 1 0 16928 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1608762278
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608762278
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_168
timestamp 1608762278
transform 1 0 16560 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1608762278
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1608762278
transform 1 0 15732 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1608762278
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 14076 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1608762278
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608762278
transform 1 0 10856 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608762278
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1608762278
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1608762278
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608762278
transform 1 0 9016 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608762278
transform 1 0 10028 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1608762278
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 6992 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_21_80
timestamp 1608762278
transform 1 0 8464 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608762278
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1608762278
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1608762278
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 3220 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1608762278
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1608762278
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1608762278
transform 1 0 2668 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1608762278
transform 1 0 1656 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608762278
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1608762278
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1608762278
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608762278
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608762278
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608762278
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_214
timestamp 1608762278
transform 1 0 20792 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1608762278
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1608762278
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608762278
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608762278
transform 1 0 20240 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762278
transform 1 0 18584 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1608762278
transform 1 0 19964 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1608762278
transform 1 0 19504 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_204
timestamp 1608762278
transform 1 0 19872 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1608762278
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 16560 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 18032 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1608762278
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608762278
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_171
timestamp 1608762278
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1608762278
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_184
timestamp 1608762278
transform 1 0 18032 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608762278
transform 1 0 16008 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1608762278
transform 1 0 15456 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608762278
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1608762278
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_165
timestamp 1608762278
transform 1 0 16284 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1608762278
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1608762278
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_165
timestamp 1608762278
transform 1 0 16284 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 14352 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608762278
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1608762278
transform 1 0 14168 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1608762278
transform 1 0 12972 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_128
timestamp 1608762278
transform 1 0 12880 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_138
timestamp 1608762278
transform 1 0 13800 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_128
timestamp 1608762278
transform 1 0 12880 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_138
timestamp 1608762278
transform 1 0 13800 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 11408 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608762278
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 12604 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1608762278
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1608762278
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 9936 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608762278
transform 1 0 8924 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608762278
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 10304 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_19_94
timestamp 1608762278
transform 1 0 9752 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1608762278
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1608762278
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1608762278
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1608762278
transform 1 0 6900 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1608762278
transform 1 0 7084 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608762278
transform 1 0 8280 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1608762278
transform 1 0 7912 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_72
timestamp 1608762278
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_83
timestamp 1608762278
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_63
timestamp 1608762278
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_74
timestamp 1608762278
transform 1 0 7912 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608762278
transform 1 0 6072 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608762278
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_47
timestamp 1608762278
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608762278
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1608762278
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_44
timestamp 1608762278
transform 1 0 5152 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_52
timestamp 1608762278
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608762278
transform 1 0 4140 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1608762278
transform 1 0 4600 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1608762278
transform 1 0 4324 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608762278
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_32
timestamp 1608762278
transform 1 0 4048 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1608762278
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1608762278
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 3220 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1608762278
transform 1 0 3680 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1608762278
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1608762278
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 2208 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1608762278
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1608762278
transform 1 0 1656 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 1472 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608762278
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608762278
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1608762278
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_10
timestamp 1608762278
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1608762278
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1608762278
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1608762278
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608762278
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608762278
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1608762278
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1608762278
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 19044 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1608762278
transform 1 0 19780 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_192
timestamp 1608762278
transform 1 0 18768 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1608762278
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1608762278
transform 1 0 17940 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_181
timestamp 1608762278
transform 1 0 17756 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608762278
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762278
transform 1 0 16284 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608762278
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1608762278
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_157
timestamp 1608762278
transform 1 0 15548 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1608762278
transform 1 0 14168 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608762278
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 13800 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_126
timestamp 1608762278
transform 1 0 12696 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_136
timestamp 1608762278
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1608762278
transform 1 0 14076 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 10856 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_122
timestamp 1608762278
transform 1 0 12328 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608762278
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608762278
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1608762278
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1608762278
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 7268 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_65
timestamp 1608762278
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_83
timestamp 1608762278
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 5612 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_43
timestamp 1608762278
transform 1 0 5060 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1608762278
transform 1 0 4232 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608762278
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_28
timestamp 1608762278
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1608762278
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762278
transform 1 0 1472 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608762278
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1608762278
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1608762278
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608762278
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1608762278
transform 1 0 20976 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1608762278
transform 1 0 19136 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1608762278
transform 1 0 20148 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_194
timestamp 1608762278
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_205
timestamp 1608762278
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 17204 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1608762278
transform 1 0 18124 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608762278
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_172
timestamp 1608762278
transform 1 0 16928 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1608762278
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1608762278
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1608762278
transform 1 0 15088 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608762278
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1608762278
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1608762278
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608762278
transform 1 0 14076 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1608762278
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1608762278
transform 1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608762278
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1608762278
transform 1 0 10948 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608762278
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608762278
transform 1 0 10120 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1608762278
transform 1 0 9660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 1608762278
transform 1 0 10028 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608762278
transform 1 0 6992 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 8188 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 7820 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_67
timestamp 1608762278
transform 1 0 7268 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_76
timestamp 1608762278
transform 1 0 8096 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608762278
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1608762278
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608762278
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1608762278
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762278
transform 1 0 4324 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1608762278
transform 1 0 3312 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_22
timestamp 1608762278
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_33
timestamp 1608762278
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608762278
transform 1 0 1472 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1608762278
transform 1 0 2300 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608762278
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1608762278
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_7
timestamp 1608762278
transform 1 0 1748 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608762278
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608762278
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1608762278
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1608762278
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1608762278
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1608762278
transform 1 0 18676 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608762278
transform 1 0 19688 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_189
timestamp 1608762278
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_200
timestamp 1608762278
transform 1 0 19504 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608762278
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1608762278
transform 1 0 17204 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_179
timestamp 1608762278
transform 1 0 17572 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 15732 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608762278
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 15456 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1608762278
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1608762278
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 12696 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_142
timestamp 1608762278
transform 1 0 14168 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608762278
transform 1 0 11684 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_113
timestamp 1608762278
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_124
timestamp 1608762278
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608762278
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608762278
transform 1 0 10672 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608762278
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1608762278
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1608762278
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1608762278
transform 1 0 7176 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608762278
transform 1 0 8188 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_64
timestamp 1608762278
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_75
timestamp 1608762278
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608762278
transform 1 0 6164 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608762278
transform 1 0 5060 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_52
timestamp 1608762278
transform 1 0 5888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1608762278
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608762278
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1608762278
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1608762278
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608762278
transform 1 0 2944 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1608762278
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608762278
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1608762278
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1608762278
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1608762278
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 20608 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608762278
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_210
timestamp 1608762278
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1608762278
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608762278
transform 1 0 18584 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1608762278
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1608762278
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1608762278
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608762278
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_174
timestamp 1608762278
transform 1 0 17112 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1608762278
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_187
timestamp 1608762278
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 14628 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608762278
transform 1 0 16284 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1608762278
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1608762278
transform 1 0 13616 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_134
timestamp 1608762278
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1608762278
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1608762278
transform 1 0 12604 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608762278
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1608762278
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1608762278
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 10488 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1608762278
transform 1 0 9476 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1608762278
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1608762278
transform 1 0 7544 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_67
timestamp 1608762278
transform 1 0 7268 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_79
timestamp 1608762278
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608762278
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608762278
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 5060 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_46
timestamp 1608762278
transform 1 0 5336 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608762278
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1608762278
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 3404 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_24
timestamp 1608762278
transform 1 0 3312 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_41
timestamp 1608762278
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 1472 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608762278
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1608762278
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1608762278
transform 1 0 2944 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608762278
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608762278
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608762278
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_213
timestamp 1608762278
transform 1 0 20700 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1608762278
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1608762278
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1608762278
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1608762278
transform 1 0 19872 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1608762278
transform 1 0 18860 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1608762278
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_191
timestamp 1608762278
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_202
timestamp 1608762278
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_193
timestamp 1608762278
transform 1 0 18860 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1608762278
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1608762278
transform 1 0 16836 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 18124 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1608762278
transform 1 0 18032 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608762278
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1608762278
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1608762278
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1608762278
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_184
timestamp 1608762278
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_179
timestamp 1608762278
transform 1 0 17572 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762278
transform 1 0 15180 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 16100 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608762278
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1608762278
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1608762278
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1608762278
transform 1 0 15272 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_162
timestamp 1608762278
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608762278
transform 1 0 12696 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 13524 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1608762278
transform 1 0 13340 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_132
timestamp 1608762278
transform 1 0 13248 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 1608762278
transform 1 0 12972 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_142
timestamp 1608762278
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 10856 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1608762278
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608762278
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_116
timestamp 1608762278
transform 1 0 11776 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_122
timestamp 1608762278
transform 1 0 12328 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608762278
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608762278
transform 1 0 9844 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608762278
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1608762278
transform 1 0 9476 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_104
timestamp 1608762278
transform 1 0 10672 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1608762278
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1608762278
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 8004 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1608762278
transform 1 0 6992 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk
timestamp 1608762278
transform 1 0 7636 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_73
timestamp 1608762278
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1608762278
transform 1 0 7084 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 5612 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608762278
transform 1 0 5612 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608762278
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_46
timestamp 1608762278
transform 1 0 5336 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_58
timestamp 1608762278
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1608762278
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_47
timestamp 1608762278
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608762278
transform 1 0 4140 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1608762278
transform 1 0 4600 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1608762278
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608762278
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_34
timestamp 1608762278
transform 1 0 4232 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1608762278
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1608762278
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1608762278
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 2760 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1608762278
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1608762278
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_18
timestamp 1608762278
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1608762278
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1608762278
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1608762278
transform 1 0 1748 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608762278
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608762278
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1608762278
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1608762278
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608762278
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608762278
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1608762278
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1608762278
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1608762278
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762278
transform 1 0 18492 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_205
timestamp 1608762278
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608762278
transform 1 0 17296 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_174
timestamp 1608762278
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_179
timestamp 1608762278
transform 1 0 17572 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_187
timestamp 1608762278
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1608762278
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1608762278
transform 1 0 16284 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608762278
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1608762278
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1608762278
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608762278
transform 1 0 14168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_12_135
timestamp 1608762278
transform 1 0 13524 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1608762278
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 12052 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_12_113
timestamp 1608762278
transform 1 0 11500 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 10028 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608762278
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1608762278
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1608762278
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608762278
transform 1 0 8464 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608762278
transform 1 0 7452 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_66
timestamp 1608762278
transform 1 0 7176 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_78
timestamp 1608762278
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_83
timestamp 1608762278
transform 1 0 8740 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1608762278
transform 1 0 5244 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_43
timestamp 1608762278
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1608762278
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 3220 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1608762278
transform 1 0 4232 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608762278
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_21
timestamp 1608762278
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1608762278
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1608762278
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 1472 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1608762278
transform 1 0 2208 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608762278
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1608762278
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1608762278
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608762278
transform 1 0 20792 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608762278
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1608762278
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_217
timestamp 1608762278
transform 1 0 21068 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608762278
transform 1 0 19780 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_200
timestamp 1608762278
transform 1 0 19504 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 18032 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608762278
transform 1 0 16560 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608762278
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1608762278
transform 1 0 16468 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_177
timestamp 1608762278
transform 1 0 17388 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608762278
transform 1 0 15272 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_150
timestamp 1608762278
transform 1 0 14904 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp 1608762278
transform 1 0 16100 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608762278
transform 1 0 14076 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1608762278
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608762278
transform 1 0 11224 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608762278
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_108
timestamp 1608762278
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1608762278
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608762278
transform 1 0 10212 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1608762278
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 8556 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608762278
transform 1 0 6992 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_73
timestamp 1608762278
transform 1 0 7820 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608762278
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608762278
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_47
timestamp 1608762278
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608762278
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1608762278
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608762278
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1608762278
transform 1 0 4600 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1608762278
transform 1 0 3128 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_26
timestamp 1608762278
transform 1 0 3496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_36
timestamp 1608762278
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762278
transform 1 0 1656 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608762278
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1608762278
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608762278
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608762278
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1608762278
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1608762278
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1608762278
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608762278
transform 1 0 18676 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1608762278
transform 1 0 19780 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1608762278
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_200
timestamp 1608762278
transform 1 0 19504 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 17020 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_171
timestamp 1608762278
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1608762278
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608762278
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_146
timestamp 1608762278
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1608762278
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_163
timestamp 1608762278
transform 1 0 16100 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_134
timestamp 1608762278
transform 1 0 13432 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608762278
transform 1 0 12604 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_113
timestamp 1608762278
transform 1 0 11500 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608762278
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608762278
transform 1 0 10672 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608762278
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1608762278
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1608762278
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1608762278
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608762278
transform 1 0 7268 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608762278
transform 1 0 8280 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1608762278
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_76
timestamp 1608762278
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762278
transform 1 0 5612 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_47
timestamp 1608762278
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1608762278
transform 1 0 4600 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608762278
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608762278
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1608762278
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1608762278
transform 1 0 2760 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1608762278
transform 1 0 1748 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608762278
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1608762278
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_16
timestamp 1608762278
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608762278
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_217
timestamp 1608762278
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608762278
transform 1 0 19228 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1608762278
transform 1 0 20240 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1608762278
transform 1 0 18860 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_206
timestamp 1608762278
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608762278
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608762278
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1608762278
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1608762278
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1608762278
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1608762278
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608762278
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_108
timestamp 1608762278
transform 1 0 11040 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608762278
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1608762278
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_96
timestamp 1608762278
transform 1 0 9936 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 8464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1608762278
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 4968 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608762278
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1608762278
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608762278
transform 1 0 3956 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_29
timestamp 1608762278
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1608762278
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762278
transform 1 0 2300 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608762278
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1608762278
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1608762278
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608762278
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608762278
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1608762278
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1608762278
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 18768 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_208
timestamp 1608762278
transform 1 0 20240 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 16560 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_184
timestamp 1608762278
transform 1 0 18032 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608762278
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1608762278
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_166
timestamp 1608762278
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1608762278
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1608762278
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1608762278
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1608762278
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608762278
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1608762278
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1608762278
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1608762278
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608762278
transform 1 0 5980 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1608762278
transform 1 0 4968 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_51
timestamp 1608762278
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1608762278
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608762278
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608762278
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1608762278
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_40
timestamp 1608762278
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1608762278
transform 1 0 2760 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608762278
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608762278
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp 1608762278
transform 1 0 2484 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608762278
transform 1 0 20700 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608762278
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608762278
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608762278
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1608762278
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1608762278
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1608762278
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_211
timestamp 1608762278
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_216
timestamp 1608762278
transform 1 0 20976 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762278
transform 1 0 19044 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1608762278
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1608762278
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_190
timestamp 1608762278
transform 1 0 18584 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_198
timestamp 1608762278
transform 1 0 19320 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1608762278
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762278
transform 1 0 18308 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608762278
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1608762278
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1608762278
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_184
timestamp 1608762278
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608762278
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1608762278
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1608762278
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1608762278
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1608762278
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1608762278
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1608762278
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1608762278
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608762278
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1608762278
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1608762278
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1608762278
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1608762278
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608762278
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1608762278
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1608762278
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1608762278
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1608762278
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1608762278
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1608762278
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1608762278
transform 1 0 5060 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608762278
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608762278
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1608762278
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_42
timestamp 1608762278
transform 1 0 4968 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_52
timestamp 1608762278
transform 1 0 5888 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1608762278
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1608762278
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608762278
transform 1 0 3220 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608762278
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608762278
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608762278
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_21
timestamp 1608762278
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_26
timestamp 1608762278
transform 1 0 3496 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_38
timestamp 1608762278
transform 1 0 4600 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762278
transform 1 0 1564 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608762278
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608762278
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608762278
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608762278
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1608762278
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608762278
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_212
timestamp 1608762278
transform 1 0 20608 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1608762278
transform 1 0 19780 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_196
timestamp 1608762278
transform 1 0 19136 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_202
timestamp 1608762278
transform 1 0 19688 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608762278
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1608762278
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1608762278
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1608762278
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1608762278
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1608762278
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608762278
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1608762278
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1608762278
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1608762278
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1608762278
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1608762278
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608762278
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608762278
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608762278
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608762278
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608762278
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608762278
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608762278
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608762278
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608762278
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608762278
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608762278
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1608762278
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1608762278
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1608762278
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1608762278
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1608762278
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608762278
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1608762278
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1608762278
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1608762278
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1608762278
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1608762278
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1608762278
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608762278
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1608762278
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1608762278
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1608762278
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608762278
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608762278
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608762278
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608762278
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608762278
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608762278
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608762278
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608762278
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608762278
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1608762278
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1608762278
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608762278
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1608762278
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1608762278
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1608762278
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1608762278
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1608762278
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608762278
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1608762278
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1608762278
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1608762278
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1608762278
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1608762278
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608762278
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608762278
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608762278
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608762278
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608762278
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608762278
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608762278
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608762278
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608762278
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608762278
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608762278
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1608762278
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1608762278
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1608762278
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1608762278
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1608762278
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608762278
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1608762278
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1608762278
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1608762278
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1608762278
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1608762278
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1608762278
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608762278
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1608762278
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608762278
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608762278
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608762278
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608762278
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608762278
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608762278
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608762278
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608762278
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608762278
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608762278
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608762278
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608762278
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608762278
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1608762278
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1608762278
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1608762278
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1608762278
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1608762278
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608762278
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608762278
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1608762278
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1608762278
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1608762278
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1608762278
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1608762278
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1608762278
transform 1 0 15180 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608762278
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608762278
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1608762278
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_147
timestamp 1608762278
transform 1 0 14628 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1608762278
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1608762278
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1608762278
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608762278
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608762278
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608762278
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608762278
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608762278
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1608762278
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1608762278
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608762278
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608762278
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608762278
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1608762278
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1608762278
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608762278
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608762278
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1608762278
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1608762278
transform 1 0 5520 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608762278
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608762278
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608762278
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608762278
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1608762278
transform 1 0 5152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_54
timestamp 1608762278
transform 1 0 6072 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1608762278
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608762278
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1608762278
transform 1 0 4600 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608762278
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608762278
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608762278
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp 1608762278
transform 1 0 3588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_35
timestamp 1608762278
transform 1 0 4324 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608762278
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608762278
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608762278
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608762278
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608762278
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1608762278
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 202 22000 258 22800 4 SC_IN_TOP
port 1 nsew
rlabel metal2 s 22558 22000 22614 22800 4 SC_OUT_TOP
port 2 nsew
rlabel metal2 s 4342 22000 4398 22800 4 Test_en_N_out
port 3 nsew
rlabel metal2 s 20442 0 20498 800 4 Test_en_S_in
port 4 nsew
rlabel metal2 s 2226 0 2282 800 4 ccff_head
port 5 nsew
rlabel metal2 s 6734 0 6790 800 4 ccff_tail
port 6 nsew
rlabel metal3 s 0 4224 800 4344 4 chanx_left_in[0]
port 7 nsew
rlabel metal3 s 0 8984 800 9104 4 chanx_left_in[10]
port 8 nsew
rlabel metal3 s 0 9392 800 9512 4 chanx_left_in[11]
port 9 nsew
rlabel metal3 s 0 9936 800 10056 4 chanx_left_in[12]
port 10 nsew
rlabel metal3 s 0 10344 800 10464 4 chanx_left_in[13]
port 11 nsew
rlabel metal3 s 0 10752 800 10872 4 chanx_left_in[14]
port 12 nsew
rlabel metal3 s 0 11296 800 11416 4 chanx_left_in[15]
port 13 nsew
rlabel metal3 s 0 11704 800 11824 4 chanx_left_in[16]
port 14 nsew
rlabel metal3 s 0 12248 800 12368 4 chanx_left_in[17]
port 15 nsew
rlabel metal3 s 0 12656 800 12776 4 chanx_left_in[18]
port 16 nsew
rlabel metal3 s 0 13200 800 13320 4 chanx_left_in[19]
port 17 nsew
rlabel metal3 s 0 4768 800 4888 4 chanx_left_in[1]
port 18 nsew
rlabel metal3 s 0 5176 800 5296 4 chanx_left_in[2]
port 19 nsew
rlabel metal3 s 0 5720 800 5840 4 chanx_left_in[3]
port 20 nsew
rlabel metal3 s 0 6128 800 6248 4 chanx_left_in[4]
port 21 nsew
rlabel metal3 s 0 6672 800 6792 4 chanx_left_in[5]
port 22 nsew
rlabel metal3 s 0 7080 800 7200 4 chanx_left_in[6]
port 23 nsew
rlabel metal3 s 0 7488 800 7608 4 chanx_left_in[7]
port 24 nsew
rlabel metal3 s 0 8032 800 8152 4 chanx_left_in[8]
port 25 nsew
rlabel metal3 s 0 8440 800 8560 4 chanx_left_in[9]
port 26 nsew
rlabel metal3 s 0 13608 800 13728 4 chanx_left_out[0]
port 27 nsew
rlabel metal3 s 0 18232 800 18352 4 chanx_left_out[10]
port 28 nsew
rlabel metal3 s 0 18776 800 18896 4 chanx_left_out[11]
port 29 nsew
rlabel metal3 s 0 19184 800 19304 4 chanx_left_out[12]
port 30 nsew
rlabel metal3 s 0 19728 800 19848 4 chanx_left_out[13]
port 31 nsew
rlabel metal3 s 0 20136 800 20256 4 chanx_left_out[14]
port 32 nsew
rlabel metal3 s 0 20544 800 20664 4 chanx_left_out[15]
port 33 nsew
rlabel metal3 s 0 21088 800 21208 4 chanx_left_out[16]
port 34 nsew
rlabel metal3 s 0 21496 800 21616 4 chanx_left_out[17]
port 35 nsew
rlabel metal3 s 0 22040 800 22160 4 chanx_left_out[18]
port 36 nsew
rlabel metal3 s 0 22448 800 22568 4 chanx_left_out[19]
port 37 nsew
rlabel metal3 s 0 14016 800 14136 4 chanx_left_out[1]
port 38 nsew
rlabel metal3 s 0 14560 800 14680 4 chanx_left_out[2]
port 39 nsew
rlabel metal3 s 0 14968 800 15088 4 chanx_left_out[3]
port 40 nsew
rlabel metal3 s 0 15512 800 15632 4 chanx_left_out[4]
port 41 nsew
rlabel metal3 s 0 15920 800 16040 4 chanx_left_out[5]
port 42 nsew
rlabel metal3 s 0 16464 800 16584 4 chanx_left_out[6]
port 43 nsew
rlabel metal3 s 0 16872 800 16992 4 chanx_left_out[7]
port 44 nsew
rlabel metal3 s 0 17280 800 17400 4 chanx_left_out[8]
port 45 nsew
rlabel metal3 s 0 17824 800 17944 4 chanx_left_out[9]
port 46 nsew
rlabel metal3 s 22000 4224 22800 4344 4 chanx_right_in[0]
port 47 nsew
rlabel metal3 s 22000 8984 22800 9104 4 chanx_right_in[10]
port 48 nsew
rlabel metal3 s 22000 9392 22800 9512 4 chanx_right_in[11]
port 49 nsew
rlabel metal3 s 22000 9936 22800 10056 4 chanx_right_in[12]
port 50 nsew
rlabel metal3 s 22000 10344 22800 10464 4 chanx_right_in[13]
port 51 nsew
rlabel metal3 s 22000 10752 22800 10872 4 chanx_right_in[14]
port 52 nsew
rlabel metal3 s 22000 11296 22800 11416 4 chanx_right_in[15]
port 53 nsew
rlabel metal3 s 22000 11704 22800 11824 4 chanx_right_in[16]
port 54 nsew
rlabel metal3 s 22000 12248 22800 12368 4 chanx_right_in[17]
port 55 nsew
rlabel metal3 s 22000 12656 22800 12776 4 chanx_right_in[18]
port 56 nsew
rlabel metal3 s 22000 13200 22800 13320 4 chanx_right_in[19]
port 57 nsew
rlabel metal3 s 22000 4768 22800 4888 4 chanx_right_in[1]
port 58 nsew
rlabel metal3 s 22000 5176 22800 5296 4 chanx_right_in[2]
port 59 nsew
rlabel metal3 s 22000 5720 22800 5840 4 chanx_right_in[3]
port 60 nsew
rlabel metal3 s 22000 6128 22800 6248 4 chanx_right_in[4]
port 61 nsew
rlabel metal3 s 22000 6672 22800 6792 4 chanx_right_in[5]
port 62 nsew
rlabel metal3 s 22000 7080 22800 7200 4 chanx_right_in[6]
port 63 nsew
rlabel metal3 s 22000 7488 22800 7608 4 chanx_right_in[7]
port 64 nsew
rlabel metal3 s 22000 8032 22800 8152 4 chanx_right_in[8]
port 65 nsew
rlabel metal3 s 22000 8440 22800 8560 4 chanx_right_in[9]
port 66 nsew
rlabel metal3 s 22000 13608 22800 13728 4 chanx_right_out[0]
port 67 nsew
rlabel metal3 s 22000 18232 22800 18352 4 chanx_right_out[10]
port 68 nsew
rlabel metal3 s 22000 18776 22800 18896 4 chanx_right_out[11]
port 69 nsew
rlabel metal3 s 22000 19184 22800 19304 4 chanx_right_out[12]
port 70 nsew
rlabel metal3 s 22000 19728 22800 19848 4 chanx_right_out[13]
port 71 nsew
rlabel metal3 s 22000 20136 22800 20256 4 chanx_right_out[14]
port 72 nsew
rlabel metal3 s 22000 20544 22800 20664 4 chanx_right_out[15]
port 73 nsew
rlabel metal3 s 22000 21088 22800 21208 4 chanx_right_out[16]
port 74 nsew
rlabel metal3 s 22000 21496 22800 21616 4 chanx_right_out[17]
port 75 nsew
rlabel metal3 s 22000 22040 22800 22160 4 chanx_right_out[18]
port 76 nsew
rlabel metal3 s 22000 22448 22800 22568 4 chanx_right_out[19]
port 77 nsew
rlabel metal3 s 22000 14016 22800 14136 4 chanx_right_out[1]
port 78 nsew
rlabel metal3 s 22000 14560 22800 14680 4 chanx_right_out[2]
port 79 nsew
rlabel metal3 s 22000 14968 22800 15088 4 chanx_right_out[3]
port 80 nsew
rlabel metal3 s 22000 15512 22800 15632 4 chanx_right_out[4]
port 81 nsew
rlabel metal3 s 22000 15920 22800 16040 4 chanx_right_out[5]
port 82 nsew
rlabel metal3 s 22000 16464 22800 16584 4 chanx_right_out[6]
port 83 nsew
rlabel metal3 s 22000 16872 22800 16992 4 chanx_right_out[7]
port 84 nsew
rlabel metal3 s 22000 17280 22800 17400 4 chanx_right_out[8]
port 85 nsew
rlabel metal3 s 22000 17824 22800 17944 4 chanx_right_out[9]
port 86 nsew
rlabel metal2 s 5630 22000 5686 22800 4 chany_top_in[0]
port 87 nsew
rlabel metal2 s 9862 22000 9918 22800 4 chany_top_in[10]
port 88 nsew
rlabel metal2 s 10322 22000 10378 22800 4 chany_top_in[11]
port 89 nsew
rlabel metal2 s 10690 22000 10746 22800 4 chany_top_in[12]
port 90 nsew
rlabel metal2 s 11150 22000 11206 22800 4 chany_top_in[13]
port 91 nsew
rlabel metal2 s 11610 22000 11666 22800 4 chany_top_in[14]
port 92 nsew
rlabel metal2 s 11978 22000 12034 22800 4 chany_top_in[15]
port 93 nsew
rlabel metal2 s 12438 22000 12494 22800 4 chany_top_in[16]
port 94 nsew
rlabel metal2 s 12806 22000 12862 22800 4 chany_top_in[17]
port 95 nsew
rlabel metal2 s 13266 22000 13322 22800 4 chany_top_in[18]
port 96 nsew
rlabel metal2 s 13634 22000 13690 22800 4 chany_top_in[19]
port 97 nsew
rlabel metal2 s 6090 22000 6146 22800 4 chany_top_in[1]
port 98 nsew
rlabel metal2 s 6458 22000 6514 22800 4 chany_top_in[2]
port 99 nsew
rlabel metal2 s 6918 22000 6974 22800 4 chany_top_in[3]
port 100 nsew
rlabel metal2 s 7378 22000 7434 22800 4 chany_top_in[4]
port 101 nsew
rlabel metal2 s 7746 22000 7802 22800 4 chany_top_in[5]
port 102 nsew
rlabel metal2 s 8206 22000 8262 22800 4 chany_top_in[6]
port 103 nsew
rlabel metal2 s 8574 22000 8630 22800 4 chany_top_in[7]
port 104 nsew
rlabel metal2 s 9034 22000 9090 22800 4 chany_top_in[8]
port 105 nsew
rlabel metal2 s 9494 22000 9550 22800 4 chany_top_in[9]
port 106 nsew
rlabel metal2 s 14094 22000 14150 22800 4 chany_top_out[0]
port 107 nsew
rlabel metal2 s 18326 22000 18382 22800 4 chany_top_out[10]
port 108 nsew
rlabel metal2 s 18786 22000 18842 22800 4 chany_top_out[11]
port 109 nsew
rlabel metal2 s 19154 22000 19210 22800 4 chany_top_out[12]
port 110 nsew
rlabel metal2 s 19614 22000 19670 22800 4 chany_top_out[13]
port 111 nsew
rlabel metal2 s 19982 22000 20038 22800 4 chany_top_out[14]
port 112 nsew
rlabel metal2 s 20442 22000 20498 22800 4 chany_top_out[15]
port 113 nsew
rlabel metal2 s 20902 22000 20958 22800 4 chany_top_out[16]
port 114 nsew
rlabel metal2 s 21270 22000 21326 22800 4 chany_top_out[17]
port 115 nsew
rlabel metal2 s 21730 22000 21786 22800 4 chany_top_out[18]
port 116 nsew
rlabel metal2 s 22098 22000 22154 22800 4 chany_top_out[19]
port 117 nsew
rlabel metal2 s 14554 22000 14610 22800 4 chany_top_out[1]
port 118 nsew
rlabel metal2 s 14922 22000 14978 22800 4 chany_top_out[2]
port 119 nsew
rlabel metal2 s 15382 22000 15438 22800 4 chany_top_out[3]
port 120 nsew
rlabel metal2 s 15750 22000 15806 22800 4 chany_top_out[4]
port 121 nsew
rlabel metal2 s 16210 22000 16266 22800 4 chany_top_out[5]
port 122 nsew
rlabel metal2 s 16670 22000 16726 22800 4 chany_top_out[6]
port 123 nsew
rlabel metal2 s 17038 22000 17094 22800 4 chany_top_out[7]
port 124 nsew
rlabel metal2 s 17498 22000 17554 22800 4 chany_top_out[8]
port 125 nsew
rlabel metal2 s 17866 22000 17922 22800 4 chany_top_out[9]
port 126 nsew
rlabel metal2 s 4802 22000 4858 22800 4 clk_3_N_out
port 127 nsew
rlabel metal2 s 15842 0 15898 800 4 clk_3_S_in
port 128 nsew
rlabel metal3 s 0 2456 800 2576 4 left_bottom_grid_pin_11_
port 129 nsew
rlabel metal3 s 0 2864 800 2984 4 left_bottom_grid_pin_13_
port 130 nsew
rlabel metal3 s 0 3408 800 3528 4 left_bottom_grid_pin_15_
port 131 nsew
rlabel metal3 s 0 3816 800 3936 4 left_bottom_grid_pin_17_
port 132 nsew
rlabel metal3 s 0 144 800 264 4 left_bottom_grid_pin_1_
port 133 nsew
rlabel metal3 s 0 552 800 672 4 left_bottom_grid_pin_3_
port 134 nsew
rlabel metal3 s 0 960 800 1080 4 left_bottom_grid_pin_5_
port 135 nsew
rlabel metal3 s 0 1504 800 1624 4 left_bottom_grid_pin_7_
port 136 nsew
rlabel metal3 s 0 1912 800 2032 4 left_bottom_grid_pin_9_
port 137 nsew
rlabel metal2 s 3974 22000 4030 22800 4 prog_clk_0_N_in
port 138 nsew
rlabel metal2 s 5262 22000 5318 22800 4 prog_clk_3_N_out
port 139 nsew
rlabel metal2 s 11334 0 11390 800 4 prog_clk_3_S_in
port 140 nsew
rlabel metal3 s 22000 2456 22800 2576 4 right_bottom_grid_pin_11_
port 141 nsew
rlabel metal3 s 22000 2864 22800 2984 4 right_bottom_grid_pin_13_
port 142 nsew
rlabel metal3 s 22000 3408 22800 3528 4 right_bottom_grid_pin_15_
port 143 nsew
rlabel metal3 s 22000 3816 22800 3936 4 right_bottom_grid_pin_17_
port 144 nsew
rlabel metal3 s 22000 144 22800 264 4 right_bottom_grid_pin_1_
port 145 nsew
rlabel metal3 s 22000 552 22800 672 4 right_bottom_grid_pin_3_
port 146 nsew
rlabel metal3 s 22000 960 22800 1080 4 right_bottom_grid_pin_5_
port 147 nsew
rlabel metal3 s 22000 1504 22800 1624 4 right_bottom_grid_pin_7_
port 148 nsew
rlabel metal3 s 22000 1912 22800 2032 4 right_bottom_grid_pin_9_
port 149 nsew
rlabel metal2 s 570 22000 626 22800 4 top_left_grid_pin_42_
port 150 nsew
rlabel metal2 s 1030 22000 1086 22800 4 top_left_grid_pin_43_
port 151 nsew
rlabel metal2 s 1398 22000 1454 22800 4 top_left_grid_pin_44_
port 152 nsew
rlabel metal2 s 1858 22000 1914 22800 4 top_left_grid_pin_45_
port 153 nsew
rlabel metal2 s 2226 22000 2282 22800 4 top_left_grid_pin_46_
port 154 nsew
rlabel metal2 s 2686 22000 2742 22800 4 top_left_grid_pin_47_
port 155 nsew
rlabel metal2 s 3146 22000 3202 22800 4 top_left_grid_pin_48_
port 156 nsew
rlabel metal2 s 3514 22000 3570 22800 4 top_left_grid_pin_49_
port 157 nsew
rlabel metal4 s 4376 2128 4696 20176 4 VPWR
port 158 nsew
rlabel metal4 s 7808 2128 8128 20176 4 VGND
port 159 nsew
<< properties >>
string FIXED_BBOX 0 0 22800 22800
string GDS_FILE /ef/openfpga/openlane/runs/sb_1__0_/results/magic/sb_1__0_.gds
string GDS_END 1224610
string GDS_START 81916
<< end >>
