magic
tech sky130A
magscale 1 2
timestamp 1609023109
<< locali >>
rect 3709 11543 3743 11713
rect 4997 10115 5031 10217
rect 3433 7395 3467 7497
rect 17601 4471 17635 4641
<< viali >>
rect 7205 14501 7239 14535
rect 15945 14501 15979 14535
rect 16865 14501 16899 14535
rect 6929 14433 6963 14467
rect 15853 14365 15887 14399
rect 16957 14365 16991 14399
rect 5917 14025 5951 14059
rect 6837 14025 6871 14059
rect 17693 14025 17727 14059
rect 8861 13957 8895 13991
rect 17325 13957 17359 13991
rect 6469 13889 6503 13923
rect 14013 13889 14047 13923
rect 16865 13889 16899 13923
rect 7113 13821 7147 13855
rect 7380 13821 7414 13855
rect 8585 13821 8619 13855
rect 13093 13821 13127 13855
rect 13277 13821 13311 13855
rect 13645 13821 13679 13855
rect 15704 13821 15738 13855
rect 17141 13821 17175 13855
rect 18061 13821 18095 13855
rect 18429 13821 18463 13855
rect 16037 13753 16071 13787
rect 16129 13753 16163 13787
rect 6285 13685 6319 13719
rect 6377 13685 6411 13719
rect 8493 13685 8527 13719
rect 15807 13685 15841 13719
rect 17601 13685 17635 13719
rect 18245 13685 18279 13719
rect 6101 13481 6135 13515
rect 6561 13481 6595 13515
rect 6929 13481 6963 13515
rect 7757 13481 7791 13515
rect 8217 13481 8251 13515
rect 8585 13481 8619 13515
rect 14473 13481 14507 13515
rect 6469 13413 6503 13447
rect 9505 13413 9539 13447
rect 4896 13345 4930 13379
rect 7297 13345 7331 13379
rect 7389 13345 7423 13379
rect 8125 13345 8159 13379
rect 8953 13345 8987 13379
rect 13360 13345 13394 13379
rect 4629 13277 4663 13311
rect 6653 13277 6687 13311
rect 7481 13277 7515 13311
rect 8309 13277 8343 13311
rect 9045 13277 9079 13311
rect 9137 13277 9171 13311
rect 13093 13277 13127 13311
rect 14565 13277 14599 13311
rect 6009 13141 6043 13175
rect 5733 12937 5767 12971
rect 5917 12937 5951 12971
rect 15853 12937 15887 12971
rect 16957 12937 16991 12971
rect 12817 12869 12851 12903
rect 6469 12801 6503 12835
rect 7389 12801 7423 12835
rect 13461 12801 13495 12835
rect 14289 12801 14323 12835
rect 14473 12801 14507 12835
rect 16773 12801 16807 12835
rect 17693 12801 17727 12835
rect 4353 12733 4387 12767
rect 7849 12733 7883 12767
rect 8116 12733 8150 12767
rect 13277 12733 13311 12767
rect 16497 12733 16531 12767
rect 17601 12733 17635 12767
rect 4620 12665 4654 12699
rect 7205 12665 7239 12699
rect 13185 12665 13219 12699
rect 14740 12665 14774 12699
rect 16589 12665 16623 12699
rect 6285 12597 6319 12631
rect 6377 12597 6411 12631
rect 6837 12597 6871 12631
rect 7297 12597 7331 12631
rect 7665 12597 7699 12631
rect 9229 12597 9263 12631
rect 13645 12597 13679 12631
rect 14013 12597 14047 12631
rect 14105 12597 14139 12631
rect 15945 12597 15979 12631
rect 16129 12597 16163 12631
rect 17141 12597 17175 12631
rect 17509 12597 17543 12631
rect 18061 12597 18095 12631
rect 5733 12393 5767 12427
rect 6193 12393 6227 12427
rect 6561 12393 6595 12427
rect 7389 12393 7423 12427
rect 10149 12393 10183 12427
rect 10701 12393 10735 12427
rect 14289 12393 14323 12427
rect 15485 12393 15519 12427
rect 15853 12393 15887 12427
rect 17693 12393 17727 12427
rect 4344 12325 4378 12359
rect 7021 12325 7055 12359
rect 8217 12325 8251 12359
rect 8585 12325 8619 12359
rect 12992 12325 13026 12359
rect 6101 12257 6135 12291
rect 6929 12257 6963 12291
rect 7757 12257 7791 12291
rect 9137 12257 9171 12291
rect 10609 12257 10643 12291
rect 14657 12257 14691 12291
rect 16313 12257 16347 12291
rect 16580 12257 16614 12291
rect 18153 12257 18187 12291
rect 2145 12189 2179 12223
rect 4077 12189 4111 12223
rect 5641 12189 5675 12223
rect 6285 12189 6319 12223
rect 7205 12189 7239 12223
rect 7849 12189 7883 12223
rect 8033 12189 8067 12223
rect 9229 12189 9263 12223
rect 9321 12189 9355 12223
rect 10885 12189 10919 12223
rect 12725 12189 12759 12223
rect 14749 12189 14783 12223
rect 14933 12189 14967 12223
rect 15945 12189 15979 12223
rect 16129 12189 16163 12223
rect 18245 12189 18279 12223
rect 18337 12189 18371 12223
rect 14105 12121 14139 12155
rect 15393 12121 15427 12155
rect 5457 12053 5491 12087
rect 8769 12053 8803 12087
rect 10241 12053 10275 12087
rect 11161 12053 11195 12087
rect 17785 12053 17819 12087
rect 3617 11849 3651 11883
rect 11253 11849 11287 11883
rect 14289 11849 14323 11883
rect 15209 11849 15243 11883
rect 16037 11849 16071 11883
rect 17785 11849 17819 11883
rect 18429 11849 18463 11883
rect 7113 11781 7147 11815
rect 10333 11781 10367 11815
rect 14105 11781 14139 11815
rect 16865 11781 16899 11815
rect 2053 11713 2087 11747
rect 2881 11713 2915 11747
rect 3709 11713 3743 11747
rect 7021 11713 7055 11747
rect 7849 11713 7883 11747
rect 8033 11713 8067 11747
rect 10977 11713 11011 11747
rect 11805 11713 11839 11747
rect 12633 11713 12667 11747
rect 13277 11713 13311 11747
rect 14013 11713 14047 11747
rect 14749 11713 14783 11747
rect 14933 11713 14967 11747
rect 15853 11713 15887 11747
rect 16681 11713 16715 11747
rect 17509 11713 17543 11747
rect 2605 11577 2639 11611
rect 3341 11577 3375 11611
rect 3801 11645 3835 11679
rect 4068 11645 4102 11679
rect 7297 11645 7331 11679
rect 8953 11645 8987 11679
rect 11621 11645 11655 11679
rect 12173 11645 12207 11679
rect 14657 11645 14691 11679
rect 15669 11645 15703 11679
rect 6653 11577 6687 11611
rect 7757 11577 7791 11611
rect 8309 11577 8343 11611
rect 9220 11577 9254 11611
rect 11713 11577 11747 11611
rect 13093 11577 13127 11611
rect 16405 11577 16439 11611
rect 1409 11509 1443 11543
rect 1777 11509 1811 11543
rect 1869 11509 1903 11543
rect 2237 11509 2271 11543
rect 2697 11509 2731 11543
rect 3065 11509 3099 11543
rect 3709 11509 3743 11543
rect 5181 11509 5215 11543
rect 6377 11509 6411 11543
rect 7389 11509 7423 11543
rect 10425 11509 10459 11543
rect 10793 11509 10827 11543
rect 10885 11509 10919 11543
rect 12725 11509 12759 11543
rect 13185 11509 13219 11543
rect 13645 11509 13679 11543
rect 15577 11509 15611 11543
rect 16497 11509 16531 11543
rect 17233 11509 17267 11543
rect 17325 11509 17359 11543
rect 3525 11305 3559 11339
rect 6837 11305 6871 11339
rect 9137 11305 9171 11339
rect 10057 11305 10091 11339
rect 10609 11305 10643 11339
rect 11069 11305 11103 11339
rect 11161 11305 11195 11339
rect 13277 11305 13311 11339
rect 13645 11305 13679 11339
rect 14105 11305 14139 11339
rect 14565 11305 14599 11339
rect 14933 11305 14967 11339
rect 16865 11305 16899 11339
rect 17509 11305 17543 11339
rect 17969 11305 18003 11339
rect 18429 11305 18463 11339
rect 2412 11237 2446 11271
rect 8002 11237 8036 11271
rect 2053 11169 2087 11203
rect 3801 11169 3835 11203
rect 5724 11169 5758 11203
rect 7297 11169 7331 11203
rect 7757 11169 7791 11203
rect 10517 11169 10551 11203
rect 11888 11169 11922 11203
rect 14473 11169 14507 11203
rect 15117 11169 15151 11203
rect 15741 11169 15775 11203
rect 16957 11169 16991 11203
rect 17877 11169 17911 11203
rect 2145 11101 2179 11135
rect 4077 11101 4111 11135
rect 4997 11101 5031 11135
rect 5457 11101 5491 11135
rect 7389 11101 7423 11135
rect 7481 11101 7515 11135
rect 10701 11101 10735 11135
rect 11621 11101 11655 11135
rect 13093 11101 13127 11135
rect 13737 11101 13771 11135
rect 13829 11101 13863 11135
rect 14657 11101 14691 11135
rect 15485 11101 15519 11135
rect 18061 11101 18095 11135
rect 1869 11033 1903 11067
rect 5273 11033 5307 11067
rect 6929 11033 6963 11067
rect 10149 11033 10183 11067
rect 13001 11033 13035 11067
rect 15393 11033 15427 11067
rect 3617 10965 3651 10999
rect 4353 10965 4387 10999
rect 4537 10965 4571 10999
rect 4905 10965 4939 10999
rect 2237 10761 2271 10795
rect 6193 10761 6227 10795
rect 6837 10761 6871 10795
rect 8861 10761 8895 10795
rect 8953 10761 8987 10795
rect 17509 10761 17543 10795
rect 6285 10693 6319 10727
rect 8493 10693 8527 10727
rect 2053 10625 2087 10659
rect 2697 10625 2731 10659
rect 2881 10625 2915 10659
rect 3801 10625 3835 10659
rect 4629 10625 4663 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 8217 10625 8251 10659
rect 9413 10625 9447 10659
rect 9597 10625 9631 10659
rect 12173 10625 12207 10659
rect 13921 10625 13955 10659
rect 1777 10557 1811 10591
rect 2605 10557 2639 10591
rect 4353 10557 4387 10591
rect 4813 10557 4847 10591
rect 6469 10557 6503 10591
rect 8033 10557 8067 10591
rect 9321 10557 9355 10591
rect 9781 10557 9815 10591
rect 11437 10557 11471 10591
rect 11897 10557 11931 10591
rect 12449 10557 12483 10591
rect 12716 10557 12750 10591
rect 14473 10557 14507 10591
rect 16129 10557 16163 10591
rect 1869 10489 1903 10523
rect 5080 10489 5114 10523
rect 8125 10489 8159 10523
rect 10048 10489 10082 10523
rect 14197 10489 14231 10523
rect 14740 10489 14774 10523
rect 16396 10489 16430 10523
rect 1409 10421 1443 10455
rect 3157 10421 3191 10455
rect 3525 10421 3559 10455
rect 3617 10421 3651 10455
rect 3985 10421 4019 10455
rect 4445 10421 4479 10455
rect 6561 10421 6595 10455
rect 7205 10421 7239 10455
rect 7665 10421 7699 10455
rect 11161 10421 11195 10455
rect 11253 10421 11287 10455
rect 11529 10421 11563 10455
rect 11989 10421 12023 10455
rect 13829 10421 13863 10455
rect 15853 10421 15887 10455
rect 16037 10421 16071 10455
rect 2789 10217 2823 10251
rect 3525 10217 3559 10251
rect 4169 10217 4203 10251
rect 4997 10217 5031 10251
rect 5089 10217 5123 10251
rect 5457 10217 5491 10251
rect 5917 10217 5951 10251
rect 6377 10217 6411 10251
rect 6929 10217 6963 10251
rect 7849 10217 7883 10251
rect 10333 10217 10367 10251
rect 10793 10217 10827 10251
rect 11621 10217 11655 10251
rect 11989 10217 12023 10251
rect 12909 10217 12943 10251
rect 15853 10217 15887 10251
rect 16221 10217 16255 10251
rect 16589 10217 16623 10251
rect 17325 10217 17359 10251
rect 17785 10217 17819 10251
rect 18153 10217 18187 10251
rect 1676 10149 1710 10183
rect 4537 10149 4571 10183
rect 6285 10149 6319 10183
rect 8208 10149 8242 10183
rect 13614 10149 13648 10183
rect 18429 10149 18463 10183
rect 2973 10081 3007 10115
rect 4997 10081 5031 10115
rect 7297 10081 7331 10115
rect 7941 10081 7975 10115
rect 9413 10081 9447 10115
rect 9965 10081 9999 10115
rect 10701 10081 10735 10115
rect 11529 10081 11563 10115
rect 12357 10081 12391 10115
rect 12449 10081 12483 10115
rect 13093 10081 13127 10115
rect 14933 10081 14967 10115
rect 15761 10081 15795 10115
rect 17693 10081 17727 10115
rect 1409 10013 1443 10047
rect 3617 10013 3651 10047
rect 3801 10013 3835 10047
rect 4629 10013 4663 10047
rect 4721 10013 4755 10047
rect 5549 10013 5583 10047
rect 5733 10013 5767 10047
rect 6561 10013 6595 10047
rect 7389 10013 7423 10047
rect 7573 10013 7607 10047
rect 10057 10013 10091 10047
rect 10977 10013 11011 10047
rect 11805 10013 11839 10047
rect 12541 10013 12575 10047
rect 13277 10013 13311 10047
rect 13369 10013 13403 10047
rect 16037 10013 16071 10047
rect 16681 10013 16715 10047
rect 16865 10013 16899 10047
rect 17877 10013 17911 10047
rect 11161 9945 11195 9979
rect 17141 9945 17175 9979
rect 3157 9877 3191 9911
rect 6745 9877 6779 9911
rect 9321 9877 9355 9911
rect 14749 9877 14783 9911
rect 15393 9877 15427 9911
rect 4813 9673 4847 9707
rect 15853 9673 15887 9707
rect 16681 9673 16715 9707
rect 4905 9605 4939 9639
rect 5917 9605 5951 9639
rect 11437 9605 11471 9639
rect 11529 9605 11563 9639
rect 13829 9605 13863 9639
rect 1961 9537 1995 9571
rect 5457 9537 5491 9571
rect 5825 9537 5859 9571
rect 6561 9537 6595 9571
rect 7481 9537 7515 9571
rect 8033 9537 8067 9571
rect 8861 9537 8895 9571
rect 9597 9537 9631 9571
rect 12081 9537 12115 9571
rect 16497 9537 16531 9571
rect 17233 9537 17267 9571
rect 1501 9469 1535 9503
rect 1593 9469 1627 9503
rect 2217 9469 2251 9503
rect 3433 9469 3467 9503
rect 7205 9469 7239 9503
rect 9413 9469 9447 9503
rect 9873 9469 9907 9503
rect 12449 9469 12483 9503
rect 12716 9469 12750 9503
rect 14197 9469 14231 9503
rect 14464 9469 14498 9503
rect 16313 9469 16347 9503
rect 18061 9469 18095 9503
rect 3678 9401 3712 9435
rect 5273 9401 5307 9435
rect 7297 9401 7331 9435
rect 8585 9401 8619 9435
rect 10140 9401 10174 9435
rect 11897 9401 11931 9435
rect 14013 9401 14047 9435
rect 17049 9401 17083 9435
rect 1777 9333 1811 9367
rect 3341 9333 3375 9367
rect 5365 9333 5399 9367
rect 6285 9333 6319 9367
rect 6377 9333 6411 9367
rect 6837 9333 6871 9367
rect 7665 9333 7699 9367
rect 8217 9333 8251 9367
rect 8677 9333 8711 9367
rect 9045 9333 9079 9367
rect 9505 9333 9539 9367
rect 11253 9333 11287 9367
rect 11989 9333 12023 9367
rect 15577 9333 15611 9367
rect 15761 9333 15795 9367
rect 16221 9333 16255 9367
rect 17141 9333 17175 9367
rect 17509 9333 17543 9367
rect 17785 9333 17819 9367
rect 2605 9129 2639 9163
rect 2973 9129 3007 9163
rect 3341 9129 3375 9163
rect 3433 9129 3467 9163
rect 4169 9129 4203 9163
rect 4537 9129 4571 9163
rect 4905 9129 4939 9163
rect 4997 9129 5031 9163
rect 8953 9129 8987 9163
rect 9045 9129 9079 9163
rect 11989 9129 12023 9163
rect 12357 9129 12391 9163
rect 15761 9129 15795 9163
rect 17969 9129 18003 9163
rect 1593 9061 1627 9095
rect 2513 9061 2547 9095
rect 4445 9061 4479 9095
rect 7104 9061 7138 9095
rect 9934 9061 9968 9095
rect 13277 9061 13311 9095
rect 15669 9061 15703 9095
rect 16856 9061 16890 9095
rect 1685 8993 1719 9027
rect 5365 8993 5399 9027
rect 5632 8993 5666 9027
rect 9413 8993 9447 9027
rect 9689 8993 9723 9027
rect 11529 8993 11563 9027
rect 13185 8993 13219 9027
rect 14749 8993 14783 9027
rect 16589 8993 16623 9027
rect 18061 8993 18095 9027
rect 18429 8993 18463 9027
rect 2697 8925 2731 8959
rect 3525 8925 3559 8959
rect 5181 8925 5215 8959
rect 6837 8925 6871 8959
rect 8309 8925 8343 8959
rect 9229 8925 9263 8959
rect 11621 8925 11655 8959
rect 11713 8925 11747 8959
rect 12449 8925 12483 8959
rect 12633 8925 12667 8959
rect 13369 8925 13403 8959
rect 14289 8925 14323 8959
rect 14841 8925 14875 8959
rect 14933 8925 14967 8959
rect 15853 8925 15887 8959
rect 6745 8857 6779 8891
rect 8217 8857 8251 8891
rect 14013 8857 14047 8891
rect 16313 8857 16347 8891
rect 1869 8789 1903 8823
rect 2145 8789 2179 8823
rect 3801 8789 3835 8823
rect 8585 8789 8619 8823
rect 11069 8789 11103 8823
rect 11161 8789 11195 8823
rect 12817 8789 12851 8823
rect 13645 8789 13679 8823
rect 14381 8789 14415 8823
rect 15301 8789 15335 8823
rect 16221 8789 16255 8823
rect 18245 8789 18279 8823
rect 2973 8585 3007 8619
rect 6101 8585 6135 8619
rect 10333 8585 10367 8619
rect 11989 8585 12023 8619
rect 17233 8585 17267 8619
rect 4169 8517 4203 8551
rect 6469 8517 6503 8551
rect 11161 8517 11195 8551
rect 12449 8517 12483 8551
rect 14105 8517 14139 8551
rect 14933 8517 14967 8551
rect 18245 8517 18279 8551
rect 1409 8449 1443 8483
rect 3709 8449 3743 8483
rect 4629 8449 4663 8483
rect 7021 8449 7055 8483
rect 7573 8449 7607 8483
rect 11713 8449 11747 8483
rect 13093 8449 13127 8483
rect 13737 8449 13771 8483
rect 13921 8449 13955 8483
rect 14565 8449 14599 8483
rect 14749 8449 14783 8483
rect 15485 8449 15519 8483
rect 3617 8381 3651 8415
rect 3985 8381 4019 8415
rect 4896 8381 4930 8415
rect 6653 8381 6687 8415
rect 7829 8381 7863 8415
rect 12173 8381 12207 8415
rect 15853 8381 15887 8415
rect 18061 8381 18095 8415
rect 18429 8381 18463 8415
rect 1676 8313 1710 8347
rect 6837 8313 6871 8347
rect 7481 8313 7515 8347
rect 9045 8313 9079 8347
rect 11069 8313 11103 8347
rect 12817 8313 12851 8347
rect 13645 8313 13679 8347
rect 15301 8313 15335 8347
rect 15393 8313 15427 8347
rect 16098 8313 16132 8347
rect 2789 8245 2823 8279
rect 3157 8245 3191 8279
rect 3525 8245 3559 8279
rect 4353 8245 4387 8279
rect 6009 8245 6043 8279
rect 6285 8245 6319 8279
rect 7297 8245 7331 8279
rect 8953 8245 8987 8279
rect 11529 8245 11563 8279
rect 11621 8245 11655 8279
rect 12909 8245 12943 8279
rect 13277 8245 13311 8279
rect 14473 8245 14507 8279
rect 2329 8041 2363 8075
rect 2421 8041 2455 8075
rect 2789 8041 2823 8075
rect 3249 8041 3283 8075
rect 3801 8041 3835 8075
rect 4445 8041 4479 8075
rect 5181 8041 5215 8075
rect 5365 8041 5399 8075
rect 5549 8041 5583 8075
rect 8677 8041 8711 8075
rect 9689 8041 9723 8075
rect 10057 8041 10091 8075
rect 10517 8041 10551 8075
rect 10885 8041 10919 8075
rect 10977 8041 11011 8075
rect 12725 8041 12759 8075
rect 16681 8041 16715 8075
rect 1501 7973 1535 8007
rect 6469 7973 6503 8007
rect 7849 7973 7883 8007
rect 9137 7973 9171 8007
rect 11590 7973 11624 8007
rect 17693 7973 17727 8007
rect 1593 7905 1627 7939
rect 3157 7905 3191 7939
rect 3617 7905 3651 7939
rect 4537 7905 4571 7939
rect 5917 7905 5951 7939
rect 6929 7905 6963 7939
rect 7021 7905 7055 7939
rect 7757 7905 7791 7939
rect 8585 7905 8619 7939
rect 10149 7905 10183 7939
rect 13277 7905 13311 7939
rect 13544 7905 13578 7939
rect 15568 7905 15602 7939
rect 17877 7905 17911 7939
rect 2605 7837 2639 7871
rect 3433 7837 3467 7871
rect 4629 7837 4663 7871
rect 6009 7837 6043 7871
rect 6101 7837 6135 7871
rect 7205 7837 7239 7871
rect 7941 7837 7975 7871
rect 8769 7837 8803 7871
rect 10333 7837 10367 7871
rect 11069 7837 11103 7871
rect 11345 7837 11379 7871
rect 12817 7837 12851 7871
rect 15301 7837 15335 7871
rect 7389 7769 7423 7803
rect 14657 7769 14691 7803
rect 18061 7769 18095 7803
rect 1777 7701 1811 7735
rect 1961 7701 1995 7735
rect 4077 7701 4111 7735
rect 4997 7701 5031 7735
rect 6561 7701 6595 7735
rect 8217 7701 8251 7735
rect 9413 7701 9447 7735
rect 13185 7701 13219 7735
rect 14749 7701 14783 7735
rect 14933 7701 14967 7735
rect 3433 7497 3467 7531
rect 6285 7497 6319 7531
rect 6837 7497 6871 7531
rect 10701 7497 10735 7531
rect 12449 7497 12483 7531
rect 14197 7497 14231 7531
rect 15853 7497 15887 7531
rect 16681 7497 16715 7531
rect 1501 7429 1535 7463
rect 9873 7429 9907 7463
rect 18245 7429 18279 7463
rect 3433 7361 3467 7395
rect 4077 7361 4111 7395
rect 4905 7361 4939 7395
rect 6469 7361 6503 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 7665 7361 7699 7395
rect 10425 7361 10459 7395
rect 11161 7361 11195 7395
rect 11253 7361 11287 7395
rect 12127 7361 12161 7395
rect 13093 7361 13127 7395
rect 13921 7361 13955 7395
rect 14657 7361 14691 7395
rect 14841 7361 14875 7395
rect 15577 7361 15611 7395
rect 16313 7361 16347 7395
rect 16405 7361 16439 7395
rect 1593 7293 1627 7327
rect 3065 7293 3099 7327
rect 3893 7293 3927 7327
rect 4353 7293 4387 7327
rect 6653 7293 6687 7327
rect 7205 7293 7239 7327
rect 8125 7293 8159 7327
rect 8392 7293 8426 7327
rect 10241 7293 10275 7327
rect 11897 7293 11931 7327
rect 12817 7293 12851 7327
rect 13829 7293 13863 7327
rect 15485 7293 15519 7327
rect 18061 7293 18095 7327
rect 18429 7293 18463 7327
rect 1860 7225 1894 7259
rect 3985 7225 4019 7259
rect 5172 7225 5206 7259
rect 13737 7225 13771 7259
rect 16221 7225 16255 7259
rect 2973 7157 3007 7191
rect 3249 7157 3283 7191
rect 3525 7157 3559 7191
rect 4537 7157 4571 7191
rect 4813 7157 4847 7191
rect 8033 7157 8067 7191
rect 9505 7157 9539 7191
rect 9781 7157 9815 7191
rect 10333 7157 10367 7191
rect 11069 7157 11103 7191
rect 11529 7157 11563 7191
rect 11989 7157 12023 7191
rect 12909 7157 12943 7191
rect 13369 7157 13403 7191
rect 14565 7157 14599 7191
rect 15025 7157 15059 7191
rect 15393 7157 15427 7191
rect 2053 6953 2087 6987
rect 4537 6953 4571 6987
rect 5641 6953 5675 6987
rect 6101 6953 6135 6987
rect 11529 6953 11563 6987
rect 12081 6953 12115 6987
rect 12633 6953 12667 6987
rect 12725 6953 12759 6987
rect 13093 6953 13127 6987
rect 13921 6953 13955 6987
rect 15485 6953 15519 6987
rect 15853 6953 15887 6987
rect 2145 6885 2179 6919
rect 5733 6885 5767 6919
rect 11713 6885 11747 6919
rect 13461 6885 13495 6919
rect 14289 6885 14323 6919
rect 17601 6885 17635 6919
rect 2780 6817 2814 6851
rect 4445 6817 4479 6851
rect 5181 6817 5215 6851
rect 6469 6817 6503 6851
rect 6929 6817 6963 6851
rect 7196 6817 7230 6851
rect 9137 6817 9171 6851
rect 9873 6817 9907 6851
rect 10149 6817 10183 6851
rect 10416 6817 10450 6851
rect 17877 6817 17911 6851
rect 18245 6817 18279 6851
rect 2329 6749 2363 6783
rect 2513 6749 2547 6783
rect 4629 6749 4663 6783
rect 5917 6749 5951 6783
rect 6561 6749 6595 6783
rect 6745 6749 6779 6783
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 12909 6749 12943 6783
rect 13553 6749 13587 6783
rect 13737 6749 13771 6783
rect 14381 6749 14415 6783
rect 14473 6749 14507 6783
rect 14933 6749 14967 6783
rect 15301 6749 15335 6783
rect 1593 6681 1627 6715
rect 3893 6681 3927 6715
rect 5273 6681 5307 6715
rect 8309 6681 8343 6715
rect 8677 6681 8711 6715
rect 14841 6681 14875 6715
rect 18429 6681 18463 6715
rect 1685 6613 1719 6647
rect 4077 6613 4111 6647
rect 4997 6613 5031 6647
rect 8401 6613 8435 6647
rect 8769 6613 8803 6647
rect 9781 6613 9815 6647
rect 11897 6613 11931 6647
rect 12265 6613 12299 6647
rect 17693 6613 17727 6647
rect 18061 6613 18095 6647
rect 2789 6409 2823 6443
rect 3617 6409 3651 6443
rect 5457 6409 5491 6443
rect 5917 6409 5951 6443
rect 8217 6409 8251 6443
rect 10241 6409 10275 6443
rect 10517 6409 10551 6443
rect 12817 6409 12851 6443
rect 13185 6409 13219 6443
rect 15393 6409 15427 6443
rect 2237 6341 2271 6375
rect 15485 6341 15519 6375
rect 1501 6273 1535 6307
rect 3433 6273 3467 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 6837 6273 6871 6307
rect 13829 6273 13863 6307
rect 1685 6205 1719 6239
rect 2053 6205 2087 6239
rect 2421 6205 2455 6239
rect 3157 6205 3191 6239
rect 3801 6205 3835 6239
rect 4068 6205 4102 6239
rect 5273 6205 5307 6239
rect 5825 6205 5859 6239
rect 6285 6205 6319 6239
rect 7104 6205 7138 6239
rect 8769 6205 8803 6239
rect 10885 6205 10919 6239
rect 11152 6205 11186 6239
rect 12633 6205 12667 6239
rect 14013 6205 14047 6239
rect 14269 6205 14303 6239
rect 18061 6205 18095 6239
rect 18429 6205 18463 6239
rect 3249 6137 3283 6171
rect 8401 6137 8435 6171
rect 9036 6137 9070 6171
rect 13553 6137 13587 6171
rect 1869 6069 1903 6103
rect 2605 6069 2639 6103
rect 5181 6069 5215 6103
rect 5641 6069 5675 6103
rect 8585 6069 8619 6103
rect 10149 6069 10183 6103
rect 10701 6069 10735 6103
rect 12265 6069 12299 6103
rect 12449 6069 12483 6103
rect 13093 6069 13127 6103
rect 13645 6069 13679 6103
rect 18245 6069 18279 6103
rect 3617 5865 3651 5899
rect 4077 5865 4111 5899
rect 4537 5865 4571 5899
rect 9321 5865 9355 5899
rect 11345 5865 11379 5899
rect 11805 5865 11839 5899
rect 12173 5865 12207 5899
rect 12265 5865 12299 5899
rect 14013 5865 14047 5899
rect 17693 5865 17727 5899
rect 1768 5797 1802 5831
rect 7205 5797 7239 5831
rect 1501 5729 1535 5763
rect 3525 5729 3559 5763
rect 4445 5729 4479 5763
rect 4905 5729 4939 5763
rect 5365 5729 5399 5763
rect 5632 5729 5666 5763
rect 7849 5729 7883 5763
rect 8585 5729 8619 5763
rect 9045 5729 9079 5763
rect 9505 5729 9539 5763
rect 9873 5729 9907 5763
rect 10140 5729 10174 5763
rect 12633 5729 12667 5763
rect 12889 5729 12923 5763
rect 14473 5729 14507 5763
rect 14933 5729 14967 5763
rect 17877 5729 17911 5763
rect 18245 5729 18279 5763
rect 3709 5661 3743 5695
rect 4629 5661 4663 5695
rect 7297 5661 7331 5695
rect 7389 5661 7423 5695
rect 8677 5661 8711 5695
rect 8769 5661 8803 5695
rect 11621 5661 11655 5695
rect 12357 5661 12391 5695
rect 14565 5661 14599 5695
rect 14749 5661 14783 5695
rect 2973 5593 3007 5627
rect 6745 5593 6779 5627
rect 7941 5593 7975 5627
rect 15301 5593 15335 5627
rect 18429 5593 18463 5627
rect 2881 5525 2915 5559
rect 3157 5525 3191 5559
rect 5089 5525 5123 5559
rect 6837 5525 6871 5559
rect 7665 5525 7699 5559
rect 8217 5525 8251 5559
rect 9781 5525 9815 5559
rect 11253 5525 11287 5559
rect 14105 5525 14139 5559
rect 18061 5525 18095 5559
rect 3065 5321 3099 5355
rect 3985 5321 4019 5355
rect 5917 5321 5951 5355
rect 9229 5321 9263 5355
rect 10885 5321 10919 5355
rect 13829 5321 13863 5355
rect 18061 5321 18095 5355
rect 4813 5253 4847 5287
rect 8309 5253 8343 5287
rect 8401 5253 8435 5287
rect 3617 5185 3651 5219
rect 3709 5185 3743 5219
rect 4629 5185 4663 5219
rect 5365 5185 5399 5219
rect 6469 5185 6503 5219
rect 8953 5185 8987 5219
rect 9781 5185 9815 5219
rect 10517 5185 10551 5219
rect 10701 5185 10735 5219
rect 11437 5185 11471 5219
rect 14013 5185 14047 5219
rect 16037 5185 16071 5219
rect 1501 5117 1535 5151
rect 1768 5117 1802 5151
rect 5181 5117 5215 5151
rect 6929 5117 6963 5151
rect 9597 5117 9631 5151
rect 10425 5117 10459 5151
rect 11345 5117 11379 5151
rect 12265 5117 12299 5151
rect 12449 5117 12483 5151
rect 14280 5117 14314 5151
rect 15945 5117 15979 5151
rect 16313 5117 16347 5151
rect 7196 5049 7230 5083
rect 9689 5049 9723 5083
rect 11253 5049 11287 5083
rect 12716 5049 12750 5083
rect 2881 4981 2915 5015
rect 3157 4981 3191 5015
rect 3525 4981 3559 5015
rect 4353 4981 4387 5015
rect 4445 4981 4479 5015
rect 5273 4981 5307 5015
rect 5641 4981 5675 5015
rect 6285 4981 6319 5015
rect 6377 4981 6411 5015
rect 8769 4981 8803 5015
rect 8861 4981 8895 5015
rect 10057 4981 10091 5015
rect 11713 4981 11747 5015
rect 12081 4981 12115 5015
rect 15393 4981 15427 5015
rect 15485 4981 15519 5015
rect 15853 4981 15887 5015
rect 1593 4777 1627 4811
rect 2053 4777 2087 4811
rect 4077 4777 4111 4811
rect 4537 4777 4571 4811
rect 5089 4777 5123 4811
rect 6285 4777 6319 4811
rect 6745 4777 6779 4811
rect 7389 4777 7423 4811
rect 8677 4777 8711 4811
rect 11529 4777 11563 4811
rect 12541 4777 12575 4811
rect 12909 4777 12943 4811
rect 13277 4777 13311 4811
rect 13737 4777 13771 4811
rect 14105 4777 14139 4811
rect 14565 4777 14599 4811
rect 2145 4709 2179 4743
rect 4445 4709 4479 4743
rect 7297 4709 7331 4743
rect 7757 4709 7791 4743
rect 9321 4709 9355 4743
rect 9956 4709 9990 4743
rect 12449 4709 12483 4743
rect 2780 4641 2814 4675
rect 4997 4641 5031 4675
rect 5457 4641 5491 4675
rect 6377 4641 6411 4675
rect 6929 4641 6963 4675
rect 7849 4641 7883 4675
rect 8585 4641 8619 4675
rect 13369 4641 13403 4675
rect 14841 4641 14875 4675
rect 17601 4641 17635 4675
rect 17877 4641 17911 4675
rect 2329 4573 2363 4607
rect 2513 4573 2547 4607
rect 4629 4573 4663 4607
rect 5549 4573 5583 4607
rect 5641 4573 5675 4607
rect 6469 4573 6503 4607
rect 8033 4573 8067 4607
rect 8769 4573 8803 4607
rect 9413 4573 9447 4607
rect 9689 4573 9723 4607
rect 11621 4573 11655 4607
rect 11713 4573 11747 4607
rect 12725 4573 12759 4607
rect 13553 4573 13587 4607
rect 14197 4573 14231 4607
rect 14289 4573 14323 4607
rect 8217 4505 8251 4539
rect 9045 4505 9079 4539
rect 15025 4505 15059 4539
rect 1685 4437 1719 4471
rect 3893 4437 3927 4471
rect 5917 4437 5951 4471
rect 11069 4437 11103 4471
rect 11161 4437 11195 4471
rect 12081 4437 12115 4471
rect 17601 4437 17635 4471
rect 17693 4437 17727 4471
rect 18061 4437 18095 4471
rect 3617 4233 3651 4267
rect 5365 4233 5399 4267
rect 6837 4233 6871 4267
rect 9045 4233 9079 4267
rect 10241 4233 10275 4267
rect 11897 4233 11931 4267
rect 12081 4233 12115 4267
rect 12725 4233 12759 4267
rect 14381 4233 14415 4267
rect 18429 4233 18463 4267
rect 5273 4165 5307 4199
rect 9137 4165 9171 4199
rect 13553 4165 13587 4199
rect 5917 4097 5951 4131
rect 6193 4097 6227 4131
rect 7389 4097 7423 4131
rect 9689 4097 9723 4131
rect 13369 4097 13403 4131
rect 14105 4097 14139 4131
rect 15025 4097 15059 4131
rect 17785 4097 17819 4131
rect 1685 4029 1719 4063
rect 2237 4029 2271 4063
rect 2493 4029 2527 4063
rect 3801 4029 3835 4063
rect 3893 4029 3927 4063
rect 5825 4029 5859 4063
rect 7665 4029 7699 4063
rect 9597 4029 9631 4063
rect 10517 4029 10551 4063
rect 10784 4029 10818 4063
rect 13093 4029 13127 4063
rect 13921 4029 13955 4063
rect 14013 4029 14047 4063
rect 18061 4029 18095 4063
rect 4160 3961 4194 3995
rect 7205 3961 7239 3995
rect 7932 3961 7966 3995
rect 13185 3961 13219 3995
rect 14841 3961 14875 3995
rect 1593 3893 1627 3927
rect 1869 3893 1903 3927
rect 2053 3893 2087 3927
rect 5733 3893 5767 3927
rect 6561 3893 6595 3927
rect 7297 3893 7331 3927
rect 9505 3893 9539 3927
rect 9965 3893 9999 3927
rect 10333 3893 10367 3927
rect 12633 3893 12667 3927
rect 14749 3893 14783 3927
rect 15301 3893 15335 3927
rect 18245 3893 18279 3927
rect 2973 3689 3007 3723
rect 4537 3689 4571 3723
rect 6101 3689 6135 3723
rect 6745 3689 6779 3723
rect 7389 3689 7423 3723
rect 9045 3689 9079 3723
rect 10425 3689 10459 3723
rect 10977 3689 11011 3723
rect 11345 3689 11379 3723
rect 14749 3689 14783 3723
rect 17693 3689 17727 3723
rect 2881 3621 2915 3655
rect 5273 3621 5307 3655
rect 7021 3621 7055 3655
rect 8677 3621 8711 3655
rect 9413 3621 9447 3655
rect 12050 3621 12084 3655
rect 13544 3621 13578 3655
rect 1593 3553 1627 3587
rect 1685 3553 1719 3587
rect 2053 3553 2087 3587
rect 2421 3553 2455 3587
rect 3341 3553 3375 3587
rect 4445 3553 4479 3587
rect 7757 3553 7791 3587
rect 8585 3553 8619 3587
rect 9229 3553 9263 3587
rect 10333 3553 10367 3587
rect 10885 3553 10919 3587
rect 11437 3553 11471 3587
rect 17509 3553 17543 3587
rect 17877 3553 17911 3587
rect 18245 3553 18279 3587
rect 3433 3485 3467 3519
rect 3617 3485 3651 3519
rect 4721 3485 4755 3519
rect 5365 3485 5399 3519
rect 5549 3485 5583 3519
rect 6193 3485 6227 3519
rect 6377 3485 6411 3519
rect 7297 3485 7331 3519
rect 7849 3485 7883 3519
rect 8033 3485 8067 3519
rect 8769 3485 8803 3519
rect 10609 3485 10643 3519
rect 11529 3485 11563 3519
rect 11805 3485 11839 3519
rect 13277 3485 13311 3519
rect 17141 3485 17175 3519
rect 2605 3417 2639 3451
rect 3893 3417 3927 3451
rect 4077 3417 4111 3451
rect 8217 3417 8251 3451
rect 13185 3417 13219 3451
rect 14657 3417 14691 3451
rect 1869 3349 1903 3383
rect 2237 3349 2271 3383
rect 4905 3349 4939 3383
rect 5733 3349 5767 3383
rect 6561 3349 6595 3383
rect 9781 3349 9815 3383
rect 9965 3349 9999 3383
rect 17325 3349 17359 3383
rect 18061 3349 18095 3383
rect 18429 3349 18463 3383
rect 2605 3145 2639 3179
rect 3065 3145 3099 3179
rect 3893 3145 3927 3179
rect 6561 3145 6595 3179
rect 8217 3145 8251 3179
rect 8401 3145 8435 3179
rect 17417 3145 17451 3179
rect 2329 3077 2363 3111
rect 2881 3077 2915 3111
rect 4721 3077 4755 3111
rect 13001 3077 13035 3111
rect 13461 3077 13495 3111
rect 3617 3009 3651 3043
rect 4445 3009 4479 3043
rect 5181 3009 5215 3043
rect 8769 3009 8803 3043
rect 9689 3009 9723 3043
rect 10333 3009 10367 3043
rect 10517 3009 10551 3043
rect 11437 3009 11471 3043
rect 11897 3009 11931 3043
rect 13185 3009 13219 3043
rect 1593 2941 1627 2975
rect 2145 2941 2179 2975
rect 2697 2941 2731 2975
rect 3433 2941 3467 2975
rect 4353 2941 4387 2975
rect 4997 2941 5031 2975
rect 6837 2941 6871 2975
rect 7093 2941 7127 2975
rect 8493 2941 8527 2975
rect 11161 2941 11195 2975
rect 11713 2941 11747 2975
rect 12449 2941 12483 2975
rect 14197 2941 14231 2975
rect 16773 2941 16807 2975
rect 16865 2941 16899 2975
rect 17601 2941 17635 2975
rect 18061 2941 18095 2975
rect 18429 2941 18463 2975
rect 1869 2873 1903 2907
rect 5448 2873 5482 2907
rect 9413 2873 9447 2907
rect 10241 2873 10275 2907
rect 12725 2873 12759 2907
rect 14473 2873 14507 2907
rect 1501 2805 1535 2839
rect 3525 2805 3559 2839
rect 4261 2805 4295 2839
rect 9045 2805 9079 2839
rect 9505 2805 9539 2839
rect 9873 2805 9907 2839
rect 10793 2805 10827 2839
rect 11253 2805 11287 2839
rect 17049 2805 17083 2839
rect 17785 2805 17819 2839
rect 18245 2805 18279 2839
rect 1501 2601 1535 2635
rect 4721 2601 4755 2635
rect 5089 2601 5123 2635
rect 9965 2601 9999 2635
rect 10425 2601 10459 2635
rect 10793 2601 10827 2635
rect 11253 2601 11287 2635
rect 11621 2601 11655 2635
rect 11989 2601 12023 2635
rect 12081 2601 12115 2635
rect 14013 2601 14047 2635
rect 16773 2601 16807 2635
rect 5181 2533 5215 2567
rect 8309 2533 8343 2567
rect 10333 2533 10367 2567
rect 1593 2465 1627 2499
rect 2145 2465 2179 2499
rect 2697 2465 2731 2499
rect 3249 2465 3283 2499
rect 3617 2465 3651 2499
rect 4077 2465 4111 2499
rect 5549 2465 5583 2499
rect 6101 2465 6135 2499
rect 6929 2465 6963 2499
rect 8033 2465 8067 2499
rect 8585 2465 8619 2499
rect 9137 2465 9171 2499
rect 11161 2465 11195 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 14381 2465 14415 2499
rect 16129 2465 16163 2499
rect 17141 2465 17175 2499
rect 17509 2465 17543 2499
rect 17877 2465 17911 2499
rect 18337 2465 18371 2499
rect 1777 2397 1811 2431
rect 2329 2397 2363 2431
rect 2973 2397 3007 2431
rect 4261 2397 4295 2431
rect 5365 2397 5399 2431
rect 5733 2397 5767 2431
rect 6285 2397 6319 2431
rect 7757 2397 7791 2431
rect 8769 2397 8803 2431
rect 9321 2397 9355 2431
rect 10609 2397 10643 2431
rect 11437 2397 11471 2431
rect 12173 2397 12207 2431
rect 12817 2397 12851 2431
rect 13369 2397 13403 2431
rect 14565 2397 14599 2431
rect 17049 2397 17083 2431
rect 3433 2261 3467 2295
rect 3801 2261 3835 2295
rect 6653 2261 6687 2295
rect 9873 2261 9907 2295
rect 13737 2261 13771 2295
rect 16313 2261 16347 2295
rect 17325 2261 17359 2295
rect 17693 2261 17727 2295
rect 18061 2261 18095 2295
<< metal1 >>
rect 3418 15716 3424 15768
rect 3476 15756 3482 15768
rect 6638 15756 6644 15768
rect 3476 15728 6644 15756
rect 3476 15716 3482 15728
rect 6638 15716 6644 15728
rect 6696 15716 6702 15768
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 18046 14600 18052 14612
rect 13320 14572 18052 14600
rect 13320 14560 13326 14572
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 7193 14535 7251 14541
rect 7193 14501 7205 14535
rect 7239 14532 7251 14535
rect 12158 14532 12164 14544
rect 7239 14504 12164 14532
rect 7239 14501 7251 14504
rect 7193 14495 7251 14501
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 14366 14492 14372 14544
rect 14424 14532 14430 14544
rect 15933 14535 15991 14541
rect 15933 14532 15945 14535
rect 14424 14504 15945 14532
rect 14424 14492 14430 14504
rect 15933 14501 15945 14504
rect 15979 14501 15991 14535
rect 15933 14495 15991 14501
rect 16853 14535 16911 14541
rect 16853 14501 16865 14535
rect 16899 14532 16911 14535
rect 18782 14532 18788 14544
rect 16899 14504 18788 14532
rect 16899 14501 16911 14504
rect 16853 14495 16911 14501
rect 18782 14492 18788 14504
rect 18840 14492 18846 14544
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 5960 14436 6929 14464
rect 5960 14424 5966 14436
rect 6917 14433 6929 14436
rect 6963 14433 6975 14467
rect 11422 14464 11428 14476
rect 6917 14427 6975 14433
rect 7024 14436 11428 14464
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 7024 14396 7052 14436
rect 11422 14424 11428 14436
rect 11480 14424 11486 14476
rect 4120 14368 7052 14396
rect 4120 14356 4126 14368
rect 15286 14356 15292 14408
rect 15344 14396 15350 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15344 14368 15853 14396
rect 15344 14356 15350 14368
rect 15841 14365 15853 14368
rect 15887 14396 15899 14399
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 15887 14368 16957 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 3786 14288 3792 14340
rect 3844 14328 3850 14340
rect 8938 14328 8944 14340
rect 3844 14300 8944 14328
rect 3844 14288 3850 14300
rect 8938 14288 8944 14300
rect 8996 14288 9002 14340
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 13262 14260 13268 14272
rect 3384 14232 13268 14260
rect 3384 14220 3390 14232
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 16206 14260 16212 14272
rect 13412 14232 16212 14260
rect 13412 14220 13418 14232
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 5902 14056 5908 14068
rect 5863 14028 5908 14056
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6788 14028 6837 14056
rect 6788 14016 6794 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 16574 14056 16580 14068
rect 6825 14019 6883 14025
rect 16040 14028 16580 14056
rect 16040 14000 16068 14028
rect 16574 14016 16580 14028
rect 16632 14056 16638 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 16632 14028 17693 14056
rect 16632 14016 16638 14028
rect 17681 14025 17693 14028
rect 17727 14025 17739 14059
rect 17681 14019 17739 14025
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 8849 13991 8907 13997
rect 8849 13988 8861 13991
rect 8260 13960 8861 13988
rect 8260 13948 8266 13960
rect 8849 13957 8861 13960
rect 8895 13988 8907 13991
rect 14734 13988 14740 14000
rect 8895 13960 14740 13988
rect 8895 13957 8907 13960
rect 8849 13951 8907 13957
rect 14734 13948 14740 13960
rect 14792 13948 14798 14000
rect 16022 13948 16028 14000
rect 16080 13948 16086 14000
rect 17313 13991 17371 13997
rect 17313 13988 17325 13991
rect 16592 13960 17325 13988
rect 5994 13880 6000 13932
rect 6052 13920 6058 13932
rect 6457 13923 6515 13929
rect 6457 13920 6469 13923
rect 6052 13892 6469 13920
rect 6052 13880 6058 13892
rect 6457 13889 6469 13892
rect 6503 13889 6515 13923
rect 6457 13883 6515 13889
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13920 14059 13923
rect 14366 13920 14372 13932
rect 14047 13892 14372 13920
rect 14047 13889 14059 13892
rect 14001 13883 14059 13889
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 16592 13920 16620 13960
rect 17313 13957 17325 13960
rect 17359 13957 17371 13991
rect 17313 13951 17371 13957
rect 16850 13920 16856 13932
rect 15856 13892 16620 13920
rect 16811 13892 16856 13920
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 7190 13852 7196 13864
rect 7147 13824 7196 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 7368 13855 7426 13861
rect 7368 13821 7380 13855
rect 7414 13852 7426 13855
rect 7742 13852 7748 13864
rect 7414 13824 7748 13852
rect 7414 13821 7426 13824
rect 7368 13815 7426 13821
rect 7742 13812 7748 13824
rect 7800 13852 7806 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 7800 13824 8585 13852
rect 7800 13812 7806 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12768 13824 13093 13852
rect 12768 13812 12774 13824
rect 13081 13821 13093 13824
rect 13127 13852 13139 13855
rect 13265 13855 13323 13861
rect 13265 13852 13277 13855
rect 13127 13824 13277 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 13265 13821 13277 13824
rect 13311 13821 13323 13855
rect 13630 13852 13636 13864
rect 13591 13824 13636 13852
rect 13265 13815 13323 13821
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 14384 13852 14412 13880
rect 15692 13855 15750 13861
rect 15692 13852 15704 13855
rect 14384 13824 15704 13852
rect 15692 13821 15704 13824
rect 15738 13821 15750 13855
rect 15692 13815 15750 13821
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 15856 13784 15884 13892
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 18046 13852 18052 13864
rect 17175 13824 17632 13852
rect 18007 13824 18052 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 16022 13784 16028 13796
rect 5592 13756 15884 13784
rect 15983 13756 16028 13784
rect 5592 13744 5598 13756
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 16117 13787 16175 13793
rect 16117 13753 16129 13787
rect 16163 13753 16175 13787
rect 16117 13747 16175 13753
rect 6086 13676 6092 13728
rect 6144 13716 6150 13728
rect 6273 13719 6331 13725
rect 6273 13716 6285 13719
rect 6144 13688 6285 13716
rect 6144 13676 6150 13688
rect 6273 13685 6285 13688
rect 6319 13685 6331 13719
rect 6273 13679 6331 13685
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6420 13688 6465 13716
rect 6420 13676 6426 13688
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 8481 13719 8539 13725
rect 8481 13716 8493 13719
rect 8444 13688 8493 13716
rect 8444 13676 8450 13688
rect 8481 13685 8493 13688
rect 8527 13685 8539 13719
rect 8481 13679 8539 13685
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 13630 13716 13636 13728
rect 10284 13688 13636 13716
rect 10284 13676 10290 13688
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 15795 13719 15853 13725
rect 15795 13685 15807 13719
rect 15841 13716 15853 13719
rect 16132 13716 16160 13747
rect 17604 13728 17632 13824
rect 18046 13812 18052 13824
rect 18104 13852 18110 13864
rect 18417 13855 18475 13861
rect 18417 13852 18429 13855
rect 18104 13824 18429 13852
rect 18104 13812 18110 13824
rect 18417 13821 18429 13824
rect 18463 13821 18475 13855
rect 18417 13815 18475 13821
rect 17586 13716 17592 13728
rect 15841 13688 16160 13716
rect 17547 13688 17592 13716
rect 15841 13685 15853 13688
rect 15795 13679 15853 13685
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 18233 13719 18291 13725
rect 18233 13685 18245 13719
rect 18279 13716 18291 13719
rect 18506 13716 18512 13728
rect 18279 13688 18512 13716
rect 18279 13685 18291 13688
rect 18233 13679 18291 13685
rect 18506 13676 18512 13688
rect 18564 13676 18570 13728
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 6549 13515 6607 13521
rect 6549 13481 6561 13515
rect 6595 13512 6607 13515
rect 6917 13515 6975 13521
rect 6917 13512 6929 13515
rect 6595 13484 6929 13512
rect 6595 13481 6607 13484
rect 6549 13475 6607 13481
rect 6917 13481 6929 13484
rect 6963 13481 6975 13515
rect 6917 13475 6975 13481
rect 7745 13515 7803 13521
rect 7745 13481 7757 13515
rect 7791 13481 7803 13515
rect 8202 13512 8208 13524
rect 8163 13484 8208 13512
rect 7745 13475 7803 13481
rect 6457 13447 6515 13453
rect 6457 13413 6469 13447
rect 6503 13444 6515 13447
rect 7760 13444 7788 13475
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 8573 13515 8631 13521
rect 8573 13481 8585 13515
rect 8619 13512 8631 13515
rect 11698 13512 11704 13524
rect 8619 13484 11704 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 14461 13515 14519 13521
rect 14461 13512 14473 13515
rect 13688 13484 14473 13512
rect 13688 13472 13694 13484
rect 14461 13481 14473 13484
rect 14507 13481 14519 13515
rect 14461 13475 14519 13481
rect 8662 13444 8668 13456
rect 6503 13416 7788 13444
rect 7944 13416 8668 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 4884 13379 4942 13385
rect 4884 13345 4896 13379
rect 4930 13376 4942 13379
rect 5718 13376 5724 13388
rect 4930 13348 5724 13376
rect 4930 13345 4942 13348
rect 4884 13339 4942 13345
rect 5718 13336 5724 13348
rect 5776 13376 5782 13388
rect 5776 13348 6684 13376
rect 5776 13336 5782 13348
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 6656 13317 6684 13348
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 6880 13348 7297 13376
rect 6880 13336 6886 13348
rect 7285 13345 7297 13348
rect 7331 13345 7343 13379
rect 7285 13339 7343 13345
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13376 7435 13379
rect 7944 13376 7972 13416
rect 8662 13404 8668 13416
rect 8720 13444 8726 13456
rect 9493 13447 9551 13453
rect 9493 13444 9505 13447
rect 8720 13416 9505 13444
rect 8720 13404 8726 13416
rect 9493 13413 9505 13416
rect 9539 13444 9551 13447
rect 13078 13444 13084 13456
rect 9539 13416 13084 13444
rect 9539 13413 9551 13416
rect 9493 13407 9551 13413
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 13170 13404 13176 13456
rect 13228 13444 13234 13456
rect 16942 13444 16948 13456
rect 13228 13416 16948 13444
rect 13228 13404 13234 13416
rect 16942 13404 16948 13416
rect 17000 13404 17006 13456
rect 8110 13376 8116 13388
rect 7423 13348 7972 13376
rect 8071 13348 8116 13376
rect 7423 13345 7435 13348
rect 7377 13339 7435 13345
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13376 8999 13379
rect 10778 13376 10784 13388
rect 8987 13348 10784 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 13348 13379 13406 13385
rect 13348 13345 13360 13379
rect 13394 13376 13406 13379
rect 13814 13376 13820 13388
rect 13394 13348 13820 13376
rect 13394 13345 13406 13348
rect 13348 13339 13406 13345
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 4396 13280 4629 13308
rect 4396 13268 4402 13280
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 6788 13280 7481 13308
rect 6788 13268 6794 13280
rect 7469 13277 7481 13280
rect 7515 13308 7527 13311
rect 8297 13311 8355 13317
rect 8297 13308 8309 13311
rect 7515 13280 8309 13308
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 8297 13277 8309 13280
rect 8343 13277 8355 13311
rect 8297 13271 8355 13277
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 9033 13311 9091 13317
rect 9033 13308 9045 13311
rect 8628 13280 9045 13308
rect 8628 13268 8634 13280
rect 9033 13277 9045 13280
rect 9079 13277 9091 13311
rect 9033 13271 9091 13277
rect 9122 13268 9128 13320
rect 9180 13308 9186 13320
rect 13081 13311 13139 13317
rect 9180 13280 9225 13308
rect 9180 13268 9186 13280
rect 13081 13277 13093 13311
rect 13127 13277 13139 13311
rect 14550 13308 14556 13320
rect 14511 13280 14556 13308
rect 13081 13271 13139 13277
rect 12710 13240 12716 13252
rect 5920 13212 12716 13240
rect 1118 13132 1124 13184
rect 1176 13172 1182 13184
rect 5920 13172 5948 13212
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 1176 13144 5948 13172
rect 1176 13132 1182 13144
rect 5994 13132 6000 13184
rect 6052 13172 6058 13184
rect 6052 13144 6097 13172
rect 6052 13132 6058 13144
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 9306 13172 9312 13184
rect 6880 13144 9312 13172
rect 6880 13132 6886 13144
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 13096 13172 13124 13271
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 14458 13172 14464 13184
rect 13096 13144 14464 13172
rect 14458 13132 14464 13144
rect 14516 13132 14522 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 3694 12928 3700 12980
rect 3752 12968 3758 12980
rect 5534 12968 5540 12980
rect 3752 12940 5540 12968
rect 3752 12928 3758 12940
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 5718 12968 5724 12980
rect 5679 12940 5724 12968
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 6362 12968 6368 12980
rect 5951 12940 6368 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 6362 12928 6368 12940
rect 6420 12928 6426 12980
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 13722 12968 13728 12980
rect 13412 12940 13728 12968
rect 13412 12928 13418 12940
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 15841 12971 15899 12977
rect 15841 12968 15853 12971
rect 14292 12940 15853 12968
rect 5736 12832 5764 12928
rect 12805 12903 12863 12909
rect 12805 12869 12817 12903
rect 12851 12900 12863 12903
rect 13906 12900 13912 12912
rect 12851 12872 13912 12900
rect 12851 12869 12863 12872
rect 12805 12863 12863 12869
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 6457 12835 6515 12841
rect 6457 12832 6469 12835
rect 5736 12804 6469 12832
rect 6457 12801 6469 12804
rect 6503 12801 6515 12835
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6457 12795 6515 12801
rect 7116 12804 7389 12832
rect 3786 12724 3792 12776
rect 3844 12764 3850 12776
rect 4338 12764 4344 12776
rect 3844 12736 4344 12764
rect 3844 12724 3850 12736
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 4608 12699 4666 12705
rect 4608 12665 4620 12699
rect 4654 12696 4666 12699
rect 6178 12696 6184 12708
rect 4654 12668 6184 12696
rect 4654 12665 4666 12668
rect 4608 12659 4666 12665
rect 6178 12656 6184 12668
rect 6236 12696 6242 12708
rect 6730 12696 6736 12708
rect 6236 12668 6736 12696
rect 6236 12656 6242 12668
rect 6730 12656 6736 12668
rect 6788 12696 6794 12708
rect 7116 12696 7144 12804
rect 7377 12801 7389 12804
rect 7423 12832 7435 12835
rect 13449 12835 13507 12841
rect 7423 12804 7972 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 7558 12764 7564 12776
rect 7340 12736 7564 12764
rect 7340 12724 7346 12736
rect 7558 12724 7564 12736
rect 7616 12764 7622 12776
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7616 12736 7849 12764
rect 7616 12724 7622 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 6788 12668 7144 12696
rect 7193 12699 7251 12705
rect 6788 12656 6794 12668
rect 7193 12665 7205 12699
rect 7239 12696 7251 12699
rect 7374 12696 7380 12708
rect 7239 12668 7380 12696
rect 7239 12665 7251 12668
rect 7193 12659 7251 12665
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 5994 12588 6000 12640
rect 6052 12628 6058 12640
rect 6273 12631 6331 12637
rect 6273 12628 6285 12631
rect 6052 12600 6285 12628
rect 6052 12588 6058 12600
rect 6273 12597 6285 12600
rect 6319 12597 6331 12631
rect 6273 12591 6331 12597
rect 6365 12631 6423 12637
rect 6365 12597 6377 12631
rect 6411 12628 6423 12631
rect 6825 12631 6883 12637
rect 6825 12628 6837 12631
rect 6411 12600 6837 12628
rect 6411 12597 6423 12600
rect 6365 12591 6423 12597
rect 6825 12597 6837 12600
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 7285 12631 7343 12637
rect 7285 12597 7297 12631
rect 7331 12628 7343 12631
rect 7466 12628 7472 12640
rect 7331 12600 7472 12628
rect 7331 12597 7343 12600
rect 7285 12591 7343 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 7650 12628 7656 12640
rect 7611 12600 7656 12628
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 7944 12628 7972 12804
rect 13449 12801 13461 12835
rect 13495 12832 13507 12835
rect 13814 12832 13820 12844
rect 13495 12804 13820 12832
rect 13495 12801 13507 12804
rect 13449 12795 13507 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14182 12792 14188 12844
rect 14240 12832 14246 12844
rect 14292 12841 14320 12940
rect 15841 12937 15853 12940
rect 15887 12937 15899 12971
rect 16942 12968 16948 12980
rect 16903 12940 16948 12968
rect 15841 12931 15899 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 14277 12835 14335 12841
rect 14277 12832 14289 12835
rect 14240 12804 14289 12832
rect 14240 12792 14246 12804
rect 14277 12801 14289 12804
rect 14323 12801 14335 12835
rect 14458 12832 14464 12844
rect 14419 12804 14464 12832
rect 14277 12795 14335 12801
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 16758 12832 16764 12844
rect 16719 12804 16764 12832
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 8104 12767 8162 12773
rect 8104 12733 8116 12767
rect 8150 12764 8162 12767
rect 8386 12764 8392 12776
rect 8150 12736 8392 12764
rect 8150 12733 8162 12736
rect 8104 12727 8162 12733
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 14366 12764 14372 12776
rect 13311 12736 14372 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 14366 12724 14372 12736
rect 14424 12724 14430 12776
rect 14476 12764 14504 12792
rect 15010 12764 15016 12776
rect 14476 12736 15016 12764
rect 15010 12724 15016 12736
rect 15068 12724 15074 12776
rect 16485 12767 16543 12773
rect 16485 12764 16497 12767
rect 15948 12736 16497 12764
rect 13173 12699 13231 12705
rect 13173 12665 13185 12699
rect 13219 12696 13231 12699
rect 14728 12699 14786 12705
rect 13219 12668 13676 12696
rect 13219 12665 13231 12668
rect 13173 12659 13231 12665
rect 13648 12637 13676 12668
rect 14728 12665 14740 12699
rect 14774 12696 14786 12699
rect 14918 12696 14924 12708
rect 14774 12668 14924 12696
rect 14774 12665 14786 12668
rect 14728 12659 14786 12665
rect 14918 12656 14924 12668
rect 14976 12656 14982 12708
rect 15948 12640 15976 12736
rect 16485 12733 16497 12736
rect 16531 12733 16543 12767
rect 16960 12764 16988 12928
rect 17678 12832 17684 12844
rect 17639 12804 17684 12832
rect 17678 12792 17684 12804
rect 17736 12792 17742 12844
rect 17589 12767 17647 12773
rect 17589 12764 17601 12767
rect 16960 12736 17601 12764
rect 16485 12727 16543 12733
rect 17589 12733 17601 12736
rect 17635 12733 17647 12767
rect 17589 12727 17647 12733
rect 16298 12656 16304 12708
rect 16356 12696 16362 12708
rect 16577 12699 16635 12705
rect 16577 12696 16589 12699
rect 16356 12668 16589 12696
rect 16356 12656 16362 12668
rect 16577 12665 16589 12668
rect 16623 12665 16635 12699
rect 16577 12659 16635 12665
rect 9217 12631 9275 12637
rect 9217 12628 9229 12631
rect 7944 12600 9229 12628
rect 9217 12597 9229 12600
rect 9263 12597 9275 12631
rect 9217 12591 9275 12597
rect 13633 12631 13691 12637
rect 13633 12597 13645 12631
rect 13679 12597 13691 12631
rect 13998 12628 14004 12640
rect 13959 12600 14004 12628
rect 13633 12591 13691 12597
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 14090 12588 14096 12640
rect 14148 12628 14154 12640
rect 15930 12628 15936 12640
rect 14148 12600 14193 12628
rect 15891 12600 15936 12628
rect 14148 12588 14154 12600
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16114 12628 16120 12640
rect 16075 12600 16120 12628
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 17126 12628 17132 12640
rect 17087 12600 17132 12628
rect 17126 12588 17132 12600
rect 17184 12588 17190 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 17497 12631 17555 12637
rect 17497 12628 17509 12631
rect 17460 12600 17509 12628
rect 17460 12588 17466 12600
rect 17497 12597 17509 12600
rect 17543 12628 17555 12631
rect 18049 12631 18107 12637
rect 18049 12628 18061 12631
rect 17543 12600 18061 12628
rect 17543 12597 17555 12600
rect 17497 12591 17555 12597
rect 18049 12597 18061 12600
rect 18095 12597 18107 12631
rect 18049 12591 18107 12597
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 5721 12427 5779 12433
rect 5721 12393 5733 12427
rect 5767 12424 5779 12427
rect 5994 12424 6000 12436
rect 5767 12396 6000 12424
rect 5767 12393 5779 12396
rect 5721 12387 5779 12393
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 6181 12427 6239 12433
rect 6181 12393 6193 12427
rect 6227 12424 6239 12427
rect 6549 12427 6607 12433
rect 6549 12424 6561 12427
rect 6227 12396 6561 12424
rect 6227 12393 6239 12396
rect 6181 12387 6239 12393
rect 6549 12393 6561 12396
rect 6595 12393 6607 12427
rect 7374 12424 7380 12436
rect 7335 12396 7380 12424
rect 6549 12387 6607 12393
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 9674 12424 9680 12436
rect 7484 12396 9680 12424
rect 3970 12316 3976 12368
rect 4028 12356 4034 12368
rect 4332 12359 4390 12365
rect 4028 12328 4292 12356
rect 4028 12316 4034 12328
rect 4264 12288 4292 12328
rect 4332 12325 4344 12359
rect 4378 12356 4390 12359
rect 5902 12356 5908 12368
rect 4378 12328 5908 12356
rect 4378 12325 4390 12328
rect 4332 12319 4390 12325
rect 5902 12316 5908 12328
rect 5960 12316 5966 12368
rect 6012 12328 6408 12356
rect 6012 12300 6040 12328
rect 5994 12288 6000 12300
rect 4264 12260 6000 12288
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12257 6147 12291
rect 6380 12288 6408 12328
rect 6454 12316 6460 12368
rect 6512 12356 6518 12368
rect 7009 12359 7067 12365
rect 7009 12356 7021 12359
rect 6512 12328 7021 12356
rect 6512 12316 6518 12328
rect 7009 12325 7021 12328
rect 7055 12356 7067 12359
rect 7484 12356 7512 12396
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10137 12427 10195 12433
rect 10137 12393 10149 12427
rect 10183 12424 10195 12427
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10183 12396 10701 12424
rect 10183 12393 10195 12396
rect 10137 12387 10195 12393
rect 10689 12393 10701 12396
rect 10735 12424 10747 12427
rect 13170 12424 13176 12436
rect 10735 12396 13176 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 14148 12396 14289 12424
rect 14148 12384 14154 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 14277 12387 14335 12393
rect 14366 12384 14372 12436
rect 14424 12424 14430 12436
rect 15473 12427 15531 12433
rect 15473 12424 15485 12427
rect 14424 12396 15485 12424
rect 14424 12384 14430 12396
rect 15473 12393 15485 12396
rect 15519 12393 15531 12427
rect 15473 12387 15531 12393
rect 15841 12427 15899 12433
rect 15841 12393 15853 12427
rect 15887 12424 15899 12427
rect 16114 12424 16120 12436
rect 15887 12396 16120 12424
rect 15887 12393 15899 12396
rect 15841 12387 15899 12393
rect 16114 12384 16120 12396
rect 16172 12384 16178 12436
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16758 12424 16764 12436
rect 16264 12396 16764 12424
rect 16264 12384 16270 12396
rect 16758 12384 16764 12396
rect 16816 12424 16822 12436
rect 17681 12427 17739 12433
rect 17681 12424 17693 12427
rect 16816 12396 17693 12424
rect 16816 12384 16822 12396
rect 17681 12393 17693 12396
rect 17727 12393 17739 12427
rect 17681 12387 17739 12393
rect 8202 12356 8208 12368
rect 7055 12328 7512 12356
rect 8163 12328 8208 12356
rect 7055 12325 7067 12328
rect 7009 12319 7067 12325
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 8573 12359 8631 12365
rect 8573 12325 8585 12359
rect 8619 12356 8631 12359
rect 8619 12328 9260 12356
rect 8619 12325 8631 12328
rect 8573 12319 8631 12325
rect 6730 12288 6736 12300
rect 6380 12260 6736 12288
rect 6089 12251 6147 12257
rect 1486 12180 1492 12232
rect 1544 12220 1550 12232
rect 2133 12223 2191 12229
rect 2133 12220 2145 12223
rect 1544 12192 2145 12220
rect 1544 12180 1550 12192
rect 2133 12189 2145 12192
rect 2179 12220 2191 12223
rect 2774 12220 2780 12232
rect 2179 12192 2780 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2774 12180 2780 12192
rect 2832 12180 2838 12232
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3844 12192 4077 12220
rect 3844 12180 3850 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5629 12223 5687 12229
rect 5629 12220 5641 12223
rect 5592 12192 5641 12220
rect 5592 12180 5598 12192
rect 5629 12189 5641 12192
rect 5675 12220 5687 12223
rect 5902 12220 5908 12232
rect 5675 12192 5908 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 5902 12180 5908 12192
rect 5960 12220 5966 12232
rect 6104 12220 6132 12251
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 6914 12288 6920 12300
rect 6875 12260 6920 12288
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 7745 12291 7803 12297
rect 7745 12288 7757 12291
rect 7024 12260 7757 12288
rect 5960 12192 6132 12220
rect 5960 12180 5966 12192
rect 6178 12180 6184 12232
rect 6236 12220 6242 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 6236 12192 6285 12220
rect 6236 12180 6242 12192
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 7024 12152 7052 12260
rect 7745 12257 7757 12260
rect 7791 12288 7803 12291
rect 8588 12288 8616 12319
rect 7791 12260 8616 12288
rect 7791 12257 7803 12260
rect 7745 12251 7803 12257
rect 9030 12248 9036 12300
rect 9088 12288 9094 12300
rect 9125 12291 9183 12297
rect 9125 12288 9137 12291
rect 9088 12260 9137 12288
rect 9088 12248 9094 12260
rect 9125 12257 9137 12260
rect 9171 12257 9183 12291
rect 9232 12288 9260 12328
rect 9306 12316 9312 12368
rect 9364 12356 9370 12368
rect 12342 12356 12348 12368
rect 9364 12328 12348 12356
rect 9364 12316 9370 12328
rect 12342 12316 12348 12328
rect 12400 12316 12406 12368
rect 12980 12359 13038 12365
rect 12980 12325 12992 12359
rect 13026 12356 13038 12359
rect 14182 12356 14188 12368
rect 13026 12328 14188 12356
rect 13026 12325 13038 12328
rect 12980 12319 13038 12325
rect 14182 12316 14188 12328
rect 14240 12356 14246 12368
rect 14240 12328 16436 12356
rect 14240 12316 14246 12328
rect 10594 12288 10600 12300
rect 9232 12260 10600 12288
rect 9125 12251 9183 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 10704 12260 13768 12288
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12189 7251 12223
rect 7193 12183 7251 12189
rect 5276 12124 7052 12152
rect 7208 12152 7236 12183
rect 7374 12180 7380 12232
rect 7432 12220 7438 12232
rect 7650 12220 7656 12232
rect 7432 12192 7656 12220
rect 7432 12180 7438 12192
rect 7650 12180 7656 12192
rect 7708 12220 7714 12232
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 7708 12192 7849 12220
rect 7708 12180 7714 12192
rect 7837 12189 7849 12192
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12220 8079 12223
rect 8386 12220 8392 12232
rect 8067 12192 8392 12220
rect 8067 12189 8079 12192
rect 8021 12183 8079 12189
rect 8036 12152 8064 12183
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 9214 12220 9220 12232
rect 9175 12192 9220 12220
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 9364 12192 9409 12220
rect 9364 12180 9370 12192
rect 9582 12180 9588 12232
rect 9640 12180 9646 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10704 12220 10732 12260
rect 9732 12192 10732 12220
rect 10873 12223 10931 12229
rect 9732 12180 9738 12192
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 10962 12220 10968 12232
rect 10919 12192 10968 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 12710 12220 12716 12232
rect 12671 12192 12716 12220
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 13740 12220 13768 12260
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 14645 12291 14703 12297
rect 14645 12288 14657 12291
rect 14424 12260 14657 12288
rect 14424 12248 14430 12260
rect 14645 12257 14657 12260
rect 14691 12257 14703 12291
rect 14645 12251 14703 12257
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 15068 12260 16313 12288
rect 15068 12248 15074 12260
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 16301 12251 16359 12257
rect 14737 12223 14795 12229
rect 13740 12192 14596 12220
rect 7208 12124 8064 12152
rect 9600 12152 9628 12180
rect 9600 12124 12756 12152
rect 2130 12044 2136 12096
rect 2188 12084 2194 12096
rect 4246 12084 4252 12096
rect 2188 12056 4252 12084
rect 2188 12044 2194 12056
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 5276 12084 5304 12124
rect 5442 12084 5448 12096
rect 4764 12056 5304 12084
rect 5403 12056 5448 12084
rect 4764 12044 4770 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 8757 12087 8815 12093
rect 8757 12053 8769 12087
rect 8803 12084 8815 12087
rect 9030 12084 9036 12096
rect 8803 12056 9036 12084
rect 8803 12053 8815 12056
rect 8757 12047 8815 12053
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 10226 12084 10232 12096
rect 10187 12056 10232 12084
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 11149 12087 11207 12093
rect 11149 12084 11161 12087
rect 10652 12056 11161 12084
rect 10652 12044 10658 12056
rect 11149 12053 11161 12056
rect 11195 12084 11207 12087
rect 12250 12084 12256 12096
rect 11195 12056 12256 12084
rect 11195 12053 11207 12056
rect 11149 12047 11207 12053
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12728 12084 12756 12124
rect 13814 12112 13820 12164
rect 13872 12152 13878 12164
rect 14093 12155 14151 12161
rect 14093 12152 14105 12155
rect 13872 12124 14105 12152
rect 13872 12112 13878 12124
rect 14093 12121 14105 12124
rect 14139 12121 14151 12155
rect 14093 12115 14151 12121
rect 14458 12084 14464 12096
rect 12728 12056 14464 12084
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 14568 12084 14596 12192
rect 14737 12189 14749 12223
rect 14783 12189 14795 12223
rect 14918 12220 14924 12232
rect 14879 12192 14924 12220
rect 14737 12183 14795 12189
rect 14752 12152 14780 12183
rect 14918 12180 14924 12192
rect 14976 12180 14982 12232
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15252 12192 15945 12220
rect 15252 12180 15258 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16117 12223 16175 12229
rect 16117 12189 16129 12223
rect 16163 12220 16175 12223
rect 16408 12220 16436 12328
rect 16666 12316 16672 12368
rect 16724 12316 16730 12368
rect 16568 12291 16626 12297
rect 16568 12257 16580 12291
rect 16614 12288 16626 12291
rect 16684 12288 16712 12316
rect 17678 12288 17684 12300
rect 16614 12260 17684 12288
rect 16614 12257 16626 12260
rect 16568 12251 16626 12257
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 18138 12288 18144 12300
rect 18099 12260 18144 12288
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 16163 12192 16436 12220
rect 16163 12189 16175 12192
rect 16117 12183 16175 12189
rect 17770 12180 17776 12232
rect 17828 12220 17834 12232
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 17828 12192 18245 12220
rect 17828 12180 17834 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 15378 12152 15384 12164
rect 14752 12124 15384 12152
rect 15378 12112 15384 12124
rect 15436 12112 15442 12164
rect 17678 12112 17684 12164
rect 17736 12152 17742 12164
rect 18340 12152 18368 12183
rect 17736 12124 18368 12152
rect 17736 12112 17742 12124
rect 14826 12084 14832 12096
rect 14568 12056 14832 12084
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 17773 12087 17831 12093
rect 17773 12084 17785 12087
rect 16172 12056 17785 12084
rect 16172 12044 16178 12056
rect 17773 12053 17785 12056
rect 17819 12053 17831 12087
rect 17773 12047 17831 12053
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 3602 11880 3608 11892
rect 3563 11852 3608 11880
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 9214 11880 9220 11892
rect 6788 11852 9220 11880
rect 6788 11840 6794 11852
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9306 11840 9312 11892
rect 9364 11880 9370 11892
rect 11241 11883 11299 11889
rect 11241 11880 11253 11883
rect 9364 11852 11253 11880
rect 9364 11840 9370 11852
rect 11241 11849 11253 11852
rect 11287 11849 11299 11883
rect 11241 11843 11299 11849
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 12584 11852 13952 11880
rect 12584 11840 12590 11852
rect 5350 11772 5356 11824
rect 5408 11812 5414 11824
rect 7101 11815 7159 11821
rect 7101 11812 7113 11815
rect 5408 11784 7113 11812
rect 5408 11772 5414 11784
rect 7101 11781 7113 11784
rect 7147 11812 7159 11815
rect 7558 11812 7564 11824
rect 7147 11784 7564 11812
rect 7147 11781 7159 11784
rect 7101 11775 7159 11781
rect 7558 11772 7564 11784
rect 7616 11812 7622 11824
rect 10318 11812 10324 11824
rect 7616 11784 7972 11812
rect 10231 11784 10324 11812
rect 7616 11772 7622 11784
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11713 2099 11747
rect 2041 11707 2099 11713
rect 2056 11676 2084 11707
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 2869 11747 2927 11753
rect 2869 11744 2881 11747
rect 2464 11716 2881 11744
rect 2464 11704 2470 11716
rect 2869 11713 2881 11716
rect 2915 11744 2927 11747
rect 3697 11747 3755 11753
rect 3697 11744 3709 11747
rect 2915 11716 3709 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 3697 11713 3709 11716
rect 3743 11713 3755 11747
rect 3697 11707 3755 11713
rect 7009 11747 7067 11753
rect 7009 11713 7021 11747
rect 7055 11744 7067 11747
rect 7837 11747 7895 11753
rect 7837 11744 7849 11747
rect 7055 11716 7849 11744
rect 7055 11713 7067 11716
rect 7009 11707 7067 11713
rect 2682 11676 2688 11688
rect 2056 11648 2688 11676
rect 2682 11636 2688 11648
rect 2740 11636 2746 11688
rect 3789 11679 3847 11685
rect 3789 11645 3801 11679
rect 3835 11676 3847 11679
rect 3878 11676 3884 11688
rect 3835 11648 3884 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4056 11679 4114 11685
rect 4056 11645 4068 11679
rect 4102 11676 4114 11679
rect 4614 11676 4620 11688
rect 4102 11648 4620 11676
rect 4102 11645 4114 11648
rect 4056 11639 4114 11645
rect 4614 11636 4620 11648
rect 4672 11676 4678 11688
rect 5442 11676 5448 11688
rect 4672 11648 5448 11676
rect 4672 11636 4678 11648
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 5592 11648 7297 11676
rect 5592 11636 5598 11648
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 1578 11568 1584 11620
rect 1636 11608 1642 11620
rect 2593 11611 2651 11617
rect 1636 11580 2544 11608
rect 1636 11568 1642 11580
rect 1394 11540 1400 11552
rect 1355 11512 1400 11540
rect 1394 11500 1400 11512
rect 1452 11500 1458 11552
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 1857 11543 1915 11549
rect 1857 11509 1869 11543
rect 1903 11540 1915 11543
rect 2225 11543 2283 11549
rect 2225 11540 2237 11543
rect 1903 11512 2237 11540
rect 1903 11509 1915 11512
rect 1857 11503 1915 11509
rect 2225 11509 2237 11512
rect 2271 11509 2283 11543
rect 2516 11540 2544 11580
rect 2593 11577 2605 11611
rect 2639 11608 2651 11611
rect 2774 11608 2780 11620
rect 2639 11580 2780 11608
rect 2639 11577 2651 11580
rect 2593 11571 2651 11577
rect 2774 11568 2780 11580
rect 2832 11568 2838 11620
rect 3329 11611 3387 11617
rect 3329 11608 3341 11611
rect 2976 11580 3341 11608
rect 2685 11543 2743 11549
rect 2685 11540 2697 11543
rect 2516 11512 2697 11540
rect 2225 11503 2283 11509
rect 2685 11509 2697 11512
rect 2731 11540 2743 11543
rect 2976 11540 3004 11580
rect 3329 11577 3341 11580
rect 3375 11608 3387 11611
rect 5810 11608 5816 11620
rect 3375 11580 5816 11608
rect 3375 11577 3387 11580
rect 3329 11571 3387 11577
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 6641 11611 6699 11617
rect 6641 11577 6653 11611
rect 6687 11608 6699 11611
rect 6914 11608 6920 11620
rect 6687 11580 6920 11608
rect 6687 11577 6699 11580
rect 6641 11571 6699 11577
rect 6914 11568 6920 11580
rect 6972 11608 6978 11620
rect 7558 11608 7564 11620
rect 6972 11580 7564 11608
rect 6972 11568 6978 11580
rect 7558 11568 7564 11580
rect 7616 11568 7622 11620
rect 2731 11512 3004 11540
rect 2731 11509 2743 11512
rect 2685 11503 2743 11509
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 3697 11543 3755 11549
rect 3108 11512 3153 11540
rect 3108 11500 3114 11512
rect 3697 11509 3709 11543
rect 3743 11540 3755 11543
rect 3786 11540 3792 11552
rect 3743 11512 3792 11540
rect 3743 11509 3755 11512
rect 3697 11503 3755 11509
rect 3786 11500 3792 11512
rect 3844 11540 3850 11552
rect 5169 11543 5227 11549
rect 5169 11540 5181 11543
rect 3844 11512 5181 11540
rect 3844 11500 3850 11512
rect 5169 11509 5181 11512
rect 5215 11509 5227 11543
rect 5169 11503 5227 11509
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 5684 11512 6377 11540
rect 5684 11500 5690 11512
rect 6365 11509 6377 11512
rect 6411 11540 6423 11543
rect 6454 11540 6460 11552
rect 6411 11512 6460 11540
rect 6411 11509 6423 11512
rect 6365 11503 6423 11509
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 7377 11543 7435 11549
rect 7377 11509 7389 11543
rect 7423 11540 7435 11543
rect 7466 11540 7472 11552
rect 7423 11512 7472 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 7668 11540 7696 11716
rect 7837 11713 7849 11716
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 7944 11688 7972 11784
rect 10318 11772 10324 11784
rect 10376 11812 10382 11824
rect 10686 11812 10692 11824
rect 10376 11784 10692 11812
rect 10376 11772 10382 11784
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 13924 11812 13952 11852
rect 13998 11840 14004 11892
rect 14056 11880 14062 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 14056 11852 14289 11880
rect 14056 11840 14062 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 15194 11880 15200 11892
rect 15155 11852 15200 11880
rect 14277 11843 14335 11849
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 16025 11883 16083 11889
rect 16025 11849 16037 11883
rect 16071 11880 16083 11883
rect 16298 11880 16304 11892
rect 16071 11852 16304 11880
rect 16071 11849 16083 11852
rect 16025 11843 16083 11849
rect 16298 11840 16304 11852
rect 16356 11840 16362 11892
rect 17126 11880 17132 11892
rect 16399 11852 17132 11880
rect 14093 11815 14151 11821
rect 14093 11812 14105 11815
rect 10796 11784 12204 11812
rect 13924 11784 14105 11812
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11744 8079 11747
rect 8386 11744 8392 11756
rect 8067 11716 8392 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 10594 11744 10600 11756
rect 10152 11716 10600 11744
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 7984 11648 8953 11676
rect 7984 11636 7990 11648
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 10152 11676 10180 11716
rect 10594 11704 10600 11716
rect 10652 11744 10658 11756
rect 10796 11744 10824 11784
rect 10962 11744 10968 11756
rect 10652 11716 10824 11744
rect 10923 11716 10968 11744
rect 10652 11704 10658 11716
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11793 11747 11851 11753
rect 11793 11744 11805 11747
rect 11112 11716 11805 11744
rect 11112 11704 11118 11716
rect 11793 11713 11805 11716
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 8941 11639 8999 11645
rect 9140 11648 10180 11676
rect 7745 11611 7803 11617
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 8297 11611 8355 11617
rect 8297 11608 8309 11611
rect 7791 11580 8309 11608
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 8297 11577 8309 11580
rect 8343 11608 8355 11611
rect 9140 11608 9168 11648
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 12176 11685 12204 11784
rect 14093 11781 14105 11784
rect 14139 11812 14151 11815
rect 14366 11812 14372 11824
rect 14139 11784 14372 11812
rect 14139 11781 14151 11784
rect 14093 11775 14151 11781
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 16399 11812 16427 11852
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17770 11880 17776 11892
rect 17731 11852 17776 11880
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 18138 11840 18144 11892
rect 18196 11880 18202 11892
rect 18417 11883 18475 11889
rect 18417 11880 18429 11883
rect 18196 11852 18429 11880
rect 18196 11840 18202 11852
rect 18417 11849 18429 11852
rect 18463 11849 18475 11883
rect 18417 11843 18475 11849
rect 15580 11784 15884 11812
rect 12618 11744 12624 11756
rect 12579 11716 12624 11744
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 13170 11704 13176 11756
rect 13228 11744 13234 11756
rect 13265 11747 13323 11753
rect 13265 11744 13277 11747
rect 13228 11716 13277 11744
rect 13228 11704 13234 11716
rect 13265 11713 13277 11716
rect 13311 11713 13323 11747
rect 13265 11707 13323 11713
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11744 14059 11747
rect 14734 11744 14740 11756
rect 14047 11716 14740 11744
rect 14047 11713 14059 11716
rect 14001 11707 14059 11713
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 14918 11744 14924 11756
rect 14831 11716 14924 11744
rect 14918 11704 14924 11716
rect 14976 11744 14982 11756
rect 15580 11744 15608 11784
rect 15856 11753 15884 11784
rect 16316 11784 16427 11812
rect 14976 11716 15608 11744
rect 15841 11747 15899 11753
rect 14976 11704 14982 11716
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16206 11744 16212 11756
rect 15887 11716 16212 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 11609 11679 11667 11685
rect 11609 11676 11621 11679
rect 10284 11648 11621 11676
rect 10284 11636 10290 11648
rect 11609 11645 11621 11648
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 12161 11679 12219 11685
rect 12161 11645 12173 11679
rect 12207 11676 12219 11679
rect 13538 11676 13544 11688
rect 12207 11648 13544 11676
rect 12207 11645 12219 11648
rect 12161 11639 12219 11645
rect 13538 11636 13544 11648
rect 13596 11636 13602 11688
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 14608 11648 14657 11676
rect 14608 11636 14614 11648
rect 14645 11645 14657 11648
rect 14691 11645 14703 11679
rect 14645 11639 14703 11645
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11676 15715 11679
rect 16114 11676 16120 11688
rect 15703 11648 16120 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 9214 11617 9220 11620
rect 8343 11580 9168 11608
rect 8343 11577 8355 11580
rect 8297 11571 8355 11577
rect 9208 11571 9220 11617
rect 9272 11608 9278 11620
rect 11701 11611 11759 11617
rect 11701 11608 11713 11611
rect 9272 11580 9308 11608
rect 10428 11580 11713 11608
rect 9214 11568 9220 11571
rect 9272 11568 9278 11580
rect 10134 11540 10140 11552
rect 7668 11512 10140 11540
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10428 11549 10456 11580
rect 11701 11577 11713 11580
rect 11747 11577 11759 11611
rect 11701 11571 11759 11577
rect 13081 11611 13139 11617
rect 13081 11577 13093 11611
rect 13127 11608 13139 11611
rect 13998 11608 14004 11620
rect 13127 11580 14004 11608
rect 13127 11577 13139 11580
rect 13081 11571 13139 11577
rect 13998 11568 14004 11580
rect 14056 11568 14062 11620
rect 10413 11543 10471 11549
rect 10413 11509 10425 11543
rect 10459 11509 10471 11543
rect 10413 11503 10471 11509
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 10652 11512 10793 11540
rect 10652 11500 10658 11512
rect 10781 11509 10793 11512
rect 10827 11509 10839 11543
rect 10781 11503 10839 11509
rect 10873 11543 10931 11549
rect 10873 11509 10885 11543
rect 10919 11540 10931 11543
rect 11054 11540 11060 11552
rect 10919 11512 11060 11540
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 12713 11543 12771 11549
rect 12713 11540 12725 11543
rect 11296 11512 12725 11540
rect 11296 11500 11302 11512
rect 12713 11509 12725 11512
rect 12759 11509 12771 11543
rect 12713 11503 12771 11509
rect 13173 11543 13231 11549
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 13262 11540 13268 11552
rect 13219 11512 13268 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 15565 11543 15623 11549
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 16316 11540 16344 11784
rect 16574 11772 16580 11824
rect 16632 11812 16638 11824
rect 16853 11815 16911 11821
rect 16853 11812 16865 11815
rect 16632 11784 16865 11812
rect 16632 11772 16638 11784
rect 16853 11781 16865 11784
rect 16899 11781 16911 11815
rect 16853 11775 16911 11781
rect 16666 11744 16672 11756
rect 16627 11716 16672 11744
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 17494 11744 17500 11756
rect 17455 11716 17500 11744
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 16393 11611 16451 11617
rect 16393 11577 16405 11611
rect 16439 11608 16451 11611
rect 16942 11608 16948 11620
rect 16439 11580 16948 11608
rect 16439 11577 16451 11580
rect 16393 11571 16451 11577
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 15611 11512 16344 11540
rect 16485 11543 16543 11549
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 16485 11509 16497 11543
rect 16531 11540 16543 11543
rect 16758 11540 16764 11552
rect 16531 11512 16764 11540
rect 16531 11509 16543 11512
rect 16485 11503 16543 11509
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 17218 11540 17224 11552
rect 17179 11512 17224 11540
rect 17218 11500 17224 11512
rect 17276 11500 17282 11552
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 17368 11512 17413 11540
rect 17368 11500 17374 11512
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 2682 11296 2688 11348
rect 2740 11336 2746 11348
rect 3513 11339 3571 11345
rect 3513 11336 3525 11339
rect 2740 11308 3525 11336
rect 2740 11296 2746 11308
rect 3513 11305 3525 11308
rect 3559 11305 3571 11339
rect 3513 11299 3571 11305
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 9125 11339 9183 11345
rect 9125 11305 9137 11339
rect 9171 11336 9183 11339
rect 9214 11336 9220 11348
rect 9171 11308 9220 11336
rect 9171 11305 9183 11308
rect 9125 11299 9183 11305
rect 2406 11277 2412 11280
rect 2400 11268 2412 11277
rect 2367 11240 2412 11268
rect 2400 11231 2412 11240
rect 2406 11228 2412 11231
rect 2464 11228 2470 11280
rect 3602 11228 3608 11280
rect 3660 11228 3666 11280
rect 1946 11160 1952 11212
rect 2004 11200 2010 11212
rect 2041 11203 2099 11209
rect 2041 11200 2053 11203
rect 2004 11172 2053 11200
rect 2004 11160 2010 11172
rect 2041 11169 2053 11172
rect 2087 11200 2099 11203
rect 2958 11200 2964 11212
rect 2087 11172 2964 11200
rect 2087 11169 2099 11172
rect 2041 11163 2099 11169
rect 2958 11160 2964 11172
rect 3016 11200 3022 11212
rect 3620 11200 3648 11228
rect 3016 11172 3648 11200
rect 3789 11203 3847 11209
rect 3016 11160 3022 11172
rect 3789 11169 3801 11203
rect 3835 11200 3847 11203
rect 5534 11200 5540 11212
rect 3835 11172 5540 11200
rect 3835 11169 3847 11172
rect 3789 11163 3847 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5718 11209 5724 11212
rect 5712 11200 5724 11209
rect 5631 11172 5724 11200
rect 5712 11163 5724 11172
rect 5776 11200 5782 11212
rect 6178 11200 6184 11212
rect 5776 11172 6184 11200
rect 5718 11160 5724 11163
rect 5776 11160 5782 11172
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6840 11200 6868 11299
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 10045 11339 10103 11345
rect 10045 11336 10057 11339
rect 9364 11308 10057 11336
rect 9364 11296 9370 11308
rect 10045 11305 10057 11308
rect 10091 11336 10103 11339
rect 10597 11339 10655 11345
rect 10597 11336 10609 11339
rect 10091 11308 10609 11336
rect 10091 11305 10103 11308
rect 10045 11299 10103 11305
rect 10597 11305 10609 11308
rect 10643 11305 10655 11339
rect 11054 11336 11060 11348
rect 11015 11308 11060 11336
rect 10597 11299 10655 11305
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 11146 11296 11152 11348
rect 11204 11336 11210 11348
rect 13262 11336 13268 11348
rect 11204 11308 11249 11336
rect 13223 11308 13268 11336
rect 11204 11296 11210 11308
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13633 11339 13691 11345
rect 13633 11305 13645 11339
rect 13679 11336 13691 11339
rect 13814 11336 13820 11348
rect 13679 11308 13820 11336
rect 13679 11305 13691 11308
rect 13633 11299 13691 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 14056 11308 14105 11336
rect 14056 11296 14062 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 14553 11339 14611 11345
rect 14553 11305 14565 11339
rect 14599 11336 14611 11339
rect 14642 11336 14648 11348
rect 14599 11308 14648 11336
rect 14599 11305 14611 11308
rect 14553 11299 14611 11305
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 14921 11339 14979 11345
rect 14921 11305 14933 11339
rect 14967 11336 14979 11339
rect 15010 11336 15016 11348
rect 14967 11308 15016 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16853 11339 16911 11345
rect 16853 11336 16865 11339
rect 16724 11308 16865 11336
rect 16724 11296 16730 11308
rect 16853 11305 16865 11308
rect 16899 11305 16911 11339
rect 16853 11299 16911 11305
rect 17218 11296 17224 11348
rect 17276 11336 17282 11348
rect 17497 11339 17555 11345
rect 17497 11336 17509 11339
rect 17276 11308 17509 11336
rect 17276 11296 17282 11308
rect 17497 11305 17509 11308
rect 17543 11305 17555 11339
rect 17497 11299 17555 11305
rect 17957 11339 18015 11345
rect 17957 11305 17969 11339
rect 18003 11336 18015 11339
rect 18414 11336 18420 11348
rect 18003 11308 18420 11336
rect 18003 11305 18015 11308
rect 17957 11299 18015 11305
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 7990 11271 8048 11277
rect 7990 11268 8002 11271
rect 7116 11240 8002 11268
rect 7116 11200 7144 11240
rect 7990 11237 8002 11240
rect 8036 11268 8048 11271
rect 8202 11268 8208 11280
rect 8036 11240 8208 11268
rect 8036 11237 8048 11240
rect 7990 11231 8048 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 9232 11268 9260 11296
rect 10686 11268 10692 11280
rect 9232 11240 10692 11268
rect 10686 11228 10692 11240
rect 10744 11268 10750 11280
rect 10962 11268 10968 11280
rect 10744 11240 10968 11268
rect 10744 11228 10750 11240
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 12802 11268 12808 11280
rect 11256 11240 12808 11268
rect 7282 11200 7288 11212
rect 6840 11172 7144 11200
rect 7243 11172 7288 11200
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11200 7803 11203
rect 7834 11200 7840 11212
rect 7791 11172 7840 11200
rect 7791 11169 7803 11172
rect 7745 11163 7803 11169
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 10502 11200 10508 11212
rect 8352 11172 10364 11200
rect 10415 11172 10508 11200
rect 8352 11160 8358 11172
rect 1486 11092 1492 11144
rect 1544 11132 1550 11144
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1544 11104 2145 11132
rect 1544 11092 1550 11104
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 1854 11064 1860 11076
rect 1815 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 2148 10996 2176 11095
rect 3602 11092 3608 11144
rect 3660 11132 3666 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3660 11104 4077 11132
rect 3660 11092 3666 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4396 11104 4997 11132
rect 4396 11092 4402 11104
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5350 11092 5356 11144
rect 5408 11132 5414 11144
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 5408 11104 5457 11132
rect 5408 11092 5414 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 7006 11092 7012 11144
rect 7064 11132 7070 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7064 11104 7389 11132
rect 7064 11092 7070 11104
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 7524 11104 7569 11132
rect 7524 11092 7530 11104
rect 8754 11092 8760 11144
rect 8812 11132 8818 11144
rect 9582 11132 9588 11144
rect 8812 11104 9588 11132
rect 8812 11092 8818 11104
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 3878 11064 3884 11076
rect 3620 11036 3884 11064
rect 3620 11005 3648 11036
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 5258 11064 5264 11076
rect 5219 11036 5264 11064
rect 5258 11024 5264 11036
rect 5316 11024 5322 11076
rect 6914 11064 6920 11076
rect 6875 11036 6920 11064
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 10137 11067 10195 11073
rect 10137 11064 10149 11067
rect 9456 11036 10149 11064
rect 9456 11024 9462 11036
rect 10137 11033 10149 11036
rect 10183 11033 10195 11067
rect 10336 11064 10364 11172
rect 10502 11160 10508 11172
rect 10560 11200 10566 11212
rect 11146 11200 11152 11212
rect 10560 11172 11152 11200
rect 10560 11160 10566 11172
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 10686 11132 10692 11144
rect 10647 11104 10692 11132
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 11256 11064 11284 11240
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 12952 11240 16427 11268
rect 12952 11228 12958 11240
rect 11876 11203 11934 11209
rect 11876 11169 11888 11203
rect 11922 11200 11934 11203
rect 11922 11172 13492 11200
rect 11922 11169 11934 11172
rect 11876 11163 11934 11169
rect 11330 11092 11336 11144
rect 11388 11132 11394 11144
rect 11609 11135 11667 11141
rect 11609 11132 11621 11135
rect 11388 11104 11621 11132
rect 11388 11092 11394 11104
rect 11609 11101 11621 11104
rect 11655 11101 11667 11135
rect 11609 11095 11667 11101
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12860 11104 13093 11132
rect 12860 11092 12866 11104
rect 13081 11101 13093 11104
rect 13127 11132 13139 11135
rect 13127 11104 13400 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 10336 11036 11284 11064
rect 12989 11067 13047 11073
rect 10137 11027 10195 11033
rect 12989 11033 13001 11067
rect 13035 11064 13047 11067
rect 13170 11064 13176 11076
rect 13035 11036 13176 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 3605 10999 3663 11005
rect 3605 10996 3617 10999
rect 2148 10968 3617 10996
rect 3605 10965 3617 10968
rect 3651 10965 3663 10999
rect 3605 10959 3663 10965
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 4341 10999 4399 11005
rect 4341 10996 4353 10999
rect 3752 10968 4353 10996
rect 3752 10956 3758 10968
rect 4341 10965 4353 10968
rect 4387 10996 4399 10999
rect 4430 10996 4436 11008
rect 4387 10968 4436 10996
rect 4387 10965 4399 10968
rect 4341 10959 4399 10965
rect 4430 10956 4436 10968
rect 4488 10956 4494 11008
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 4890 10996 4896 11008
rect 4580 10968 4625 10996
rect 4851 10968 4896 10996
rect 4580 10956 4586 10968
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 13262 10996 13268 11008
rect 5132 10968 13268 10996
rect 5132 10956 5138 10968
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 13372 10996 13400 11104
rect 13464 11064 13492 11172
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 14461 11203 14519 11209
rect 14461 11200 14473 11203
rect 13964 11172 14473 11200
rect 13964 11160 13970 11172
rect 14461 11169 14473 11172
rect 14507 11169 14519 11203
rect 15102 11200 15108 11212
rect 15063 11172 15108 11200
rect 14461 11163 14519 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 15729 11203 15787 11209
rect 15729 11200 15741 11203
rect 15620 11172 15741 11200
rect 15620 11160 15626 11172
rect 15729 11169 15741 11172
rect 15775 11169 15787 11203
rect 16399 11200 16427 11240
rect 16942 11200 16948 11212
rect 16399 11172 16948 11200
rect 15729 11163 15787 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17862 11200 17868 11212
rect 17823 11172 17868 11200
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 13722 11132 13728 11144
rect 13683 11104 13728 11132
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13817 11135 13875 11141
rect 13817 11101 13829 11135
rect 13863 11132 13875 11135
rect 13998 11132 14004 11144
rect 13863 11104 14004 11132
rect 13863 11101 13875 11104
rect 13817 11095 13875 11101
rect 13832 11064 13860 11095
rect 13998 11092 14004 11104
rect 14056 11132 14062 11144
rect 14645 11135 14703 11141
rect 14645 11132 14657 11135
rect 14056 11104 14657 11132
rect 14056 11092 14062 11104
rect 14645 11101 14657 11104
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 15473 11135 15531 11141
rect 15473 11132 15485 11135
rect 15068 11104 15485 11132
rect 15068 11092 15074 11104
rect 15473 11101 15485 11104
rect 15519 11101 15531 11135
rect 15473 11095 15531 11101
rect 17770 11092 17776 11144
rect 17828 11132 17834 11144
rect 18049 11135 18107 11141
rect 18049 11132 18061 11135
rect 17828 11104 18061 11132
rect 17828 11092 17834 11104
rect 18049 11101 18061 11104
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 13464 11036 13860 11064
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 15381 11067 15439 11073
rect 15381 11064 15393 11067
rect 14884 11036 15393 11064
rect 14884 11024 14890 11036
rect 15381 11033 15393 11036
rect 15427 11064 15439 11067
rect 15427 11036 15516 11064
rect 15427 11033 15439 11036
rect 15381 11027 15439 11033
rect 13814 10996 13820 11008
rect 13372 10968 13820 10996
rect 13814 10956 13820 10968
rect 13872 10956 13878 11008
rect 15488 10996 15516 11036
rect 16758 10996 16764 11008
rect 15488 10968 16764 10996
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 2225 10795 2283 10801
rect 2225 10792 2237 10795
rect 1820 10764 2237 10792
rect 1820 10752 1826 10764
rect 2225 10761 2237 10764
rect 2271 10761 2283 10795
rect 2225 10755 2283 10761
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 5074 10792 5080 10804
rect 3476 10764 5080 10792
rect 3476 10752 3482 10764
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 6178 10792 6184 10804
rect 5592 10764 5856 10792
rect 6091 10764 6184 10792
rect 5592 10752 5598 10764
rect 2958 10724 2964 10736
rect 2700 10696 2964 10724
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2700 10665 2728 10696
rect 2958 10684 2964 10696
rect 3016 10684 3022 10736
rect 5828 10724 5856 10764
rect 6178 10752 6184 10764
rect 6236 10792 6242 10804
rect 6825 10795 6883 10801
rect 6236 10764 6408 10792
rect 6236 10752 6242 10764
rect 6273 10727 6331 10733
rect 6273 10724 6285 10727
rect 5828 10696 6285 10724
rect 6273 10693 6285 10696
rect 6319 10693 6331 10727
rect 6380 10724 6408 10764
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 7006 10792 7012 10804
rect 6871 10764 7012 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 7466 10792 7472 10804
rect 7116 10764 7472 10792
rect 7116 10724 7144 10764
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 8846 10792 8852 10804
rect 8807 10764 8852 10792
rect 8846 10752 8852 10764
rect 8904 10752 8910 10804
rect 8941 10795 8999 10801
rect 8941 10761 8953 10795
rect 8987 10792 8999 10795
rect 9122 10792 9128 10804
rect 8987 10764 9128 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 17494 10792 17500 10804
rect 9600 10764 17356 10792
rect 17455 10764 17500 10792
rect 8481 10727 8539 10733
rect 8481 10724 8493 10727
rect 6380 10696 7144 10724
rect 7300 10696 8493 10724
rect 6273 10687 6331 10693
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 3786 10656 3792 10668
rect 2915 10628 3792 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 4614 10656 4620 10668
rect 4575 10628 4620 10656
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 7300 10665 7328 10696
rect 8481 10693 8493 10696
rect 8527 10724 8539 10727
rect 9600 10724 9628 10764
rect 8527 10696 9628 10724
rect 8527 10693 8539 10696
rect 8481 10687 8539 10693
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 17328 10724 17356 10764
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 17678 10724 17684 10736
rect 11388 10696 12112 10724
rect 17328 10696 17684 10724
rect 11388 10684 11394 10696
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 5868 10628 7297 10656
rect 5868 10616 5874 10628
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7558 10656 7564 10668
rect 7515 10628 7564 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8202 10656 8208 10668
rect 8163 10628 8208 10656
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 9398 10656 9404 10668
rect 9359 10628 9404 10656
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1452 10560 1777 10588
rect 1452 10548 1458 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 3050 10588 3056 10600
rect 2639 10560 3056 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 4706 10588 4712 10600
rect 4387 10560 4712 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10588 4859 10591
rect 6454 10588 6460 10600
rect 4847 10560 4927 10588
rect 6415 10560 6460 10588
rect 4847 10557 4859 10560
rect 4801 10551 4859 10557
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 2958 10520 2964 10532
rect 1903 10492 2964 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 1397 10455 1455 10461
rect 1397 10421 1409 10455
rect 1443 10452 1455 10455
rect 1670 10452 1676 10464
rect 1443 10424 1676 10452
rect 1443 10421 1455 10424
rect 1397 10415 1455 10421
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 3142 10452 3148 10464
rect 3103 10424 3148 10452
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3418 10412 3424 10464
rect 3476 10452 3482 10464
rect 3513 10455 3571 10461
rect 3513 10452 3525 10455
rect 3476 10424 3525 10452
rect 3476 10412 3482 10424
rect 3513 10421 3525 10424
rect 3559 10421 3571 10455
rect 3513 10415 3571 10421
rect 3605 10455 3663 10461
rect 3605 10421 3617 10455
rect 3651 10452 3663 10455
rect 3973 10455 4031 10461
rect 3973 10452 3985 10455
rect 3651 10424 3985 10452
rect 3651 10421 3663 10424
rect 3605 10415 3663 10421
rect 3973 10421 3985 10424
rect 4019 10421 4031 10455
rect 4430 10452 4436 10464
rect 4391 10424 4436 10452
rect 3973 10415 4031 10421
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 4899 10452 4927 10560
rect 6454 10548 6460 10560
rect 6512 10548 6518 10600
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 6972 10560 8033 10588
rect 6972 10548 6978 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 8846 10548 8852 10600
rect 8904 10588 8910 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 8904 10560 9321 10588
rect 8904 10548 8910 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 5074 10529 5080 10532
rect 5068 10520 5080 10529
rect 5035 10492 5080 10520
rect 5068 10483 5080 10492
rect 5074 10480 5080 10483
rect 5132 10480 5138 10532
rect 5166 10480 5172 10532
rect 5224 10520 5230 10532
rect 8113 10523 8171 10529
rect 8113 10520 8125 10523
rect 5224 10492 8125 10520
rect 5224 10480 5230 10492
rect 8113 10489 8125 10492
rect 8159 10489 8171 10523
rect 9600 10520 9628 10619
rect 9766 10588 9772 10600
rect 9727 10560 9772 10588
rect 9766 10548 9772 10560
rect 9824 10588 9830 10600
rect 11330 10588 11336 10600
rect 9824 10560 11336 10588
rect 9824 10548 9830 10560
rect 9674 10520 9680 10532
rect 9587 10492 9680 10520
rect 8113 10483 8171 10489
rect 9674 10480 9680 10492
rect 9732 10520 9738 10532
rect 10036 10523 10094 10529
rect 10036 10520 10048 10523
rect 9732 10492 10048 10520
rect 9732 10480 9738 10492
rect 10036 10489 10048 10492
rect 10082 10520 10094 10523
rect 10318 10520 10324 10532
rect 10082 10492 10324 10520
rect 10082 10489 10094 10492
rect 10036 10483 10094 10489
rect 10318 10480 10324 10492
rect 10376 10520 10382 10532
rect 10594 10520 10600 10532
rect 10376 10492 10600 10520
rect 10376 10480 10382 10492
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 6546 10452 6552 10464
rect 4856 10424 4927 10452
rect 6507 10424 6552 10452
rect 4856 10412 4862 10424
rect 6546 10412 6552 10424
rect 6604 10452 6610 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 6604 10424 7205 10452
rect 6604 10412 6610 10424
rect 7193 10421 7205 10424
rect 7239 10452 7251 10455
rect 7374 10452 7380 10464
rect 7239 10424 7380 10452
rect 7239 10421 7251 10424
rect 7193 10415 7251 10421
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7653 10455 7711 10461
rect 7653 10421 7665 10455
rect 7699 10452 7711 10455
rect 7834 10452 7840 10464
rect 7699 10424 7840 10452
rect 7699 10421 7711 10424
rect 7653 10415 7711 10421
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 9490 10452 9496 10464
rect 9364 10424 9496 10452
rect 9364 10412 9370 10424
rect 9490 10412 9496 10424
rect 9548 10452 9554 10464
rect 11256 10461 11284 10560
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 11425 10591 11483 10597
rect 11425 10557 11437 10591
rect 11471 10588 11483 10591
rect 11606 10588 11612 10600
rect 11471 10560 11612 10588
rect 11471 10557 11483 10560
rect 11425 10551 11483 10557
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 12084 10588 12112 10696
rect 17678 10684 17684 10696
rect 17736 10724 17742 10736
rect 18966 10724 18972 10736
rect 17736 10696 18972 10724
rect 17736 10684 17742 10696
rect 18966 10684 18972 10696
rect 19024 10684 19030 10736
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10656 12219 10659
rect 13906 10656 13912 10668
rect 12207 10628 12572 10656
rect 13867 10628 13912 10656
rect 12207 10625 12219 10628
rect 12161 10619 12219 10625
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 11940 10560 11985 10588
rect 12084 10560 12449 10588
rect 11940 10548 11946 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12544 10588 12572 10628
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 12704 10591 12762 10597
rect 12704 10588 12716 10591
rect 12544 10560 12716 10588
rect 12437 10551 12495 10557
rect 12704 10557 12716 10560
rect 12750 10588 12762 10591
rect 13170 10588 13176 10600
rect 12750 10560 13176 10588
rect 12750 10557 12762 10560
rect 12704 10551 12762 10557
rect 12158 10520 12164 10532
rect 12084 10492 12164 10520
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 9548 10424 11161 10452
rect 9548 10412 9554 10424
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11149 10415 11207 10421
rect 11241 10455 11299 10461
rect 11241 10421 11253 10455
rect 11287 10421 11299 10455
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11241 10415 11299 10421
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 11977 10455 12035 10461
rect 11977 10421 11989 10455
rect 12023 10452 12035 10455
rect 12084 10452 12112 10492
rect 12158 10480 12164 10492
rect 12216 10480 12222 10532
rect 12452 10520 12480 10551
rect 13170 10548 13176 10560
rect 13228 10548 13234 10600
rect 14274 10548 14280 10600
rect 14332 10588 14338 10600
rect 14461 10591 14519 10597
rect 14461 10588 14473 10591
rect 14332 10560 14473 10588
rect 14332 10548 14338 10560
rect 14461 10557 14473 10560
rect 14507 10588 14519 10591
rect 15010 10588 15016 10600
rect 14507 10560 15016 10588
rect 14507 10557 14519 10560
rect 14461 10551 14519 10557
rect 15010 10548 15016 10560
rect 15068 10588 15074 10600
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 15068 10560 16129 10588
rect 15068 10548 15074 10560
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 12618 10520 12624 10532
rect 12452 10492 12624 10520
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 13722 10520 13728 10532
rect 13556 10492 13728 10520
rect 12023 10424 12112 10452
rect 12023 10421 12035 10424
rect 11977 10415 12035 10421
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 13556 10452 13584 10492
rect 13722 10480 13728 10492
rect 13780 10520 13786 10532
rect 14185 10523 14243 10529
rect 14185 10520 14197 10523
rect 13780 10492 14197 10520
rect 13780 10480 13786 10492
rect 14185 10489 14197 10492
rect 14231 10489 14243 10523
rect 14185 10483 14243 10489
rect 14728 10523 14786 10529
rect 14728 10489 14740 10523
rect 14774 10520 14786 10523
rect 16384 10523 16442 10529
rect 14774 10492 16344 10520
rect 14774 10489 14786 10492
rect 14728 10483 14786 10489
rect 13814 10452 13820 10464
rect 12492 10424 13584 10452
rect 13775 10424 13820 10452
rect 12492 10412 12498 10424
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 15562 10412 15568 10464
rect 15620 10452 15626 10464
rect 15841 10455 15899 10461
rect 15841 10452 15853 10455
rect 15620 10424 15853 10452
rect 15620 10412 15626 10424
rect 15841 10421 15853 10424
rect 15887 10421 15899 10455
rect 16022 10452 16028 10464
rect 15983 10424 16028 10452
rect 15841 10415 15899 10421
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16316 10452 16344 10492
rect 16384 10489 16396 10523
rect 16430 10520 16442 10523
rect 16574 10520 16580 10532
rect 16430 10492 16580 10520
rect 16430 10489 16442 10492
rect 16384 10483 16442 10489
rect 16574 10480 16580 10492
rect 16632 10480 16638 10532
rect 16666 10452 16672 10464
rect 16316 10424 16672 10452
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2096 10220 2789 10248
rect 2096 10208 2102 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 3513 10251 3571 10257
rect 3513 10217 3525 10251
rect 3559 10248 3571 10251
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 3559 10220 4169 10248
rect 3559 10217 3571 10220
rect 3513 10211 3571 10217
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 4157 10211 4215 10217
rect 4430 10208 4436 10260
rect 4488 10248 4494 10260
rect 4985 10251 5043 10257
rect 4985 10248 4997 10251
rect 4488 10220 4997 10248
rect 4488 10208 4494 10220
rect 4985 10217 4997 10220
rect 5031 10217 5043 10251
rect 4985 10211 5043 10217
rect 5077 10251 5135 10257
rect 5077 10217 5089 10251
rect 5123 10248 5135 10251
rect 5166 10248 5172 10260
rect 5123 10220 5172 10248
rect 5123 10217 5135 10220
rect 5077 10211 5135 10217
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 5445 10251 5503 10257
rect 5445 10217 5457 10251
rect 5491 10248 5503 10251
rect 5905 10251 5963 10257
rect 5905 10248 5917 10251
rect 5491 10220 5917 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 5905 10217 5917 10220
rect 5951 10217 5963 10251
rect 6362 10248 6368 10260
rect 6323 10220 6368 10248
rect 5905 10211 5963 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 7282 10248 7288 10260
rect 6963 10220 7288 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7524 10220 7849 10248
rect 7524 10208 7530 10220
rect 7837 10217 7849 10220
rect 7883 10248 7895 10251
rect 10318 10248 10324 10260
rect 7883 10220 9628 10248
rect 10279 10220 10324 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 1664 10183 1722 10189
rect 1664 10149 1676 10183
rect 1710 10180 1722 10183
rect 2682 10180 2688 10192
rect 1710 10152 2688 10180
rect 1710 10149 1722 10152
rect 1664 10143 1722 10149
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 4338 10140 4344 10192
rect 4396 10180 4402 10192
rect 4525 10183 4583 10189
rect 4525 10180 4537 10183
rect 4396 10152 4537 10180
rect 4396 10140 4402 10152
rect 4525 10149 4537 10152
rect 4571 10149 4583 10183
rect 6178 10180 6184 10192
rect 4525 10143 4583 10149
rect 4623 10152 6184 10180
rect 2590 10072 2596 10124
rect 2648 10112 2654 10124
rect 2961 10115 3019 10121
rect 2961 10112 2973 10115
rect 2648 10084 2973 10112
rect 2648 10072 2654 10084
rect 2961 10081 2973 10084
rect 3007 10112 3019 10115
rect 3418 10112 3424 10124
rect 3007 10084 3424 10112
rect 3007 10081 3019 10084
rect 2961 10075 3019 10081
rect 3418 10072 3424 10084
rect 3476 10112 3482 10124
rect 4623 10112 4651 10152
rect 6178 10140 6184 10152
rect 6236 10180 6242 10192
rect 6273 10183 6331 10189
rect 6273 10180 6285 10183
rect 6236 10152 6285 10180
rect 6236 10140 6242 10152
rect 6273 10149 6285 10152
rect 6319 10149 6331 10183
rect 6273 10143 6331 10149
rect 7374 10140 7380 10192
rect 7432 10180 7438 10192
rect 8196 10183 8254 10189
rect 7432 10152 8156 10180
rect 7432 10140 7438 10152
rect 3476 10084 4651 10112
rect 4985 10115 5043 10121
rect 3476 10072 3482 10084
rect 4985 10081 4997 10115
rect 5031 10112 5043 10115
rect 6914 10112 6920 10124
rect 5031 10084 5856 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10013 3663 10047
rect 3786 10044 3792 10056
rect 3747 10016 3792 10044
rect 3605 10007 3663 10013
rect 3620 9976 3648 10007
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4212 10016 4629 10044
rect 4212 10004 4218 10016
rect 4430 9976 4436 9988
rect 3620 9948 4436 9976
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 3145 9911 3203 9917
rect 3145 9877 3157 9911
rect 3191 9908 3203 9911
rect 3418 9908 3424 9920
rect 3191 9880 3424 9908
rect 3191 9877 3203 9880
rect 3145 9871 3203 9877
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 4540 9908 4568 10016
rect 4617 10013 4629 10016
rect 4663 10013 4675 10047
rect 4617 10007 4675 10013
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 5534 10044 5540 10056
rect 4764 10016 4809 10044
rect 5495 10016 5540 10044
rect 4764 10004 4770 10016
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5718 10044 5724 10056
rect 5679 10016 5724 10044
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 5828 10044 5856 10084
rect 6380 10084 6920 10112
rect 6380 10044 6408 10084
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10112 7343 10115
rect 7650 10112 7656 10124
rect 7331 10084 7656 10112
rect 7331 10081 7343 10084
rect 7285 10075 7343 10081
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 7926 10112 7932 10124
rect 7887 10084 7932 10112
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 8128 10112 8156 10152
rect 8196 10149 8208 10183
rect 8242 10180 8254 10183
rect 9490 10180 9496 10192
rect 8242 10152 9496 10180
rect 8242 10149 8254 10152
rect 8196 10143 8254 10149
rect 9490 10140 9496 10152
rect 9548 10140 9554 10192
rect 9600 10180 9628 10220
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 10781 10251 10839 10257
rect 10781 10217 10793 10251
rect 10827 10248 10839 10251
rect 11514 10248 11520 10260
rect 10827 10220 11520 10248
rect 10827 10217 10839 10220
rect 10781 10211 10839 10217
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11655 10220 11989 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 11977 10217 11989 10220
rect 12023 10217 12035 10251
rect 11977 10211 12035 10217
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12124 10220 12909 10248
rect 12124 10208 12130 10220
rect 12897 10217 12909 10220
rect 12943 10248 12955 10251
rect 15102 10248 15108 10260
rect 12943 10220 15108 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15841 10251 15899 10257
rect 15841 10217 15853 10251
rect 15887 10248 15899 10251
rect 16209 10251 16267 10257
rect 16209 10248 16221 10251
rect 15887 10220 16221 10248
rect 15887 10217 15899 10220
rect 15841 10211 15899 10217
rect 16209 10217 16221 10220
rect 16255 10217 16267 10251
rect 16577 10251 16635 10257
rect 16577 10248 16589 10251
rect 16209 10211 16267 10217
rect 16316 10220 16589 10248
rect 10870 10180 10876 10192
rect 9600 10152 10876 10180
rect 10870 10140 10876 10152
rect 10928 10140 10934 10192
rect 13602 10183 13660 10189
rect 13602 10180 13614 10183
rect 10980 10152 13614 10180
rect 9398 10112 9404 10124
rect 8128 10084 8984 10112
rect 9359 10084 9404 10112
rect 5828 10016 6408 10044
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10013 6607 10047
rect 7374 10044 7380 10056
rect 7335 10016 7380 10044
rect 6549 10007 6607 10013
rect 5074 9936 5080 9988
rect 5132 9976 5138 9988
rect 6564 9976 6592 10007
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 7558 10044 7564 10056
rect 7519 10016 7564 10044
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7006 9976 7012 9988
rect 5132 9948 7012 9976
rect 5132 9936 5138 9948
rect 7006 9936 7012 9948
rect 7064 9976 7070 9988
rect 7576 9976 7604 10004
rect 7064 9948 7604 9976
rect 8956 9976 8984 10084
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 9953 10115 10011 10121
rect 9953 10081 9965 10115
rect 9999 10112 10011 10115
rect 10410 10112 10416 10124
rect 9999 10084 10416 10112
rect 9999 10081 10011 10084
rect 9953 10075 10011 10081
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 9968 10044 9996 10075
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 10735 10084 10916 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 9272 10016 9996 10044
rect 10045 10047 10103 10053
rect 9272 10004 9278 10016
rect 10045 10013 10057 10047
rect 10091 10044 10103 10047
rect 10226 10044 10232 10056
rect 10091 10016 10232 10044
rect 10091 10013 10103 10016
rect 10045 10007 10103 10013
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10686 9976 10692 9988
rect 8956 9948 10692 9976
rect 7064 9936 7070 9948
rect 10686 9936 10692 9948
rect 10744 9936 10750 9988
rect 10888 9976 10916 10084
rect 10980 10053 11008 10152
rect 13602 10149 13614 10152
rect 13648 10180 13660 10183
rect 13814 10180 13820 10192
rect 13648 10152 13820 10180
rect 13648 10149 13660 10152
rect 13602 10143 13660 10149
rect 13814 10140 13820 10152
rect 13872 10140 13878 10192
rect 13906 10140 13912 10192
rect 13964 10180 13970 10192
rect 16022 10180 16028 10192
rect 13964 10152 16028 10180
rect 13964 10140 13970 10152
rect 16022 10140 16028 10152
rect 16080 10180 16086 10192
rect 16316 10180 16344 10220
rect 16577 10217 16589 10220
rect 16623 10217 16635 10251
rect 17310 10248 17316 10260
rect 17271 10220 17316 10248
rect 16577 10211 16635 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17678 10208 17684 10260
rect 17736 10248 17742 10260
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 17736 10220 17785 10248
rect 17736 10208 17742 10220
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 16666 10180 16672 10192
rect 16080 10152 16344 10180
rect 16408 10152 16672 10180
rect 16080 10140 16086 10152
rect 11514 10112 11520 10124
rect 11475 10084 11520 10112
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 12342 10112 12348 10124
rect 12303 10084 12348 10112
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 12483 10084 12664 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 10965 10047 11023 10053
rect 10965 10013 10977 10047
rect 11011 10013 11023 10047
rect 11238 10044 11244 10056
rect 10965 10007 11023 10013
rect 11072 10016 11244 10044
rect 11072 9976 11100 10016
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 11793 10047 11851 10053
rect 11793 10013 11805 10047
rect 11839 10044 11851 10047
rect 12066 10044 12072 10056
rect 11839 10016 12072 10044
rect 11839 10013 11851 10016
rect 11793 10007 11851 10013
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12526 10044 12532 10056
rect 12487 10016 12532 10044
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 12636 10044 12664 10084
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 13081 10115 13139 10121
rect 13081 10112 13093 10115
rect 12860 10084 13093 10112
rect 12860 10072 12866 10084
rect 13081 10081 13093 10084
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 14550 10072 14556 10124
rect 14608 10112 14614 10124
rect 14921 10115 14979 10121
rect 14921 10112 14933 10115
rect 14608 10084 14933 10112
rect 14608 10072 14614 10084
rect 14921 10081 14933 10084
rect 14967 10081 14979 10115
rect 14921 10075 14979 10081
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15712 10084 15761 10112
rect 15712 10072 15718 10084
rect 15749 10081 15761 10084
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 12986 10044 12992 10056
rect 12636 10016 12992 10044
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 13262 10044 13268 10056
rect 13223 10016 13268 10044
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 16025 10047 16083 10053
rect 16025 10013 16037 10047
rect 16071 10044 16083 10047
rect 16408 10044 16436 10152
rect 16666 10140 16672 10152
rect 16724 10180 16730 10192
rect 17494 10180 17500 10192
rect 16724 10152 17500 10180
rect 16724 10140 16730 10152
rect 17494 10140 17500 10152
rect 17552 10140 17558 10192
rect 17788 10180 17816 10211
rect 17862 10208 17868 10260
rect 17920 10248 17926 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 17920 10220 18153 10248
rect 17920 10208 17926 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18141 10211 18199 10217
rect 18417 10183 18475 10189
rect 18417 10180 18429 10183
rect 17788 10152 18429 10180
rect 18417 10149 18429 10152
rect 18463 10149 18475 10183
rect 18417 10143 18475 10149
rect 17126 10072 17132 10124
rect 17184 10112 17190 10124
rect 17678 10112 17684 10124
rect 17184 10084 17684 10112
rect 17184 10072 17190 10084
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 16666 10044 16672 10056
rect 16071 10016 16436 10044
rect 16627 10016 16672 10044
rect 16071 10013 16083 10016
rect 16025 10007 16083 10013
rect 10888 9948 11100 9976
rect 11149 9979 11207 9985
rect 11149 9945 11161 9979
rect 11195 9976 11207 9979
rect 11882 9976 11888 9988
rect 11195 9948 11888 9976
rect 11195 9945 11207 9948
rect 11149 9939 11207 9945
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 12894 9936 12900 9988
rect 12952 9976 12958 9988
rect 13372 9976 13400 10007
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 17770 10044 17776 10056
rect 16899 10016 17776 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 15010 9976 15016 9988
rect 12952 9948 13400 9976
rect 14292 9948 15016 9976
rect 12952 9936 12958 9948
rect 5350 9908 5356 9920
rect 4540 9880 5356 9908
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 6733 9911 6791 9917
rect 6733 9908 6745 9911
rect 6144 9880 6745 9908
rect 6144 9868 6150 9880
rect 6733 9877 6745 9880
rect 6779 9877 6791 9911
rect 6733 9871 6791 9877
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7466 9908 7472 9920
rect 6972 9880 7472 9908
rect 6972 9868 6978 9880
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 9306 9908 9312 9920
rect 9267 9880 9312 9908
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 10410 9908 10416 9920
rect 9456 9880 10416 9908
rect 9456 9868 9462 9880
rect 10410 9868 10416 9880
rect 10468 9868 10474 9920
rect 12250 9868 12256 9920
rect 12308 9908 12314 9920
rect 14292 9908 14320 9948
rect 15010 9936 15016 9948
rect 15068 9936 15074 9988
rect 16574 9936 16580 9988
rect 16632 9976 16638 9988
rect 16868 9976 16896 10007
rect 17770 10004 17776 10016
rect 17828 10044 17834 10056
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 17828 10016 17877 10044
rect 17828 10004 17834 10016
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 17126 9976 17132 9988
rect 16632 9948 16896 9976
rect 17087 9948 17132 9976
rect 16632 9936 16638 9948
rect 17126 9936 17132 9948
rect 17184 9936 17190 9988
rect 14734 9908 14740 9920
rect 12308 9880 14320 9908
rect 14695 9880 14740 9908
rect 12308 9868 12314 9880
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 15378 9908 15384 9920
rect 15339 9880 15384 9908
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 16298 9868 16304 9920
rect 16356 9908 16362 9920
rect 18046 9908 18052 9920
rect 16356 9880 18052 9908
rect 16356 9868 16362 9880
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4801 9707 4859 9713
rect 4801 9704 4813 9707
rect 4396 9676 4813 9704
rect 4396 9664 4402 9676
rect 4801 9673 4813 9676
rect 4847 9673 4859 9707
rect 8110 9704 8116 9716
rect 4801 9667 4859 9673
rect 7208 9676 8116 9704
rect 4430 9596 4436 9648
rect 4488 9636 4494 9648
rect 4893 9639 4951 9645
rect 4893 9636 4905 9639
rect 4488 9608 4905 9636
rect 4488 9596 4494 9608
rect 4893 9605 4905 9608
rect 4939 9605 4951 9639
rect 4893 9599 4951 9605
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5905 9639 5963 9645
rect 5905 9636 5917 9639
rect 5592 9608 5917 9636
rect 5592 9596 5598 9608
rect 5905 9605 5917 9608
rect 5951 9605 5963 9639
rect 5905 9599 5963 9605
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 1949 9571 2007 9577
rect 1949 9568 1961 9571
rect 1452 9540 1961 9568
rect 1452 9528 1458 9540
rect 1949 9537 1961 9540
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9500 1547 9503
rect 1578 9500 1584 9512
rect 1535 9472 1584 9500
rect 1535 9469 1547 9472
rect 1489 9463 1547 9469
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 1964 9432 1992 9531
rect 4706 9528 4712 9580
rect 4764 9568 4770 9580
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 4764 9540 5457 9568
rect 4764 9528 4770 9540
rect 5445 9537 5457 9540
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 6178 9568 6184 9580
rect 5859 9540 6184 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9568 6607 9571
rect 7006 9568 7012 9580
rect 6595 9540 7012 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7208 9568 7236 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 11330 9704 11336 9716
rect 8904 9676 11336 9704
rect 8904 9664 8910 9676
rect 11330 9664 11336 9676
rect 11388 9664 11394 9716
rect 12250 9704 12256 9716
rect 11440 9676 12256 9704
rect 11440 9648 11468 9676
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 12452 9676 13400 9704
rect 8202 9636 8208 9648
rect 7852 9608 8208 9636
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 7208 9540 7328 9568
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2205 9503 2263 9509
rect 2205 9500 2217 9503
rect 2096 9472 2217 9500
rect 2096 9460 2102 9472
rect 2205 9469 2217 9472
rect 2251 9469 2263 9503
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 2205 9463 2263 9469
rect 3252 9472 3433 9500
rect 3252 9432 3280 9472
rect 3421 9469 3433 9472
rect 3467 9500 3479 9503
rect 4430 9500 4436 9512
rect 3467 9472 4436 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 4430 9460 4436 9472
rect 4488 9500 4494 9512
rect 4798 9500 4804 9512
rect 4488 9472 4804 9500
rect 4488 9460 4494 9472
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 5276 9472 7205 9500
rect 3694 9441 3700 9444
rect 3666 9435 3700 9441
rect 3666 9432 3678 9435
rect 1964 9404 3280 9432
rect 3344 9404 3678 9432
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 3050 9364 3056 9376
rect 1811 9336 3056 9364
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3344 9373 3372 9404
rect 3666 9401 3678 9404
rect 3752 9432 3758 9444
rect 3752 9404 3814 9432
rect 3666 9395 3700 9401
rect 3694 9392 3700 9395
rect 3752 9392 3758 9404
rect 5074 9392 5080 9444
rect 5132 9432 5138 9444
rect 5276 9441 5304 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 7300 9441 7328 9540
rect 7392 9540 7481 9568
rect 7392 9444 7420 9540
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 5261 9435 5319 9441
rect 5261 9432 5273 9435
rect 5132 9404 5273 9432
rect 5132 9392 5138 9404
rect 5261 9401 5273 9404
rect 5307 9401 5319 9435
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 5261 9395 5319 9401
rect 6104 9404 7297 9432
rect 6104 9376 6132 9404
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 7285 9395 7343 9401
rect 7374 9392 7380 9444
rect 7432 9392 7438 9444
rect 7742 9392 7748 9444
rect 7800 9432 7806 9444
rect 7852 9432 7880 9608
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 11422 9636 11428 9648
rect 8536 9608 9904 9636
rect 11383 9608 11428 9636
rect 8536 9596 8542 9608
rect 8018 9568 8024 9580
rect 7979 9540 8024 9568
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9568 8907 9571
rect 9490 9568 9496 9580
rect 8895 9540 9496 9568
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 9585 9571 9643 9577
rect 9585 9537 9597 9571
rect 9631 9568 9643 9571
rect 9674 9568 9680 9580
rect 9631 9540 9680 9568
rect 9631 9537 9643 9540
rect 9585 9531 9643 9537
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 9876 9568 9904 9608
rect 11422 9596 11428 9608
rect 11480 9596 11486 9648
rect 11517 9639 11575 9645
rect 11517 9605 11529 9639
rect 11563 9636 11575 9639
rect 11974 9636 11980 9648
rect 11563 9608 11980 9636
rect 11563 9605 11575 9608
rect 11517 9599 11575 9605
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 12452 9636 12480 9676
rect 12084 9608 12480 9636
rect 13372 9636 13400 9676
rect 14200 9676 15148 9704
rect 14200 9648 14228 9676
rect 13817 9639 13875 9645
rect 13817 9636 13829 9639
rect 13372 9608 13829 9636
rect 12084 9580 12112 9608
rect 13817 9605 13829 9608
rect 13863 9636 13875 9639
rect 13998 9636 14004 9648
rect 13863 9608 14004 9636
rect 13863 9605 13875 9608
rect 13817 9599 13875 9605
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 14182 9596 14188 9648
rect 14240 9596 14246 9648
rect 15120 9636 15148 9676
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 15841 9707 15899 9713
rect 15841 9704 15853 9707
rect 15712 9676 15853 9704
rect 15712 9664 15718 9676
rect 15841 9673 15853 9676
rect 15887 9673 15899 9707
rect 16666 9704 16672 9716
rect 16627 9676 16672 9704
rect 15841 9667 15899 9673
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 15746 9636 15752 9648
rect 15120 9608 15752 9636
rect 15746 9596 15752 9608
rect 15804 9596 15810 9648
rect 12066 9568 12072 9580
rect 9876 9540 9987 9568
rect 12027 9540 12072 9568
rect 8036 9500 8064 9528
rect 9398 9500 9404 9512
rect 8036 9472 9404 9500
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9824 9472 9873 9500
rect 9824 9460 9830 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9959 9500 9987 9540
rect 12066 9528 12072 9540
rect 12124 9528 12130 9580
rect 16485 9571 16543 9577
rect 16485 9537 16497 9571
rect 16531 9568 16543 9571
rect 16574 9568 16580 9580
rect 16531 9540 16580 9568
rect 16531 9537 16543 9540
rect 16485 9531 16543 9537
rect 16574 9528 16580 9540
rect 16632 9528 16638 9580
rect 17218 9568 17224 9580
rect 17179 9540 17224 9568
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 11606 9500 11612 9512
rect 9959 9472 11612 9500
rect 9861 9463 9919 9469
rect 7800 9404 7880 9432
rect 8573 9435 8631 9441
rect 7800 9392 7806 9404
rect 8573 9401 8585 9435
rect 8619 9432 8631 9435
rect 9674 9432 9680 9444
rect 8619 9404 9680 9432
rect 8619 9401 8631 9404
rect 8573 9395 8631 9401
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 3329 9367 3387 9373
rect 3329 9333 3341 9367
rect 3375 9333 3387 9367
rect 3329 9327 3387 9333
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 4614 9364 4620 9376
rect 4212 9336 4620 9364
rect 4212 9324 4218 9336
rect 4614 9324 4620 9336
rect 4672 9364 4678 9376
rect 5353 9367 5411 9373
rect 5353 9364 5365 9367
rect 4672 9336 5365 9364
rect 4672 9324 4678 9336
rect 5353 9333 5365 9336
rect 5399 9364 5411 9367
rect 6086 9364 6092 9376
rect 5399 9336 6092 9364
rect 5399 9333 5411 9336
rect 5353 9327 5411 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6270 9364 6276 9376
rect 6231 9336 6276 9364
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 6411 9336 6837 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6825 9333 6837 9336
rect 6871 9333 6883 9367
rect 7650 9364 7656 9376
rect 7611 9336 7656 9364
rect 6825 9327 6883 9333
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 8202 9364 8208 9376
rect 8163 9336 8208 9364
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8665 9367 8723 9373
rect 8665 9333 8677 9367
rect 8711 9364 8723 9367
rect 9033 9367 9091 9373
rect 9033 9364 9045 9367
rect 8711 9336 9045 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 9033 9333 9045 9336
rect 9079 9333 9091 9367
rect 9033 9327 9091 9333
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9493 9367 9551 9373
rect 9493 9364 9505 9367
rect 9272 9336 9505 9364
rect 9272 9324 9278 9336
rect 9493 9333 9505 9336
rect 9539 9364 9551 9367
rect 9766 9364 9772 9376
rect 9539 9336 9772 9364
rect 9539 9333 9551 9336
rect 9493 9327 9551 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 9876 9364 9904 9463
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 12158 9500 12164 9512
rect 11716 9472 12164 9500
rect 10128 9435 10186 9441
rect 10128 9401 10140 9435
rect 10174 9432 10186 9435
rect 10870 9432 10876 9444
rect 10174 9404 10876 9432
rect 10174 9401 10186 9404
rect 10128 9395 10186 9401
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 11716 9432 11744 9472
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 12710 9509 12716 9512
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12704 9463 12716 9509
rect 12768 9500 12774 9512
rect 14185 9503 14243 9509
rect 12768 9472 12804 9500
rect 11882 9432 11888 9444
rect 11020 9404 11744 9432
rect 11843 9404 11888 9432
rect 11020 9392 11026 9404
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 12452 9432 12480 9463
rect 12710 9460 12716 9463
rect 12768 9460 12774 9472
rect 14185 9469 14197 9503
rect 14231 9500 14243 9503
rect 14274 9500 14280 9512
rect 14231 9472 14280 9500
rect 14231 9469 14243 9472
rect 14185 9463 14243 9469
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 14452 9503 14510 9509
rect 14452 9469 14464 9503
rect 14498 9500 14510 9503
rect 14734 9500 14740 9512
rect 14498 9472 14740 9500
rect 14498 9469 14510 9472
rect 14452 9463 14510 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 15252 9472 16313 9500
rect 15252 9460 15258 9472
rect 16301 9469 16313 9472
rect 16347 9500 16359 9503
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 16347 9472 18061 9500
rect 16347 9469 16359 9472
rect 16301 9463 16359 9469
rect 18049 9469 18061 9472
rect 18095 9500 18107 9503
rect 18138 9500 18144 9512
rect 18095 9472 18144 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 12894 9432 12900 9444
rect 12452 9404 12900 9432
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 14001 9435 14059 9441
rect 14001 9401 14013 9435
rect 14047 9432 14059 9435
rect 17037 9435 17095 9441
rect 17037 9432 17049 9435
rect 14047 9404 17049 9432
rect 14047 9401 14059 9404
rect 14001 9395 14059 9401
rect 17037 9401 17049 9404
rect 17083 9432 17095 9435
rect 17083 9404 17816 9432
rect 17083 9401 17095 9404
rect 17037 9395 17095 9401
rect 10042 9364 10048 9376
rect 9876 9336 10048 9364
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 10594 9364 10600 9376
rect 10376 9336 10600 9364
rect 10376 9324 10382 9336
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 10744 9336 11253 9364
rect 10744 9324 10750 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11974 9364 11980 9376
rect 11935 9336 11980 9364
rect 11241 9327 11299 9333
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 12342 9324 12348 9376
rect 12400 9364 12406 9376
rect 14016 9364 14044 9395
rect 17788 9376 17816 9404
rect 12400 9336 14044 9364
rect 12400 9324 12406 9336
rect 15102 9324 15108 9376
rect 15160 9364 15166 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 15160 9336 15577 9364
rect 15160 9324 15166 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 15746 9364 15752 9376
rect 15659 9336 15752 9364
rect 15565 9327 15623 9333
rect 15746 9324 15752 9336
rect 15804 9364 15810 9376
rect 16209 9367 16267 9373
rect 16209 9364 16221 9367
rect 15804 9336 16221 9364
rect 15804 9324 15810 9336
rect 16209 9333 16221 9336
rect 16255 9364 16267 9367
rect 16666 9364 16672 9376
rect 16255 9336 16672 9364
rect 16255 9333 16267 9336
rect 16209 9327 16267 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 17126 9364 17132 9376
rect 17087 9336 17132 9364
rect 17126 9324 17132 9336
rect 17184 9364 17190 9376
rect 17497 9367 17555 9373
rect 17497 9364 17509 9367
rect 17184 9336 17509 9364
rect 17184 9324 17190 9336
rect 17497 9333 17509 9336
rect 17543 9333 17555 9367
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 17497 9327 17555 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 2590 9160 2596 9172
rect 2551 9132 2596 9160
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 2958 9160 2964 9172
rect 2919 9132 2964 9160
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 3142 9120 3148 9172
rect 3200 9160 3206 9172
rect 3329 9163 3387 9169
rect 3329 9160 3341 9163
rect 3200 9132 3341 9160
rect 3200 9120 3206 9132
rect 3329 9129 3341 9132
rect 3375 9129 3387 9163
rect 3329 9123 3387 9129
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 4154 9160 4160 9172
rect 3476 9132 3521 9160
rect 4115 9132 4160 9160
rect 3476 9120 3482 9132
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 4890 9160 4896 9172
rect 4724 9132 4896 9160
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 2501 9095 2559 9101
rect 2501 9092 2513 9095
rect 1627 9064 2513 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 2501 9061 2513 9064
rect 2547 9061 2559 9095
rect 2501 9055 2559 9061
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 9024 1731 9027
rect 1946 9024 1952 9036
rect 1719 8996 1952 9024
rect 1719 8993 1731 8996
rect 1673 8987 1731 8993
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 2516 9024 2544 9055
rect 2682 9052 2688 9104
rect 2740 9092 2746 9104
rect 4433 9095 4491 9101
rect 2740 9064 3556 9092
rect 2740 9052 2746 9064
rect 2866 9024 2872 9036
rect 2516 8996 2872 9024
rect 2866 8984 2872 8996
rect 2924 9024 2930 9036
rect 3418 9024 3424 9036
rect 2924 8996 3424 9024
rect 2924 8984 2930 8996
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 2774 8956 2780 8968
rect 2731 8928 2780 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 3528 8965 3556 9064
rect 4433 9061 4445 9095
rect 4479 9092 4491 9095
rect 4724 9092 4752 9132
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 4985 9163 5043 9169
rect 4985 9129 4997 9163
rect 5031 9160 5043 9163
rect 5166 9160 5172 9172
rect 5031 9132 5172 9160
rect 5031 9129 5043 9132
rect 4985 9123 5043 9129
rect 5166 9120 5172 9132
rect 5224 9160 5230 9172
rect 5224 9132 7512 9160
rect 5224 9120 5230 9132
rect 4479 9064 4752 9092
rect 4479 9061 4491 9064
rect 4433 9055 4491 9061
rect 4798 9052 4804 9104
rect 4856 9092 4862 9104
rect 7092 9095 7150 9101
rect 7092 9092 7104 9095
rect 4856 9064 5396 9092
rect 4856 9052 4862 9064
rect 5368 9033 5396 9064
rect 6840 9064 7104 9092
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 8993 5411 9027
rect 5353 8987 5411 8993
rect 5620 9027 5678 9033
rect 5620 8993 5632 9027
rect 5666 9024 5678 9027
rect 5994 9024 6000 9036
rect 5666 8996 6000 9024
rect 5666 8993 5678 8996
rect 5620 8987 5678 8993
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 6840 9024 6868 9064
rect 7092 9061 7104 9064
rect 7138 9092 7150 9095
rect 7374 9092 7380 9104
rect 7138 9064 7380 9092
rect 7138 9061 7150 9064
rect 7092 9055 7150 9061
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 7484 9092 7512 9132
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8260 9132 8953 9160
rect 8260 9120 8266 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 9030 9120 9036 9172
rect 9088 9160 9094 9172
rect 11790 9160 11796 9172
rect 9088 9132 9133 9160
rect 9232 9132 11796 9160
rect 9088 9120 9094 9132
rect 9232 9092 9260 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 11974 9160 11980 9172
rect 11935 9132 11980 9160
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12342 9160 12348 9172
rect 12303 9132 12348 9160
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 15194 9160 15200 9172
rect 14200 9132 15200 9160
rect 7484 9064 9260 9092
rect 9306 9052 9312 9104
rect 9364 9092 9370 9104
rect 9922 9095 9980 9101
rect 9922 9092 9934 9095
rect 9364 9064 9934 9092
rect 9364 9052 9370 9064
rect 9922 9061 9934 9064
rect 9968 9061 9980 9095
rect 9922 9055 9980 9061
rect 10042 9052 10048 9104
rect 10100 9052 10106 9104
rect 12526 9052 12532 9104
rect 12584 9092 12590 9104
rect 13265 9095 13323 9101
rect 12584 9064 12664 9092
rect 12584 9052 12590 9064
rect 7466 9024 7472 9036
rect 6748 8996 6868 9024
rect 6932 8996 7472 9024
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 1854 8820 1860 8832
rect 1815 8792 1860 8820
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 2130 8820 2136 8832
rect 2091 8792 2136 8820
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 3786 8820 3792 8832
rect 3747 8792 3792 8820
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 5184 8820 5212 8919
rect 6748 8897 6776 8996
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8956 6883 8959
rect 6932 8956 6960 8996
rect 7466 8984 7472 8996
rect 7524 9024 7530 9036
rect 7926 9024 7932 9036
rect 7524 8996 7932 9024
rect 7524 8984 7530 8996
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 8444 8996 9413 9024
rect 8444 8984 8450 8996
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 10060 9024 10088 9052
rect 9723 8996 10088 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 8294 8956 8300 8968
rect 6871 8928 6960 8956
rect 8255 8928 8300 8956
rect 6871 8925 6883 8928
rect 6825 8919 6883 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9306 8956 9312 8968
rect 9263 8928 9312 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 9416 8956 9444 8987
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11517 9027 11575 9033
rect 11517 9024 11529 9027
rect 11204 8996 11529 9024
rect 11204 8984 11210 8996
rect 11517 8993 11529 8996
rect 11563 8993 11575 9027
rect 11517 8987 11575 8993
rect 9416 8928 9536 8956
rect 6733 8891 6791 8897
rect 6733 8857 6745 8891
rect 6779 8857 6791 8891
rect 8205 8891 8263 8897
rect 8205 8888 8217 8891
rect 6733 8851 6791 8857
rect 7935 8860 8217 8888
rect 7190 8820 7196 8832
rect 5184 8792 7196 8820
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 7935 8820 7963 8860
rect 8205 8857 8217 8860
rect 8251 8857 8263 8891
rect 8205 8851 8263 8857
rect 8570 8820 8576 8832
rect 7616 8792 7963 8820
rect 8531 8792 8576 8820
rect 7616 8780 7622 8792
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 9508 8820 9536 8928
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11112 8928 11621 8956
rect 11112 8916 11118 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8925 11759 8959
rect 11701 8919 11759 8925
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 12526 8956 12532 8968
rect 12483 8928 12532 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 11716 8888 11744 8919
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 12636 8965 12664 9064
rect 13265 9061 13277 9095
rect 13311 9092 13323 9095
rect 13722 9092 13728 9104
rect 13311 9064 13728 9092
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 13170 9024 13176 9036
rect 13131 8996 13176 9024
rect 13170 8984 13176 8996
rect 13228 9024 13234 9036
rect 13630 9024 13636 9036
rect 13228 8996 13636 9024
rect 13228 8984 13234 8996
rect 13630 8984 13636 8996
rect 13688 9024 13694 9036
rect 14200 9024 14228 9132
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 15378 9120 15384 9172
rect 15436 9160 15442 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 15436 9132 15761 9160
rect 15436 9120 15442 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 15749 9123 15807 9129
rect 16022 9120 16028 9172
rect 16080 9160 16086 9172
rect 16390 9160 16396 9172
rect 16080 9132 16396 9160
rect 16080 9120 16086 9132
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 17957 9163 18015 9169
rect 17957 9160 17969 9163
rect 17920 9132 17969 9160
rect 17920 9120 17926 9132
rect 17957 9129 17969 9132
rect 18003 9129 18015 9163
rect 17957 9123 18015 9129
rect 14274 9052 14280 9104
rect 14332 9092 14338 9104
rect 15657 9095 15715 9101
rect 14332 9064 15424 9092
rect 14332 9052 14338 9064
rect 13688 8996 14228 9024
rect 13688 8984 13694 8996
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 14700 8996 14749 9024
rect 14700 8984 14706 8996
rect 14737 8993 14749 8996
rect 14783 9024 14795 9027
rect 15396 9024 15424 9064
rect 15657 9061 15669 9095
rect 15703 9092 15715 9095
rect 16114 9092 16120 9104
rect 15703 9064 16120 9092
rect 15703 9061 15715 9064
rect 15657 9055 15715 9061
rect 16114 9052 16120 9064
rect 16172 9052 16178 9104
rect 16844 9095 16902 9101
rect 16844 9061 16856 9095
rect 16890 9092 16902 9095
rect 17218 9092 17224 9104
rect 16890 9064 17224 9092
rect 16890 9061 16902 9064
rect 16844 9055 16902 9061
rect 17218 9052 17224 9064
rect 17276 9052 17282 9104
rect 16390 9024 16396 9036
rect 14783 8996 15056 9024
rect 15396 8996 16396 9024
rect 14783 8993 14795 8996
rect 14737 8987 14795 8993
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8956 12679 8959
rect 12710 8956 12716 8968
rect 12667 8928 12716 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 12710 8916 12716 8928
rect 12768 8956 12774 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 12768 8928 13369 8956
rect 12768 8916 12774 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 14826 8956 14832 8968
rect 14323 8928 14832 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 14921 8959 14979 8965
rect 14921 8925 14933 8959
rect 14967 8925 14979 8959
rect 15028 8956 15056 8996
rect 16390 8984 16396 8996
rect 16448 9024 16454 9036
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 16448 8996 16589 9024
rect 16448 8984 16454 8996
rect 16577 8993 16589 8996
rect 16623 8993 16635 9027
rect 16577 8987 16635 8993
rect 16666 8984 16672 9036
rect 16724 9024 16730 9036
rect 18049 9027 18107 9033
rect 18049 9024 18061 9027
rect 16724 8996 18061 9024
rect 16724 8984 16730 8996
rect 18049 8993 18061 8996
rect 18095 9024 18107 9027
rect 18417 9027 18475 9033
rect 18417 9024 18429 9027
rect 18095 8996 18429 9024
rect 18095 8993 18107 8996
rect 18049 8987 18107 8993
rect 18417 8993 18429 8996
rect 18463 8993 18475 9027
rect 18417 8987 18475 8993
rect 15470 8956 15476 8968
rect 15028 8928 15476 8956
rect 14921 8919 14979 8925
rect 14001 8891 14059 8897
rect 14001 8888 14013 8891
rect 10744 8860 11744 8888
rect 13372 8860 14013 8888
rect 10744 8848 10750 8860
rect 13372 8832 13400 8860
rect 14001 8857 14013 8860
rect 14047 8888 14059 8891
rect 14458 8888 14464 8900
rect 14047 8860 14464 8888
rect 14047 8857 14059 8860
rect 14001 8851 14059 8857
rect 14458 8848 14464 8860
rect 14516 8848 14522 8900
rect 14734 8848 14740 8900
rect 14792 8888 14798 8900
rect 14936 8888 14964 8919
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 15562 8916 15568 8968
rect 15620 8956 15626 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 15620 8928 15853 8956
rect 15620 8916 15626 8928
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 14792 8860 14964 8888
rect 14792 8848 14798 8860
rect 15378 8848 15384 8900
rect 15436 8888 15442 8900
rect 16301 8891 16359 8897
rect 16301 8888 16313 8891
rect 15436 8860 16313 8888
rect 15436 8848 15442 8860
rect 16301 8857 16313 8860
rect 16347 8857 16359 8891
rect 16301 8851 16359 8857
rect 10594 8820 10600 8832
rect 9508 8792 10600 8820
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10928 8792 11069 8820
rect 10928 8780 10934 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8820 11207 8823
rect 11790 8820 11796 8832
rect 11195 8792 11796 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 11882 8780 11888 8832
rect 11940 8820 11946 8832
rect 12805 8823 12863 8829
rect 12805 8820 12817 8823
rect 11940 8792 12817 8820
rect 11940 8780 11946 8792
rect 12805 8789 12817 8792
rect 12851 8789 12863 8823
rect 12805 8783 12863 8789
rect 13354 8780 13360 8832
rect 13412 8780 13418 8832
rect 13630 8820 13636 8832
rect 13591 8792 13636 8820
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14182 8820 14188 8832
rect 13872 8792 14188 8820
rect 13872 8780 13878 8792
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 14369 8823 14427 8829
rect 14369 8789 14381 8823
rect 14415 8820 14427 8823
rect 14550 8820 14556 8832
rect 14415 8792 14556 8820
rect 14415 8789 14427 8792
rect 14369 8783 14427 8789
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 15286 8820 15292 8832
rect 15247 8792 15292 8820
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 16209 8823 16267 8829
rect 16209 8820 16221 8823
rect 15528 8792 16221 8820
rect 15528 8780 15534 8792
rect 16209 8789 16221 8792
rect 16255 8820 16267 8823
rect 16574 8820 16580 8832
rect 16255 8792 16580 8820
rect 16255 8789 16267 8792
rect 16209 8783 16267 8789
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 18233 8823 18291 8829
rect 18233 8789 18245 8823
rect 18279 8820 18291 8823
rect 18322 8820 18328 8832
rect 18279 8792 18328 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 2958 8616 2964 8628
rect 2648 8588 2964 8616
rect 2648 8576 2654 8588
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 4430 8576 4436 8628
rect 4488 8576 4494 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 6089 8619 6147 8625
rect 6089 8616 6101 8619
rect 5408 8588 6101 8616
rect 5408 8576 5414 8588
rect 6089 8585 6101 8588
rect 6135 8616 6147 8619
rect 6270 8616 6276 8628
rect 6135 8588 6276 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 10321 8619 10379 8625
rect 10321 8616 10333 8619
rect 7576 8588 10333 8616
rect 3418 8508 3424 8560
rect 3476 8548 3482 8560
rect 4157 8551 4215 8557
rect 4157 8548 4169 8551
rect 3476 8520 4169 8548
rect 3476 8508 3482 8520
rect 4157 8517 4169 8520
rect 4203 8517 4215 8551
rect 4157 8511 4215 8517
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 3694 8480 3700 8492
rect 3655 8452 3700 8480
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 4448 8480 4476 8576
rect 5718 8508 5724 8560
rect 5776 8548 5782 8560
rect 6454 8548 6460 8560
rect 5776 8520 6460 8548
rect 5776 8508 5782 8520
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 7576 8548 7604 8588
rect 10321 8585 10333 8588
rect 10367 8585 10379 8619
rect 10321 8579 10379 8585
rect 11977 8619 12035 8625
rect 11977 8585 11989 8619
rect 12023 8616 12035 8619
rect 12618 8616 12624 8628
rect 12023 8588 12624 8616
rect 12023 8585 12035 8588
rect 11977 8579 12035 8585
rect 6656 8520 7604 8548
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4448 8452 4629 8480
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5684 8452 6592 8480
rect 5684 8440 5690 8452
rect 2774 8372 2780 8424
rect 2832 8372 2838 8424
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3605 8415 3663 8421
rect 3605 8412 3617 8415
rect 3016 8384 3617 8412
rect 3016 8372 3022 8384
rect 3605 8381 3617 8384
rect 3651 8381 3663 8415
rect 3970 8412 3976 8424
rect 3931 8384 3976 8412
rect 3605 8375 3663 8381
rect 1664 8347 1722 8353
rect 1664 8313 1676 8347
rect 1710 8344 1722 8347
rect 2792 8344 2820 8372
rect 3418 8344 3424 8356
rect 1710 8316 3424 8344
rect 1710 8313 1722 8316
rect 1664 8307 1722 8313
rect 3418 8304 3424 8316
rect 3476 8304 3482 8356
rect 3620 8344 3648 8375
rect 3970 8372 3976 8384
rect 4028 8372 4034 8424
rect 4884 8415 4942 8421
rect 4884 8381 4896 8415
rect 4930 8412 4942 8415
rect 5810 8412 5816 8424
rect 4930 8384 5816 8412
rect 4930 8381 4942 8384
rect 4884 8375 4942 8381
rect 5810 8372 5816 8384
rect 5868 8372 5874 8424
rect 6454 8344 6460 8356
rect 3620 8316 6460 8344
rect 6454 8304 6460 8316
rect 6512 8304 6518 8356
rect 6564 8344 6592 8452
rect 6656 8421 6684 8520
rect 7006 8480 7012 8492
rect 6967 8452 7012 8480
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7524 8452 7573 8480
rect 7524 8440 7530 8452
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 10134 8480 10140 8492
rect 8812 8452 10140 8480
rect 8812 8440 8818 8452
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7817 8415 7875 8421
rect 7817 8412 7829 8415
rect 7248 8384 7829 8412
rect 7248 8372 7254 8384
rect 7817 8381 7829 8384
rect 7863 8412 7875 8415
rect 10336 8412 10364 8579
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 17218 8616 17224 8628
rect 17179 8588 17224 8616
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 11149 8551 11207 8557
rect 11149 8517 11161 8551
rect 11195 8548 11207 8551
rect 11790 8548 11796 8560
rect 11195 8520 11796 8548
rect 11195 8517 11207 8520
rect 11149 8511 11207 8517
rect 11790 8508 11796 8520
rect 11848 8508 11854 8560
rect 12437 8551 12495 8557
rect 12437 8517 12449 8551
rect 12483 8548 12495 8551
rect 13170 8548 13176 8560
rect 12483 8520 13176 8548
rect 12483 8517 12495 8520
rect 12437 8511 12495 8517
rect 13170 8508 13176 8520
rect 13228 8508 13234 8560
rect 14093 8551 14151 8557
rect 14093 8548 14105 8551
rect 13740 8520 14105 8548
rect 10502 8440 10508 8492
rect 10560 8480 10566 8492
rect 11054 8480 11060 8492
rect 10560 8452 11060 8480
rect 10560 8440 10566 8452
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 11514 8440 11520 8492
rect 11572 8480 11578 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11572 8452 11713 8480
rect 11572 8440 11578 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 12250 8480 12256 8492
rect 12032 8452 12256 8480
rect 12032 8440 12038 8452
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 13740 8489 13768 8520
rect 14093 8517 14105 8520
rect 14139 8517 14151 8551
rect 14093 8511 14151 8517
rect 14182 8508 14188 8560
rect 14240 8548 14246 8560
rect 14921 8551 14979 8557
rect 14240 8520 14780 8548
rect 14240 8508 14246 8520
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8449 13783 8483
rect 13906 8480 13912 8492
rect 13867 8452 13912 8480
rect 13725 8443 13783 8449
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 7863 8384 10272 8412
rect 10336 8384 12173 8412
rect 7863 8381 7875 8384
rect 7817 8375 7875 8381
rect 6730 8344 6736 8356
rect 6564 8316 6736 8344
rect 6730 8304 6736 8316
rect 6788 8344 6794 8356
rect 6825 8347 6883 8353
rect 6825 8344 6837 8347
rect 6788 8316 6837 8344
rect 6788 8304 6794 8316
rect 6825 8313 6837 8316
rect 6871 8313 6883 8347
rect 7466 8344 7472 8356
rect 7379 8316 7472 8344
rect 6825 8307 6883 8313
rect 7466 8304 7472 8316
rect 7524 8344 7530 8356
rect 8662 8344 8668 8356
rect 7524 8316 8668 8344
rect 7524 8304 7530 8316
rect 8662 8304 8668 8316
rect 8720 8304 8726 8356
rect 9030 8344 9036 8356
rect 8991 8316 9036 8344
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 10244 8344 10272 8384
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 13096 8412 13124 8443
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 14550 8480 14556 8492
rect 14511 8452 14556 8480
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14752 8489 14780 8520
rect 14921 8517 14933 8551
rect 14967 8548 14979 8551
rect 15654 8548 15660 8560
rect 14967 8520 15660 8548
rect 14967 8517 14979 8520
rect 14921 8511 14979 8517
rect 15654 8508 15660 8520
rect 15712 8508 15718 8560
rect 17862 8508 17868 8560
rect 17920 8548 17926 8560
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 17920 8520 18245 8548
rect 17920 8508 17926 8520
rect 18233 8517 18245 8520
rect 18279 8517 18291 8551
rect 18233 8511 18291 8517
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8480 14795 8483
rect 15102 8480 15108 8492
rect 14783 8452 15108 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 15102 8440 15108 8452
rect 15160 8480 15166 8492
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15160 8452 15485 8480
rect 15160 8440 15166 8452
rect 15473 8449 15485 8452
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 15562 8440 15568 8492
rect 15620 8480 15626 8492
rect 15620 8452 15884 8480
rect 15620 8440 15626 8452
rect 15856 8421 15884 8452
rect 15841 8415 15899 8421
rect 13096 8384 15608 8412
rect 12161 8375 12219 8381
rect 10686 8344 10692 8356
rect 10244 8316 10692 8344
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 11057 8347 11115 8353
rect 11057 8313 11069 8347
rect 11103 8344 11115 8347
rect 11422 8344 11428 8356
rect 11103 8316 11428 8344
rect 11103 8313 11115 8316
rect 11057 8307 11115 8313
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 2866 8276 2872 8288
rect 2823 8248 2872 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3142 8276 3148 8288
rect 3103 8248 3148 8276
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 3513 8279 3571 8285
rect 3513 8245 3525 8279
rect 3559 8276 3571 8279
rect 3694 8276 3700 8288
rect 3559 8248 3700 8276
rect 3559 8245 3571 8248
rect 3513 8239 3571 8245
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 4246 8236 4252 8288
rect 4304 8276 4310 8288
rect 4341 8279 4399 8285
rect 4341 8276 4353 8279
rect 4304 8248 4353 8276
rect 4304 8236 4310 8248
rect 4341 8245 4353 8248
rect 4387 8245 4399 8279
rect 5994 8276 6000 8288
rect 5955 8248 6000 8276
rect 4341 8239 4399 8245
rect 5994 8236 6000 8248
rect 6052 8236 6058 8288
rect 6270 8276 6276 8288
rect 6231 8248 6276 8276
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 7285 8279 7343 8285
rect 7285 8245 7297 8279
rect 7331 8276 7343 8279
rect 8386 8276 8392 8288
rect 7331 8248 8392 8276
rect 7331 8245 7343 8248
rect 7285 8239 7343 8245
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 8938 8276 8944 8288
rect 8899 8248 8944 8276
rect 8938 8236 8944 8248
rect 8996 8236 9002 8288
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 11072 8276 11100 8307
rect 11422 8304 11428 8316
rect 11480 8344 11486 8356
rect 12526 8344 12532 8356
rect 11480 8316 12532 8344
rect 11480 8304 11486 8316
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 12805 8347 12863 8353
rect 12805 8313 12817 8347
rect 12851 8344 12863 8347
rect 13633 8347 13691 8353
rect 12851 8316 13584 8344
rect 12851 8313 12863 8316
rect 12805 8307 12863 8313
rect 9272 8248 11100 8276
rect 9272 8236 9278 8248
rect 11238 8236 11244 8288
rect 11296 8276 11302 8288
rect 11517 8279 11575 8285
rect 11517 8276 11529 8279
rect 11296 8248 11529 8276
rect 11296 8236 11302 8248
rect 11517 8245 11529 8248
rect 11563 8245 11575 8279
rect 11517 8239 11575 8245
rect 11606 8236 11612 8288
rect 11664 8276 11670 8288
rect 12897 8279 12955 8285
rect 11664 8248 11709 8276
rect 11664 8236 11670 8248
rect 12897 8245 12909 8279
rect 12943 8276 12955 8279
rect 13265 8279 13323 8285
rect 13265 8276 13277 8279
rect 12943 8248 13277 8276
rect 12943 8245 12955 8248
rect 12897 8239 12955 8245
rect 13265 8245 13277 8248
rect 13311 8245 13323 8279
rect 13556 8276 13584 8316
rect 13633 8313 13645 8347
rect 13679 8344 13691 8347
rect 14182 8344 14188 8356
rect 13679 8316 14188 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 14182 8304 14188 8316
rect 14240 8304 14246 8356
rect 14918 8304 14924 8356
rect 14976 8344 14982 8356
rect 15289 8347 15347 8353
rect 15289 8344 15301 8347
rect 14976 8316 15301 8344
rect 14976 8304 14982 8316
rect 15289 8313 15301 8316
rect 15335 8313 15347 8347
rect 15289 8307 15347 8313
rect 15378 8304 15384 8356
rect 15436 8344 15442 8356
rect 15580 8344 15608 8384
rect 15841 8381 15853 8415
rect 15887 8412 15899 8415
rect 16390 8412 16396 8424
rect 15887 8384 16396 8412
rect 15887 8381 15899 8384
rect 15841 8375 15899 8381
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 17678 8372 17684 8424
rect 17736 8412 17742 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17736 8384 18061 8412
rect 17736 8372 17742 8384
rect 18049 8381 18061 8384
rect 18095 8412 18107 8415
rect 18417 8415 18475 8421
rect 18417 8412 18429 8415
rect 18095 8384 18429 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18417 8381 18429 8384
rect 18463 8381 18475 8415
rect 18417 8375 18475 8381
rect 16086 8347 16144 8353
rect 16086 8344 16098 8347
rect 15436 8316 15481 8344
rect 15580 8316 16098 8344
rect 15436 8304 15442 8316
rect 16086 8313 16098 8316
rect 16132 8344 16144 8347
rect 16666 8344 16672 8356
rect 16132 8316 16672 8344
rect 16132 8313 16144 8316
rect 16086 8307 16144 8313
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 14366 8276 14372 8288
rect 13556 8248 14372 8276
rect 13265 8239 13323 8245
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 14516 8248 14561 8276
rect 14516 8236 14522 8248
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 2188 8044 2329 8072
rect 2188 8032 2194 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 2317 8035 2375 8041
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2455 8044 2789 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 2777 8035 2835 8041
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 3237 8075 3295 8081
rect 3237 8072 3249 8075
rect 3200 8044 3249 8072
rect 3200 8032 3206 8044
rect 3237 8041 3249 8044
rect 3283 8041 3295 8075
rect 3786 8072 3792 8084
rect 3747 8044 3792 8072
rect 3237 8035 3295 8041
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4396 8044 4445 8072
rect 4396 8032 4402 8044
rect 4433 8041 4445 8044
rect 4479 8072 4491 8075
rect 4798 8072 4804 8084
rect 4479 8044 4804 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 5166 8072 5172 8084
rect 5127 8044 5172 8072
rect 5166 8032 5172 8044
rect 5224 8072 5230 8084
rect 5353 8075 5411 8081
rect 5353 8072 5365 8075
rect 5224 8044 5365 8072
rect 5224 8032 5230 8044
rect 5353 8041 5365 8044
rect 5399 8041 5411 8075
rect 5353 8035 5411 8041
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 8665 8075 8723 8081
rect 8665 8072 8677 8075
rect 5583 8044 8677 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 8665 8041 8677 8044
rect 8711 8041 8723 8075
rect 9674 8072 9680 8084
rect 9635 8044 9680 8072
rect 8665 8035 8723 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10226 8072 10232 8084
rect 10091 8044 10232 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 10502 8072 10508 8084
rect 10463 8044 10508 8072
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10652 8044 10885 8072
rect 10652 8032 10658 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 10965 8075 11023 8081
rect 10965 8041 10977 8075
rect 11011 8072 11023 8075
rect 11422 8072 11428 8084
rect 11011 8044 11428 8072
rect 11011 8041 11023 8044
rect 10965 8035 11023 8041
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 12710 8072 12716 8084
rect 12671 8044 12716 8072
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 16666 8072 16672 8084
rect 16627 8044 16672 8072
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 1489 8007 1547 8013
rect 1489 7973 1501 8007
rect 1535 8004 1547 8007
rect 5626 8004 5632 8016
rect 1535 7976 3188 8004
rect 1535 7973 1547 7976
rect 1489 7967 1547 7973
rect 1578 7936 1584 7948
rect 1539 7908 1584 7936
rect 1578 7896 1584 7908
rect 1636 7896 1642 7948
rect 3160 7945 3188 7976
rect 3620 7976 5632 8004
rect 3620 7945 3648 7976
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 5810 7964 5816 8016
rect 5868 8004 5874 8016
rect 6457 8007 6515 8013
rect 5868 7976 6132 8004
rect 5868 7964 5874 7976
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 3605 7939 3663 7945
rect 3191 7908 3556 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 3528 7880 3556 7908
rect 3605 7905 3617 7939
rect 3651 7905 3663 7939
rect 3605 7899 3663 7905
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 4525 7939 4583 7945
rect 4525 7936 4537 7939
rect 4396 7908 4537 7936
rect 4396 7896 4402 7908
rect 4525 7905 4537 7908
rect 4571 7936 4583 7939
rect 4571 7908 4752 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2866 7868 2872 7880
rect 2639 7840 2872 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 3418 7868 3424 7880
rect 3331 7840 3424 7868
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3694 7868 3700 7880
rect 3568 7840 3700 7868
rect 3568 7828 3574 7840
rect 3694 7828 3700 7840
rect 3752 7828 3758 7880
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4488 7840 4629 7868
rect 4488 7828 4494 7840
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 3436 7800 3464 7828
rect 3602 7800 3608 7812
rect 3436 7772 3608 7800
rect 3602 7760 3608 7772
rect 3660 7800 3666 7812
rect 4448 7800 4476 7828
rect 3660 7772 4476 7800
rect 4724 7800 4752 7908
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 5905 7939 5963 7945
rect 5905 7936 5917 7939
rect 5592 7908 5917 7936
rect 5592 7896 5598 7908
rect 5905 7905 5917 7908
rect 5951 7905 5963 7939
rect 5905 7899 5963 7905
rect 5994 7868 6000 7880
rect 5955 7840 6000 7868
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6104 7877 6132 7976
rect 6457 7973 6469 8007
rect 6503 8004 6515 8007
rect 6638 8004 6644 8016
rect 6503 7976 6644 8004
rect 6503 7973 6515 7976
rect 6457 7967 6515 7973
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 7837 8007 7895 8013
rect 7837 8004 7849 8007
rect 6788 7976 7849 8004
rect 6788 7964 6794 7976
rect 7837 7973 7849 7976
rect 7883 8004 7895 8007
rect 8294 8004 8300 8016
rect 7883 7976 8300 8004
rect 7883 7973 7895 7976
rect 7837 7967 7895 7973
rect 8294 7964 8300 7976
rect 8352 8004 8358 8016
rect 9125 8007 9183 8013
rect 8352 7976 8708 8004
rect 8352 7964 8358 7976
rect 6656 7936 6684 7964
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6656 7908 6929 7936
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7936 7067 7939
rect 7466 7936 7472 7948
rect 7055 7908 7472 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7708 7908 7757 7936
rect 7708 7896 7714 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 7745 7899 7803 7905
rect 8018 7896 8024 7948
rect 8076 7936 8082 7948
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 8076 7908 8585 7936
rect 8076 7896 8082 7908
rect 8573 7905 8585 7908
rect 8619 7905 8631 7939
rect 8680 7936 8708 7976
rect 9125 7973 9137 8007
rect 9171 8004 9183 8007
rect 9171 7976 10640 8004
rect 9171 7973 9183 7976
rect 9125 7967 9183 7973
rect 10137 7939 10195 7945
rect 10137 7936 10149 7939
rect 8680 7908 10149 7936
rect 8573 7899 8631 7905
rect 10137 7905 10149 7908
rect 10183 7936 10195 7939
rect 10502 7936 10508 7948
rect 10183 7908 10508 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 10612 7936 10640 7976
rect 11514 7964 11520 8016
rect 11572 8013 11578 8016
rect 11572 8007 11636 8013
rect 11572 7973 11590 8007
rect 11624 7973 11636 8007
rect 11572 7967 11636 7973
rect 11572 7964 11578 7967
rect 14918 7964 14924 8016
rect 14976 8004 14982 8016
rect 17681 8007 17739 8013
rect 17681 8004 17693 8007
rect 14976 7976 17693 8004
rect 14976 7964 14982 7976
rect 17681 7973 17693 7976
rect 17727 7973 17739 8007
rect 17681 7967 17739 7973
rect 11422 7936 11428 7948
rect 10612 7908 11428 7936
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7936 13323 7939
rect 13354 7936 13360 7948
rect 13311 7908 13360 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 13532 7939 13590 7945
rect 13532 7905 13544 7939
rect 13578 7936 13590 7939
rect 13814 7936 13820 7948
rect 13578 7908 13820 7936
rect 13578 7905 13590 7908
rect 13532 7899 13590 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 15556 7939 15614 7945
rect 15556 7936 15568 7939
rect 13964 7908 15568 7936
rect 13964 7896 13970 7908
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7868 7251 7871
rect 7926 7868 7932 7880
rect 7239 7840 7932 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 8754 7868 8760 7880
rect 8715 7840 8760 7868
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 10318 7868 10324 7880
rect 10279 7840 10324 7868
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10410 7828 10416 7880
rect 10468 7868 10474 7880
rect 11054 7868 11060 7880
rect 10468 7840 11060 7868
rect 10468 7828 10474 7840
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 5258 7800 5264 7812
rect 4724 7772 5264 7800
rect 3660 7760 3666 7772
rect 5258 7760 5264 7772
rect 5316 7800 5322 7812
rect 5316 7772 6684 7800
rect 5316 7760 5322 7772
rect 1762 7732 1768 7744
rect 1723 7704 1768 7732
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7732 2007 7735
rect 2130 7732 2136 7744
rect 1995 7704 2136 7732
rect 1995 7701 2007 7704
rect 1949 7695 2007 7701
rect 2130 7692 2136 7704
rect 2188 7692 2194 7744
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 3384 7704 4077 7732
rect 3384 7692 3390 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 4856 7704 4997 7732
rect 4856 7692 4862 7704
rect 4985 7701 4997 7704
rect 5031 7732 5043 7735
rect 6178 7732 6184 7744
rect 5031 7704 6184 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 6546 7732 6552 7744
rect 6507 7704 6552 7732
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 6656 7732 6684 7772
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 7377 7803 7435 7809
rect 7377 7800 7389 7803
rect 7064 7772 7389 7800
rect 7064 7760 7070 7772
rect 7377 7769 7389 7772
rect 7423 7769 7435 7803
rect 10042 7800 10048 7812
rect 7377 7763 7435 7769
rect 7484 7772 10048 7800
rect 7484 7732 7512 7772
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 8202 7732 8208 7744
rect 6656 7704 7512 7732
rect 8163 7704 8208 7732
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 9214 7732 9220 7744
rect 8352 7704 9220 7732
rect 8352 7692 8358 7704
rect 9214 7692 9220 7704
rect 9272 7732 9278 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 9272 7704 9413 7732
rect 9272 7692 9278 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 10962 7732 10968 7744
rect 9548 7704 10968 7732
rect 9548 7692 9554 7704
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11348 7732 11376 7831
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 12805 7871 12863 7877
rect 12805 7868 12817 7871
rect 12400 7840 12817 7868
rect 12400 7828 12406 7840
rect 12805 7837 12817 7840
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 14660 7809 14688 7908
rect 15556 7905 15568 7908
rect 15602 7936 15614 7939
rect 16390 7936 16396 7948
rect 15602 7908 16396 7936
rect 15602 7905 15614 7908
rect 15556 7899 15614 7905
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 17696 7936 17724 7967
rect 17865 7939 17923 7945
rect 17865 7936 17877 7939
rect 17696 7908 17877 7936
rect 17865 7905 17877 7908
rect 17911 7905 17923 7939
rect 17865 7899 17923 7905
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 14645 7803 14703 7809
rect 14645 7769 14657 7803
rect 14691 7769 14703 7803
rect 14645 7763 14703 7769
rect 11112 7704 11376 7732
rect 11112 7692 11118 7704
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 13173 7735 13231 7741
rect 13173 7732 13185 7735
rect 12860 7704 13185 7732
rect 12860 7692 12866 7704
rect 13173 7701 13185 7704
rect 13219 7732 13231 7735
rect 14274 7732 14280 7744
rect 13219 7704 14280 7732
rect 13219 7701 13231 7704
rect 13173 7695 13231 7701
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 14734 7732 14740 7744
rect 14608 7704 14740 7732
rect 14608 7692 14614 7704
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 14918 7732 14924 7744
rect 14879 7704 14924 7732
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15304 7732 15332 7831
rect 18046 7800 18052 7812
rect 18007 7772 18052 7800
rect 18046 7760 18052 7772
rect 18104 7760 18110 7812
rect 15562 7732 15568 7744
rect 15304 7704 15568 7732
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 3421 7531 3479 7537
rect 3421 7497 3433 7531
rect 3467 7528 3479 7531
rect 5166 7528 5172 7540
rect 3467 7500 5172 7528
rect 3467 7497 3479 7500
rect 3421 7491 3479 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 6273 7531 6331 7537
rect 6273 7528 6285 7531
rect 5868 7500 6285 7528
rect 5868 7488 5874 7500
rect 6273 7497 6285 7500
rect 6319 7497 6331 7531
rect 6273 7491 6331 7497
rect 6825 7531 6883 7537
rect 6825 7497 6837 7531
rect 6871 7528 6883 7531
rect 8018 7528 8024 7540
rect 6871 7500 8024 7528
rect 6871 7497 6883 7500
rect 6825 7491 6883 7497
rect 1489 7463 1547 7469
rect 1489 7429 1501 7463
rect 1535 7460 1547 7463
rect 1578 7460 1584 7472
rect 1535 7432 1584 7460
rect 1535 7429 1547 7432
rect 1489 7423 1547 7429
rect 1578 7420 1584 7432
rect 1636 7420 1642 7472
rect 6288 7460 6316 7491
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 11238 7528 11244 7540
rect 10735 7500 11244 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 12437 7531 12495 7537
rect 12437 7528 12449 7531
rect 11992 7500 12449 7528
rect 9861 7463 9919 7469
rect 6288 7432 7420 7460
rect 3421 7395 3479 7401
rect 3421 7392 3433 7395
rect 3068 7364 3433 7392
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7324 1639 7327
rect 2406 7324 2412 7336
rect 1627 7296 2412 7324
rect 1627 7293 1639 7296
rect 1581 7287 1639 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 3068 7333 3096 7364
rect 3421 7361 3433 7364
rect 3467 7361 3479 7395
rect 3421 7355 3479 7361
rect 3602 7352 3608 7404
rect 3660 7392 3666 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 3660 7364 4077 7392
rect 3660 7352 3666 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4890 7392 4896 7404
rect 4851 7364 4896 7392
rect 4065 7355 4123 7361
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 6454 7392 6460 7404
rect 6415 7364 6460 7392
rect 6454 7352 6460 7364
rect 6512 7352 6518 7404
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 7392 7401 7420 7432
rect 9861 7429 9873 7463
rect 9907 7460 9919 7463
rect 11054 7460 11060 7472
rect 9907 7432 11060 7460
rect 9907 7429 9919 7432
rect 9861 7423 9919 7429
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 11992 7460 12020 7500
rect 12437 7497 12449 7500
rect 12483 7497 12495 7531
rect 14182 7528 14188 7540
rect 14143 7500 14188 7528
rect 12437 7491 12495 7497
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 14366 7488 14372 7540
rect 14424 7528 14430 7540
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 14424 7500 15853 7528
rect 14424 7488 14430 7500
rect 15841 7497 15853 7500
rect 15887 7497 15899 7531
rect 15841 7491 15899 7497
rect 16482 7488 16488 7540
rect 16540 7528 16546 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 16540 7500 16681 7528
rect 16540 7488 16546 7500
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 16669 7491 16727 7497
rect 11155 7432 12020 7460
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 6604 7364 7297 7392
rect 6604 7352 6610 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 7377 7355 7435 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 8036 7364 8248 7392
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7324 3939 7327
rect 4246 7324 4252 7336
rect 3927 7296 4252 7324
rect 3927 7293 3939 7296
rect 3881 7287 3939 7293
rect 4246 7284 4252 7296
rect 4304 7284 4310 7336
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7324 4399 7327
rect 6270 7324 6276 7336
rect 4387 7296 6276 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 6270 7284 6276 7296
rect 6328 7284 6334 7336
rect 6362 7284 6368 7336
rect 6420 7324 6426 7336
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6420 7296 6653 7324
rect 6420 7284 6426 7296
rect 6641 7293 6653 7296
rect 6687 7293 6699 7327
rect 6641 7287 6699 7293
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 7064 7296 7205 7324
rect 7064 7284 7070 7296
rect 7193 7293 7205 7296
rect 7239 7293 7251 7327
rect 8036 7324 8064 7364
rect 7193 7287 7251 7293
rect 7576 7296 8064 7324
rect 8113 7327 8171 7333
rect 1848 7259 1906 7265
rect 1848 7225 1860 7259
rect 1894 7256 1906 7259
rect 2866 7256 2872 7268
rect 1894 7228 2872 7256
rect 1894 7225 1906 7228
rect 1848 7219 1906 7225
rect 2866 7216 2872 7228
rect 2924 7256 2930 7268
rect 3418 7256 3424 7268
rect 2924 7228 3424 7256
rect 2924 7216 2930 7228
rect 3418 7216 3424 7228
rect 3476 7216 3482 7268
rect 3973 7259 4031 7265
rect 3973 7225 3985 7259
rect 4019 7256 4031 7259
rect 5160 7259 5218 7265
rect 4019 7228 5120 7256
rect 4019 7225 4031 7228
rect 3973 7219 4031 7225
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 2961 7191 3019 7197
rect 2961 7188 2973 7191
rect 2832 7160 2973 7188
rect 2832 7148 2838 7160
rect 2961 7157 2973 7160
rect 3007 7157 3019 7191
rect 3234 7188 3240 7200
rect 3195 7160 3240 7188
rect 2961 7151 3019 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 3510 7188 3516 7200
rect 3471 7160 3516 7188
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4062 7148 4068 7200
rect 4120 7188 4126 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 4120 7160 4537 7188
rect 4120 7148 4126 7160
rect 4525 7157 4537 7160
rect 4571 7157 4583 7191
rect 4798 7188 4804 7200
rect 4759 7160 4804 7188
rect 4525 7151 4583 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 5092 7188 5120 7228
rect 5160 7225 5172 7259
rect 5206 7256 5218 7259
rect 5810 7256 5816 7268
rect 5206 7228 5816 7256
rect 5206 7225 5218 7228
rect 5160 7219 5218 7225
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 6288 7256 6316 7284
rect 7576 7256 7604 7296
rect 8113 7293 8125 7327
rect 8159 7293 8171 7327
rect 8113 7287 8171 7293
rect 6288 7228 7604 7256
rect 7650 7216 7656 7268
rect 7708 7256 7714 7268
rect 8128 7256 8156 7287
rect 7708 7228 8156 7256
rect 8220 7256 8248 7364
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10410 7392 10416 7404
rect 10100 7364 10416 7392
rect 10100 7352 10106 7364
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 11155 7401 11183 7432
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 13446 7460 13452 7472
rect 12584 7432 13452 7460
rect 12584 7420 12590 7432
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 15010 7460 15016 7472
rect 14660 7432 15016 7460
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 11241 7395 11299 7401
rect 11241 7361 11253 7395
rect 11287 7361 11299 7395
rect 11241 7355 11299 7361
rect 12115 7395 12173 7401
rect 12115 7361 12127 7395
rect 12161 7392 12173 7395
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 12161 7364 13093 7392
rect 12161 7361 12173 7364
rect 12115 7355 12173 7361
rect 13081 7361 13093 7364
rect 13127 7392 13139 7395
rect 13906 7392 13912 7404
rect 13127 7364 13912 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 8380 7327 8438 7333
rect 8380 7293 8392 7327
rect 8426 7324 8438 7327
rect 8938 7324 8944 7336
rect 8426 7296 8944 7324
rect 8426 7293 8438 7296
rect 8380 7287 8438 7293
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 10226 7324 10232 7336
rect 10187 7296 10232 7324
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 11256 7324 11284 7355
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 14660 7401 14688 7432
rect 15010 7420 15016 7432
rect 15068 7420 15074 7472
rect 18230 7460 18236 7472
rect 18191 7432 18236 7460
rect 18230 7420 18236 7432
rect 18288 7420 18294 7472
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7392 14887 7395
rect 15102 7392 15108 7404
rect 14875 7364 15108 7392
rect 14875 7361 14887 7364
rect 14829 7355 14887 7361
rect 15102 7352 15108 7364
rect 15160 7392 15166 7404
rect 15565 7395 15623 7401
rect 15565 7392 15577 7395
rect 15160 7364 15577 7392
rect 15160 7352 15166 7364
rect 15565 7361 15577 7364
rect 15611 7361 15623 7395
rect 15565 7355 15623 7361
rect 15654 7352 15660 7404
rect 15712 7392 15718 7404
rect 16301 7395 16359 7401
rect 16301 7392 16313 7395
rect 15712 7364 16313 7392
rect 15712 7352 15718 7364
rect 16301 7361 16313 7364
rect 16347 7361 16359 7395
rect 16301 7355 16359 7361
rect 16390 7352 16396 7404
rect 16448 7392 16454 7404
rect 16448 7364 16493 7392
rect 16448 7352 16454 7364
rect 11330 7324 11336 7336
rect 11256 7296 11336 7324
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 11885 7327 11943 7333
rect 11885 7293 11897 7327
rect 11931 7324 11943 7327
rect 12802 7324 12808 7336
rect 11931 7296 12112 7324
rect 12763 7296 12808 7324
rect 11931 7293 11943 7296
rect 11885 7287 11943 7293
rect 11146 7256 11152 7268
rect 8220 7228 11152 7256
rect 7708 7216 7714 7228
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 12084 7256 12112 7296
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 13817 7327 13875 7333
rect 13817 7293 13829 7327
rect 13863 7293 13875 7327
rect 15470 7324 15476 7336
rect 15383 7296 15476 7324
rect 13817 7287 13875 7293
rect 12342 7256 12348 7268
rect 11256 7228 11560 7256
rect 12084 7228 12348 7256
rect 5626 7188 5632 7200
rect 5092 7160 5632 7188
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 8018 7188 8024 7200
rect 7979 7160 8024 7188
rect 8018 7148 8024 7160
rect 8076 7148 8082 7200
rect 9490 7188 9496 7200
rect 9451 7160 9496 7188
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 9769 7191 9827 7197
rect 9769 7157 9781 7191
rect 9815 7188 9827 7191
rect 10321 7191 10379 7197
rect 10321 7188 10333 7191
rect 9815 7160 10333 7188
rect 9815 7157 9827 7160
rect 9769 7151 9827 7157
rect 10321 7157 10333 7160
rect 10367 7188 10379 7191
rect 10410 7188 10416 7200
rect 10367 7160 10416 7188
rect 10367 7157 10379 7160
rect 10321 7151 10379 7157
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 11057 7191 11115 7197
rect 11057 7157 11069 7191
rect 11103 7188 11115 7191
rect 11256 7188 11284 7228
rect 11532 7197 11560 7228
rect 12342 7216 12348 7228
rect 12400 7216 12406 7268
rect 13722 7256 13728 7268
rect 13683 7228 13728 7256
rect 13722 7216 13728 7228
rect 13780 7216 13786 7268
rect 11103 7160 11284 7188
rect 11517 7191 11575 7197
rect 11103 7157 11115 7160
rect 11057 7151 11115 7157
rect 11517 7157 11529 7191
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 11977 7191 12035 7197
rect 11977 7157 11989 7191
rect 12023 7188 12035 7191
rect 12158 7188 12164 7200
rect 12023 7160 12164 7188
rect 12023 7157 12035 7160
rect 11977 7151 12035 7157
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12308 7160 12909 7188
rect 12308 7148 12314 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 13354 7188 13360 7200
rect 13315 7160 13360 7188
rect 12897 7151 12955 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 13630 7148 13636 7200
rect 13688 7188 13694 7200
rect 13832 7188 13860 7287
rect 15470 7284 15476 7296
rect 15528 7324 15534 7336
rect 16482 7324 16488 7336
rect 15528 7296 16488 7324
rect 15528 7284 15534 7296
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 17954 7284 17960 7336
rect 18012 7324 18018 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 18012 7296 18061 7324
rect 18012 7284 18018 7296
rect 18049 7293 18061 7296
rect 18095 7324 18107 7327
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18095 7296 18429 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 16209 7259 16267 7265
rect 16209 7256 16221 7259
rect 15028 7228 16221 7256
rect 14550 7188 14556 7200
rect 13688 7160 13860 7188
rect 14511 7160 14556 7188
rect 13688 7148 13694 7160
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 15028 7197 15056 7228
rect 16209 7225 16221 7228
rect 16255 7225 16267 7259
rect 16209 7219 16267 7225
rect 15013 7191 15071 7197
rect 15013 7157 15025 7191
rect 15059 7157 15071 7191
rect 15378 7188 15384 7200
rect 15339 7160 15384 7188
rect 15013 7151 15071 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 2041 6987 2099 6993
rect 2041 6953 2053 6987
rect 2087 6984 2099 6987
rect 2866 6984 2872 6996
rect 2087 6956 2872 6984
rect 2087 6953 2099 6956
rect 2041 6947 2099 6953
rect 2866 6944 2872 6956
rect 2924 6944 2930 6996
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 4525 6987 4583 6993
rect 4525 6984 4537 6987
rect 3660 6956 4537 6984
rect 3660 6944 3666 6956
rect 4525 6953 4537 6956
rect 4571 6984 4583 6987
rect 4614 6984 4620 6996
rect 4571 6956 4620 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 5629 6987 5687 6993
rect 5629 6984 5641 6987
rect 4856 6956 5641 6984
rect 4856 6944 4862 6956
rect 5629 6953 5641 6956
rect 5675 6984 5687 6987
rect 5902 6984 5908 6996
rect 5675 6956 5908 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6089 6987 6147 6993
rect 6089 6984 6101 6987
rect 6052 6956 6101 6984
rect 6052 6944 6058 6956
rect 6089 6953 6101 6956
rect 6135 6953 6147 6987
rect 11238 6984 11244 6996
rect 6089 6947 6147 6953
rect 6288 6956 7512 6984
rect 2130 6916 2136 6928
rect 2091 6888 2136 6916
rect 2130 6876 2136 6888
rect 2188 6876 2194 6928
rect 4338 6916 4344 6928
rect 2240 6888 4344 6916
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 2240 6848 2268 6888
rect 4338 6876 4344 6888
rect 4396 6876 4402 6928
rect 4706 6876 4712 6928
rect 4764 6916 4770 6928
rect 5721 6919 5779 6925
rect 5721 6916 5733 6919
rect 4764 6888 5733 6916
rect 4764 6876 4770 6888
rect 5721 6885 5733 6888
rect 5767 6885 5779 6919
rect 5920 6916 5948 6944
rect 6288 6916 6316 6956
rect 5920 6888 6316 6916
rect 7484 6916 7512 6956
rect 9232 6956 11244 6984
rect 9232 6916 9260 6956
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 11514 6984 11520 6996
rect 11475 6956 11520 6984
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12621 6987 12679 6993
rect 12621 6984 12633 6987
rect 12124 6956 12633 6984
rect 12124 6944 12130 6956
rect 12621 6953 12633 6956
rect 12667 6953 12679 6987
rect 12621 6947 12679 6953
rect 12713 6987 12771 6993
rect 12713 6953 12725 6987
rect 12759 6984 12771 6987
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 12759 6956 13093 6984
rect 12759 6953 12771 6956
rect 12713 6947 12771 6953
rect 13081 6953 13093 6956
rect 13127 6953 13139 6987
rect 13081 6947 13139 6953
rect 7484 6888 9260 6916
rect 5721 6879 5779 6885
rect 11146 6876 11152 6928
rect 11204 6916 11210 6928
rect 11701 6919 11759 6925
rect 11701 6916 11713 6919
rect 11204 6888 11713 6916
rect 11204 6876 11210 6888
rect 11701 6885 11713 6888
rect 11747 6916 11759 6919
rect 12158 6916 12164 6928
rect 11747 6888 12164 6916
rect 11747 6885 11759 6888
rect 11701 6879 11759 6885
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 2774 6857 2780 6860
rect 2768 6848 2780 6857
rect 1912 6820 2268 6848
rect 2332 6820 2780 6848
rect 1912 6808 1918 6820
rect 2332 6789 2360 6820
rect 2768 6811 2780 6820
rect 2832 6848 2838 6860
rect 4433 6851 4491 6857
rect 2832 6820 2916 6848
rect 2774 6808 2780 6811
rect 2832 6808 2838 6820
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 4798 6848 4804 6860
rect 4479 6820 4804 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 4798 6808 4804 6820
rect 4856 6848 4862 6860
rect 5074 6848 5080 6860
rect 4856 6820 5080 6848
rect 4856 6808 4862 6820
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6848 5227 6851
rect 5215 6820 5672 6848
rect 5215 6817 5227 6820
rect 5169 6811 5227 6817
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6749 2375 6783
rect 2317 6743 2375 6749
rect 2406 6740 2412 6792
rect 2464 6780 2470 6792
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 2464 6752 2513 6780
rect 2464 6740 2470 6752
rect 2501 6749 2513 6752
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 1762 6712 1768 6724
rect 1627 6684 1768 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 1762 6672 1768 6684
rect 1820 6672 1826 6724
rect 3881 6715 3939 6721
rect 3881 6681 3893 6715
rect 3927 6712 3939 6715
rect 4338 6712 4344 6724
rect 3927 6684 4344 6712
rect 3927 6681 3939 6684
rect 3881 6675 3939 6681
rect 4338 6672 4344 6684
rect 4396 6712 4402 6724
rect 4632 6712 4660 6743
rect 4396 6684 4660 6712
rect 5261 6715 5319 6721
rect 4396 6672 4402 6684
rect 5261 6681 5273 6715
rect 5307 6712 5319 6715
rect 5534 6712 5540 6724
rect 5307 6684 5540 6712
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 5644 6712 5672 6820
rect 6362 6808 6368 6860
rect 6420 6848 6426 6860
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 6420 6820 6469 6848
rect 6420 6808 6426 6820
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 7190 6857 7196 6860
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 6880 6820 6929 6848
rect 6880 6808 6886 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 7184 6848 7196 6857
rect 7151 6820 7196 6848
rect 6917 6811 6975 6817
rect 7184 6811 7196 6820
rect 7190 6808 7196 6811
rect 7248 6808 7254 6860
rect 9122 6848 9128 6860
rect 9083 6820 9128 6848
rect 9122 6808 9128 6820
rect 9180 6848 9186 6860
rect 9861 6851 9919 6857
rect 9861 6848 9873 6851
rect 9180 6820 9873 6848
rect 9180 6808 9186 6820
rect 9861 6817 9873 6820
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10226 6848 10232 6860
rect 10183 6820 10232 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 10404 6851 10462 6857
rect 10404 6817 10416 6851
rect 10450 6848 10462 6851
rect 11330 6848 11336 6860
rect 10450 6820 11336 6848
rect 10450 6817 10462 6820
rect 10404 6811 10462 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 12636 6848 12664 6947
rect 13262 6944 13268 6996
rect 13320 6984 13326 6996
rect 13320 6956 13492 6984
rect 13320 6944 13326 6956
rect 13464 6925 13492 6956
rect 13630 6944 13636 6996
rect 13688 6984 13694 6996
rect 13909 6987 13967 6993
rect 13909 6984 13921 6987
rect 13688 6956 13921 6984
rect 13688 6944 13694 6956
rect 13909 6953 13921 6956
rect 13955 6953 13967 6987
rect 13909 6947 13967 6953
rect 14016 6956 15056 6984
rect 13449 6919 13507 6925
rect 13449 6885 13461 6919
rect 13495 6916 13507 6919
rect 14016 6916 14044 6956
rect 13495 6888 14044 6916
rect 14277 6919 14335 6925
rect 13495 6885 13507 6888
rect 13449 6879 13507 6885
rect 14277 6885 14289 6919
rect 14323 6885 14335 6919
rect 14277 6879 14335 6885
rect 14090 6848 14096 6860
rect 12636 6820 14096 6848
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 14292 6792 14320 6879
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 15028 6916 15056 6956
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 15473 6987 15531 6993
rect 15473 6984 15485 6987
rect 15436 6956 15485 6984
rect 15436 6944 15442 6956
rect 15473 6953 15485 6956
rect 15519 6953 15531 6987
rect 15473 6947 15531 6953
rect 15841 6987 15899 6993
rect 15841 6953 15853 6987
rect 15887 6984 15899 6987
rect 16114 6984 16120 6996
rect 15887 6956 16120 6984
rect 15887 6953 15899 6956
rect 15841 6947 15899 6953
rect 15856 6916 15884 6947
rect 16114 6944 16120 6956
rect 16172 6944 16178 6996
rect 14424 6888 14688 6916
rect 15028 6888 15884 6916
rect 17589 6919 17647 6925
rect 14424 6876 14430 6888
rect 14660 6848 14688 6888
rect 17589 6885 17601 6919
rect 17635 6916 17647 6919
rect 17635 6888 18276 6916
rect 17635 6885 17647 6888
rect 17589 6879 17647 6885
rect 17604 6848 17632 6879
rect 18248 6857 18276 6888
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 14384 6820 14596 6848
rect 14660 6820 17632 6848
rect 17696 6820 17877 6848
rect 5902 6780 5908 6792
rect 5815 6752 5908 6780
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 6549 6783 6607 6789
rect 6549 6780 6561 6783
rect 6328 6752 6561 6780
rect 6328 6740 6334 6752
rect 6549 6749 6561 6752
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 9217 6783 9275 6789
rect 6779 6752 6868 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 5718 6712 5724 6724
rect 5644 6684 5724 6712
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 5920 6712 5948 6740
rect 6840 6712 6868 6752
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 10042 6780 10048 6792
rect 9447 6752 10048 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 5920 6684 6868 6712
rect 1673 6647 1731 6653
rect 1673 6613 1685 6647
rect 1719 6644 1731 6647
rect 2222 6644 2228 6656
rect 1719 6616 2228 6644
rect 1719 6613 1731 6616
rect 1673 6607 1731 6613
rect 2222 6604 2228 6616
rect 2280 6604 2286 6656
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6644 4123 6647
rect 4522 6644 4528 6656
rect 4111 6616 4528 6644
rect 4111 6613 4123 6616
rect 4065 6607 4123 6613
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 4985 6647 5043 6653
rect 4985 6613 4997 6647
rect 5031 6644 5043 6647
rect 5810 6644 5816 6656
rect 5031 6616 5816 6644
rect 5031 6613 5043 6616
rect 4985 6607 5043 6613
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 6840 6644 6868 6684
rect 7926 6672 7932 6724
rect 7984 6712 7990 6724
rect 8297 6715 8355 6721
rect 8297 6712 8309 6715
rect 7984 6684 8309 6712
rect 7984 6672 7990 6684
rect 8297 6681 8309 6684
rect 8343 6681 8355 6715
rect 8297 6675 8355 6681
rect 8665 6715 8723 6721
rect 8665 6681 8677 6715
rect 8711 6712 8723 6715
rect 9232 6712 9260 6743
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 11204 6752 12909 6780
rect 11204 6740 11210 6752
rect 12897 6749 12909 6752
rect 12943 6780 12955 6783
rect 12943 6752 13032 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 9582 6712 9588 6724
rect 8711 6684 9588 6712
rect 8711 6681 8723 6684
rect 8665 6675 8723 6681
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 11164 6684 12664 6712
rect 7944 6644 7972 6672
rect 8386 6644 8392 6656
rect 6840 6616 7972 6644
rect 8347 6616 8392 6644
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 9674 6644 9680 6656
rect 8803 6616 9680 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 11164 6644 11192 6684
rect 9815 6616 11192 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 11885 6647 11943 6653
rect 11885 6644 11897 6647
rect 11572 6616 11897 6644
rect 11572 6604 11578 6616
rect 11885 6613 11897 6616
rect 11931 6644 11943 6647
rect 12066 6644 12072 6656
rect 11931 6616 12072 6644
rect 11931 6613 11943 6616
rect 11885 6607 11943 6613
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 12253 6647 12311 6653
rect 12253 6644 12265 6647
rect 12216 6616 12265 6644
rect 12216 6604 12222 6616
rect 12253 6613 12265 6616
rect 12299 6613 12311 6647
rect 12636 6644 12664 6684
rect 12802 6644 12808 6656
rect 12636 6616 12808 6644
rect 12253 6607 12311 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 13004 6644 13032 6752
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13136 6752 13553 6780
rect 13136 6740 13142 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13740 6712 13768 6743
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 14384 6789 14412 6820
rect 14369 6783 14427 6789
rect 14369 6749 14381 6783
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 13814 6712 13820 6724
rect 13727 6684 13820 6712
rect 13814 6672 13820 6684
rect 13872 6712 13878 6724
rect 14476 6712 14504 6743
rect 13872 6684 14504 6712
rect 14568 6712 14596 6820
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 14921 6783 14979 6789
rect 14921 6780 14933 6783
rect 14700 6752 14933 6780
rect 14700 6740 14706 6752
rect 14921 6749 14933 6752
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 15068 6752 15301 6780
rect 15068 6740 15074 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 14826 6712 14832 6724
rect 14568 6684 14832 6712
rect 13872 6672 13878 6684
rect 14826 6672 14832 6684
rect 14884 6712 14890 6724
rect 16942 6712 16948 6724
rect 14884 6684 16948 6712
rect 14884 6672 14890 6684
rect 16942 6672 16948 6684
rect 17000 6672 17006 6724
rect 13906 6644 13912 6656
rect 13004 6616 13912 6644
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 14642 6644 14648 6656
rect 14332 6616 14648 6644
rect 14332 6604 14338 6616
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 17494 6604 17500 6656
rect 17552 6644 17558 6656
rect 17696 6653 17724 6820
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 18233 6851 18291 6857
rect 18233 6817 18245 6851
rect 18279 6817 18291 6851
rect 18233 6811 18291 6817
rect 18414 6712 18420 6724
rect 18375 6684 18420 6712
rect 18414 6672 18420 6684
rect 18472 6672 18478 6724
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17552 6616 17693 6644
rect 17552 6604 17558 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 18046 6644 18052 6656
rect 18007 6616 18052 6644
rect 17681 6607 17739 6613
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 2866 6440 2872 6452
rect 2823 6412 2872 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 3602 6440 3608 6452
rect 3563 6412 3608 6440
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 3712 6412 5457 6440
rect 2225 6375 2283 6381
rect 2225 6341 2237 6375
rect 2271 6372 2283 6375
rect 2958 6372 2964 6384
rect 2271 6344 2964 6372
rect 2271 6341 2283 6344
rect 2225 6335 2283 6341
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 3712 6372 3740 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 5905 6443 5963 6449
rect 5905 6409 5917 6443
rect 5951 6440 5963 6443
rect 6270 6440 6276 6452
rect 5951 6412 6276 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 7190 6440 7196 6452
rect 6564 6412 7196 6440
rect 3068 6344 3740 6372
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6304 1547 6307
rect 1535 6276 2452 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 1762 6236 1768 6248
rect 1719 6208 1768 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 2424 6245 2452 6276
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3068 6304 3096 6344
rect 3418 6304 3424 6316
rect 2832 6276 3096 6304
rect 3379 6276 3424 6304
rect 2832 6264 2838 6276
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 6365 6307 6423 6313
rect 5132 6276 6316 6304
rect 5132 6264 5138 6276
rect 2041 6239 2099 6245
rect 2041 6236 2053 6239
rect 2004 6208 2053 6236
rect 2004 6196 2010 6208
rect 2041 6205 2053 6208
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2498 6236 2504 6248
rect 2455 6208 2504 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3510 6236 3516 6248
rect 3191 6208 3516 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 4056 6239 4114 6245
rect 4056 6205 4068 6239
rect 4102 6236 4114 6239
rect 4338 6236 4344 6248
rect 4102 6208 4344 6236
rect 4102 6205 4114 6208
rect 4056 6199 4114 6205
rect 3237 6171 3295 6177
rect 3237 6137 3249 6171
rect 3283 6168 3295 6171
rect 3326 6168 3332 6180
rect 3283 6140 3332 6168
rect 3283 6137 3295 6140
rect 3237 6131 3295 6137
rect 3326 6128 3332 6140
rect 3384 6128 3390 6180
rect 3418 6128 3424 6180
rect 3476 6168 3482 6180
rect 3804 6168 3832 6199
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 5626 6236 5632 6248
rect 5307 6208 5632 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5626 6196 5632 6208
rect 5684 6236 5690 6248
rect 5813 6239 5871 6245
rect 5684 6208 5764 6236
rect 5684 6196 5690 6208
rect 4890 6168 4896 6180
rect 3476 6140 3832 6168
rect 3476 6128 3482 6140
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1452 6072 1869 6100
rect 1452 6060 1458 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 1857 6063 1915 6069
rect 2593 6103 2651 6109
rect 2593 6069 2605 6103
rect 2639 6100 2651 6103
rect 2774 6100 2780 6112
rect 2639 6072 2780 6100
rect 2639 6069 2651 6072
rect 2593 6063 2651 6069
rect 2774 6060 2780 6072
rect 2832 6060 2838 6112
rect 3804 6100 3832 6140
rect 4540 6140 4896 6168
rect 4540 6100 4568 6140
rect 4890 6128 4896 6140
rect 4948 6168 4954 6180
rect 5736 6168 5764 6208
rect 5813 6205 5825 6239
rect 5859 6236 5871 6239
rect 5902 6236 5908 6248
rect 5859 6208 5908 6236
rect 5859 6205 5871 6208
rect 5813 6199 5871 6205
rect 5902 6196 5908 6208
rect 5960 6196 5966 6248
rect 6288 6245 6316 6276
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 6454 6304 6460 6316
rect 6411 6276 6460 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 6564 6313 6592 6412
rect 7190 6400 7196 6412
rect 7248 6440 7254 6452
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 7248 6412 8217 6440
rect 7248 6400 7254 6412
rect 8205 6409 8217 6412
rect 8251 6409 8263 6443
rect 8205 6403 8263 6409
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 10229 6443 10287 6449
rect 10229 6440 10241 6443
rect 9180 6412 10241 6440
rect 9180 6400 9186 6412
rect 10229 6409 10241 6412
rect 10275 6409 10287 6443
rect 10502 6440 10508 6452
rect 10463 6412 10508 6440
rect 10229 6403 10287 6409
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 11514 6440 11520 6452
rect 10888 6412 11520 6440
rect 9950 6332 9956 6384
rect 10008 6372 10014 6384
rect 10888 6372 10916 6412
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12805 6443 12863 6449
rect 12805 6440 12817 6443
rect 12492 6412 12817 6440
rect 12492 6400 12498 6412
rect 12805 6409 12817 6412
rect 12851 6440 12863 6443
rect 13078 6440 13084 6452
rect 12851 6412 13084 6440
rect 12851 6409 12863 6412
rect 12805 6403 12863 6409
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13722 6440 13728 6452
rect 13219 6412 13728 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 15381 6443 15439 6449
rect 15381 6440 15393 6443
rect 13964 6412 15393 6440
rect 13964 6400 13970 6412
rect 15381 6409 15393 6412
rect 15427 6409 15439 6443
rect 15381 6403 15439 6409
rect 10008 6344 10916 6372
rect 10008 6332 10014 6344
rect 15010 6332 15016 6384
rect 15068 6372 15074 6384
rect 15473 6375 15531 6381
rect 15473 6372 15485 6375
rect 15068 6344 15485 6372
rect 15068 6332 15074 6344
rect 15473 6341 15485 6344
rect 15519 6341 15531 6375
rect 15473 6335 15531 6341
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6822 6304 6828 6316
rect 6696 6276 6828 6304
rect 6696 6264 6702 6276
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 10042 6304 10048 6316
rect 9784 6276 10048 6304
rect 6273 6239 6331 6245
rect 6273 6205 6285 6239
rect 6319 6236 6331 6239
rect 6730 6236 6736 6248
rect 6319 6208 6736 6236
rect 6319 6205 6331 6208
rect 6273 6199 6331 6205
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 7092 6239 7150 6245
rect 7092 6205 7104 6239
rect 7138 6236 7150 6239
rect 7466 6236 7472 6248
rect 7138 6208 7472 6236
rect 7138 6205 7150 6208
rect 7092 6199 7150 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 7708 6208 8769 6236
rect 7708 6196 7714 6208
rect 8757 6205 8769 6208
rect 8803 6205 8815 6239
rect 9784 6236 9812 6276
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 13814 6304 13820 6316
rect 13775 6276 13820 6304
rect 13814 6264 13820 6276
rect 13872 6304 13878 6316
rect 13872 6276 14136 6304
rect 13872 6264 13878 6276
rect 8757 6199 8815 6205
rect 8864 6208 9812 6236
rect 4948 6140 5672 6168
rect 5736 6140 6776 6168
rect 4948 6128 4954 6140
rect 3804 6072 4568 6100
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 5644 6109 5672 6140
rect 5828 6112 5856 6140
rect 6748 6112 6776 6140
rect 6914 6128 6920 6180
rect 6972 6168 6978 6180
rect 8389 6171 8447 6177
rect 8389 6168 8401 6171
rect 6972 6140 8401 6168
rect 6972 6128 6978 6140
rect 8389 6137 8401 6140
rect 8435 6168 8447 6171
rect 8864 6168 8892 6208
rect 9858 6196 9864 6248
rect 9916 6236 9922 6248
rect 10226 6236 10232 6248
rect 9916 6208 10232 6236
rect 9916 6196 9922 6208
rect 10226 6196 10232 6208
rect 10284 6236 10290 6248
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10284 6208 10885 6236
rect 10284 6196 10290 6208
rect 10873 6205 10885 6208
rect 10919 6236 10931 6239
rect 10962 6236 10968 6248
rect 10919 6208 10968 6236
rect 10919 6205 10931 6208
rect 10873 6199 10931 6205
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 11146 6245 11152 6248
rect 11140 6236 11152 6245
rect 11107 6208 11152 6236
rect 11140 6199 11152 6208
rect 11146 6196 11152 6199
rect 11204 6196 11210 6248
rect 12618 6236 12624 6248
rect 12579 6208 12624 6236
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 13446 6196 13452 6248
rect 13504 6236 13510 6248
rect 13722 6236 13728 6248
rect 13504 6208 13728 6236
rect 13504 6196 13510 6208
rect 13722 6196 13728 6208
rect 13780 6236 13786 6248
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13780 6208 14013 6236
rect 13780 6196 13786 6208
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14108 6236 14136 6276
rect 14257 6239 14315 6245
rect 14257 6236 14269 6239
rect 14108 6208 14269 6236
rect 14001 6199 14059 6205
rect 14257 6205 14269 6208
rect 14303 6205 14315 6239
rect 14257 6199 14315 6205
rect 17954 6196 17960 6248
rect 18012 6236 18018 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 18012 6208 18061 6236
rect 18012 6196 18018 6208
rect 18049 6205 18061 6208
rect 18095 6236 18107 6239
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 18095 6208 18429 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 8435 6140 8892 6168
rect 9024 6171 9082 6177
rect 8435 6137 8447 6140
rect 8389 6131 8447 6137
rect 9024 6137 9036 6171
rect 9070 6168 9082 6171
rect 9490 6168 9496 6180
rect 9070 6140 9496 6168
rect 9070 6137 9082 6140
rect 9024 6131 9082 6137
rect 9490 6128 9496 6140
rect 9548 6128 9554 6180
rect 10594 6168 10600 6180
rect 9600 6140 10600 6168
rect 5169 6103 5227 6109
rect 5169 6100 5181 6103
rect 4672 6072 5181 6100
rect 4672 6060 4678 6072
rect 5169 6069 5181 6072
rect 5215 6069 5227 6103
rect 5169 6063 5227 6069
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6069 5687 6103
rect 5629 6063 5687 6069
rect 5810 6060 5816 6112
rect 5868 6060 5874 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 8018 6100 8024 6112
rect 6788 6072 8024 6100
rect 6788 6060 6794 6072
rect 8018 6060 8024 6072
rect 8076 6100 8082 6112
rect 8573 6103 8631 6109
rect 8573 6100 8585 6103
rect 8076 6072 8585 6100
rect 8076 6060 8082 6072
rect 8573 6069 8585 6072
rect 8619 6100 8631 6103
rect 9600 6100 9628 6140
rect 10594 6128 10600 6140
rect 10652 6128 10658 6180
rect 11054 6128 11060 6180
rect 11112 6168 11118 6180
rect 11974 6168 11980 6180
rect 11112 6140 11980 6168
rect 11112 6128 11118 6140
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 12066 6128 12072 6180
rect 12124 6168 12130 6180
rect 12124 6140 12480 6168
rect 12124 6128 12130 6140
rect 10134 6100 10140 6112
rect 8619 6072 9628 6100
rect 10095 6072 10140 6100
rect 8619 6069 8631 6072
rect 8573 6063 8631 6069
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10689 6103 10747 6109
rect 10689 6100 10701 6103
rect 10284 6072 10701 6100
rect 10284 6060 10290 6072
rect 10689 6069 10701 6072
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 12253 6103 12311 6109
rect 12253 6100 12265 6103
rect 11388 6072 12265 6100
rect 11388 6060 11394 6072
rect 12253 6069 12265 6072
rect 12299 6100 12311 6103
rect 12342 6100 12348 6112
rect 12299 6072 12348 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 12452 6109 12480 6140
rect 12802 6128 12808 6180
rect 12860 6168 12866 6180
rect 13541 6171 13599 6177
rect 13541 6168 13553 6171
rect 12860 6140 13553 6168
rect 12860 6128 12866 6140
rect 13541 6137 13553 6140
rect 13587 6168 13599 6171
rect 14366 6168 14372 6180
rect 13587 6140 14372 6168
rect 13587 6137 13599 6140
rect 13541 6131 13599 6137
rect 14366 6128 14372 6140
rect 14424 6168 14430 6180
rect 15010 6168 15016 6180
rect 14424 6140 15016 6168
rect 14424 6128 14430 6140
rect 15010 6128 15016 6140
rect 15068 6128 15074 6180
rect 12437 6103 12495 6109
rect 12437 6069 12449 6103
rect 12483 6069 12495 6103
rect 12437 6063 12495 6069
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 13081 6103 13139 6109
rect 13081 6100 13093 6103
rect 12676 6072 13093 6100
rect 12676 6060 12682 6072
rect 13081 6069 13093 6072
rect 13127 6100 13139 6103
rect 13633 6103 13691 6109
rect 13633 6100 13645 6103
rect 13127 6072 13645 6100
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 13633 6069 13645 6072
rect 13679 6100 13691 6103
rect 14458 6100 14464 6112
rect 13679 6072 14464 6100
rect 13679 6069 13691 6072
rect 13633 6063 13691 6069
rect 14458 6060 14464 6072
rect 14516 6100 14522 6112
rect 17218 6100 17224 6112
rect 14516 6072 17224 6100
rect 14516 6060 14522 6072
rect 17218 6060 17224 6072
rect 17276 6060 17282 6112
rect 18230 6100 18236 6112
rect 18191 6072 18236 6100
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 2406 5896 2412 5908
rect 1596 5868 2412 5896
rect 1596 5772 1624 5868
rect 2406 5856 2412 5868
rect 2464 5896 2470 5908
rect 3418 5896 3424 5908
rect 2464 5868 3424 5896
rect 2464 5856 2470 5868
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3651 5868 4077 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4522 5896 4528 5908
rect 4483 5868 4528 5896
rect 4065 5859 4123 5865
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 6638 5896 6644 5908
rect 5368 5868 6644 5896
rect 1756 5831 1814 5837
rect 1756 5797 1768 5831
rect 1802 5828 1814 5831
rect 1802 5800 4568 5828
rect 1802 5797 1814 5800
rect 1756 5791 1814 5797
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5760 1547 5763
rect 1578 5760 1584 5772
rect 1535 5732 1584 5760
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 1578 5720 1584 5732
rect 1636 5720 1642 5772
rect 3510 5760 3516 5772
rect 3471 5732 3516 5760
rect 3510 5720 3516 5732
rect 3568 5720 3574 5772
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 3697 5695 3755 5701
rect 3697 5692 3709 5695
rect 2884 5664 3709 5692
rect 2884 5568 2912 5664
rect 3697 5661 3709 5664
rect 3743 5661 3755 5695
rect 3697 5655 3755 5661
rect 2961 5627 3019 5633
rect 2961 5593 2973 5627
rect 3007 5624 3019 5627
rect 4448 5624 4476 5723
rect 4540 5692 4568 5800
rect 5368 5769 5396 5868
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 9309 5899 9367 5905
rect 9309 5865 9321 5899
rect 9355 5896 9367 5899
rect 9858 5896 9864 5908
rect 9355 5868 9864 5896
rect 9355 5865 9367 5868
rect 9309 5859 9367 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 11146 5896 11152 5908
rect 10100 5868 11152 5896
rect 10100 5856 10106 5868
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 11333 5899 11391 5905
rect 11333 5896 11345 5899
rect 11296 5868 11345 5896
rect 11296 5856 11302 5868
rect 11333 5865 11345 5868
rect 11379 5865 11391 5899
rect 11333 5859 11391 5865
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 11793 5899 11851 5905
rect 11793 5896 11805 5899
rect 11664 5868 11805 5896
rect 11664 5856 11670 5868
rect 11793 5865 11805 5868
rect 11839 5865 11851 5899
rect 12158 5896 12164 5908
rect 12119 5868 12164 5896
rect 11793 5859 11851 5865
rect 12158 5856 12164 5868
rect 12216 5856 12222 5908
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 13354 5896 13360 5908
rect 12299 5868 13360 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 14001 5899 14059 5905
rect 14001 5896 14013 5899
rect 13872 5868 14013 5896
rect 13872 5856 13878 5868
rect 14001 5865 14013 5868
rect 14047 5865 14059 5899
rect 14001 5859 14059 5865
rect 14090 5856 14096 5908
rect 14148 5896 14154 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 14148 5868 17693 5896
rect 14148 5856 14154 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 7098 5828 7104 5840
rect 5460 5800 7104 5828
rect 4893 5763 4951 5769
rect 4893 5729 4905 5763
rect 4939 5729 4951 5763
rect 4893 5723 4951 5729
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5729 5411 5763
rect 5353 5723 5411 5729
rect 4614 5692 4620 5704
rect 4527 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4908 5692 4936 5723
rect 5460 5692 5488 5800
rect 7098 5788 7104 5800
rect 7156 5788 7162 5840
rect 7193 5831 7251 5837
rect 7193 5797 7205 5831
rect 7239 5828 7251 5831
rect 9214 5828 9220 5840
rect 7239 5800 9220 5828
rect 7239 5797 7251 5800
rect 7193 5791 7251 5797
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 12066 5828 12072 5840
rect 9508 5800 12072 5828
rect 5626 5769 5632 5772
rect 5620 5723 5632 5769
rect 5684 5760 5690 5772
rect 5684 5732 5720 5760
rect 5626 5720 5632 5723
rect 5684 5720 5690 5732
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 9508 5769 9536 5800
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 12636 5800 13032 5828
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 5960 5732 7849 5760
rect 5960 5720 5966 5732
rect 7837 5729 7849 5732
rect 7883 5729 7895 5763
rect 7837 5723 7895 5729
rect 8573 5763 8631 5769
rect 8573 5729 8585 5763
rect 8619 5760 8631 5763
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8619 5732 9045 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 9033 5729 9045 5732
rect 9079 5729 9091 5763
rect 9033 5723 9091 5729
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5729 9551 5763
rect 9858 5760 9864 5772
rect 9819 5732 9864 5760
rect 9493 5723 9551 5729
rect 9858 5720 9864 5732
rect 9916 5720 9922 5772
rect 10134 5769 10140 5772
rect 10128 5760 10140 5769
rect 10047 5732 10140 5760
rect 10128 5723 10140 5732
rect 10192 5760 10198 5772
rect 11514 5760 11520 5772
rect 10192 5732 11520 5760
rect 10134 5720 10140 5723
rect 10192 5720 10198 5732
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12636 5769 12664 5800
rect 12621 5763 12679 5769
rect 12621 5760 12633 5763
rect 12492 5732 12633 5760
rect 12492 5720 12498 5732
rect 12621 5729 12633 5732
rect 12667 5729 12679 5763
rect 12621 5723 12679 5729
rect 12710 5720 12716 5772
rect 12768 5760 12774 5772
rect 12877 5763 12935 5769
rect 12877 5760 12889 5763
rect 12768 5732 12889 5760
rect 12768 5720 12774 5732
rect 12877 5729 12889 5732
rect 12923 5729 12935 5763
rect 13004 5760 13032 5800
rect 13630 5760 13636 5772
rect 13004 5732 13636 5760
rect 12877 5723 12935 5729
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 13906 5720 13912 5772
rect 13964 5760 13970 5772
rect 14461 5763 14519 5769
rect 14461 5760 14473 5763
rect 13964 5732 14473 5760
rect 13964 5720 13970 5732
rect 14461 5729 14473 5732
rect 14507 5760 14519 5763
rect 14921 5763 14979 5769
rect 14921 5760 14933 5763
rect 14507 5732 14933 5760
rect 14507 5729 14519 5732
rect 14461 5723 14519 5729
rect 14921 5729 14933 5732
rect 14967 5760 14979 5763
rect 17494 5760 17500 5772
rect 14967 5732 17500 5760
rect 14967 5729 14979 5732
rect 14921 5723 14979 5729
rect 17494 5720 17500 5732
rect 17552 5720 17558 5772
rect 17696 5760 17724 5859
rect 17865 5763 17923 5769
rect 17865 5760 17877 5763
rect 17696 5732 17877 5760
rect 17865 5729 17877 5732
rect 17911 5729 17923 5763
rect 18230 5760 18236 5772
rect 18191 5732 18236 5760
rect 17865 5723 17923 5729
rect 18230 5720 18236 5732
rect 18288 5720 18294 5772
rect 7282 5692 7288 5704
rect 4908 5664 5488 5692
rect 7243 5664 7288 5692
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5692 7435 5695
rect 7466 5692 7472 5704
rect 7423 5664 7472 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 5350 5624 5356 5636
rect 3007 5596 5356 5624
rect 3007 5593 3019 5596
rect 2961 5587 3019 5593
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 6733 5627 6791 5633
rect 6733 5593 6745 5627
rect 6779 5624 6791 5627
rect 7392 5624 7420 5655
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 8665 5695 8723 5701
rect 8665 5692 8677 5695
rect 8536 5664 8677 5692
rect 8536 5652 8542 5664
rect 8665 5661 8677 5664
rect 8711 5661 8723 5695
rect 8665 5655 8723 5661
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 8812 5664 8857 5692
rect 8812 5652 8818 5664
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 11330 5692 11336 5704
rect 10928 5664 11336 5692
rect 10928 5652 10934 5664
rect 11330 5652 11336 5664
rect 11388 5692 11394 5704
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11388 5664 11621 5692
rect 11388 5652 11394 5664
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 12342 5692 12348 5704
rect 12303 5664 12348 5692
rect 11609 5655 11667 5661
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 14550 5692 14556 5704
rect 14511 5664 14556 5692
rect 14550 5652 14556 5664
rect 14608 5652 14614 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 15010 5692 15016 5704
rect 14783 5664 15016 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 7929 5627 7987 5633
rect 7929 5624 7941 5627
rect 6779 5596 7420 5624
rect 7484 5596 7941 5624
rect 6779 5593 6791 5596
rect 6733 5587 6791 5593
rect 2866 5556 2872 5568
rect 2827 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 3050 5516 3056 5568
rect 3108 5556 3114 5568
rect 3145 5559 3203 5565
rect 3145 5556 3157 5559
rect 3108 5528 3157 5556
rect 3108 5516 3114 5528
rect 3145 5525 3157 5528
rect 3191 5525 3203 5559
rect 3145 5519 3203 5525
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 3752 5528 5089 5556
rect 3752 5516 3758 5528
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5077 5519 5135 5525
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 6825 5559 6883 5565
rect 6825 5556 6837 5559
rect 5592 5528 6837 5556
rect 5592 5516 5598 5528
rect 6825 5525 6837 5528
rect 6871 5525 6883 5559
rect 6825 5519 6883 5525
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7484 5556 7512 5596
rect 7929 5593 7941 5596
rect 7975 5624 7987 5627
rect 9858 5624 9864 5636
rect 7975 5596 9864 5624
rect 7975 5593 7987 5596
rect 7929 5587 7987 5593
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 11146 5584 11152 5636
rect 11204 5624 11210 5636
rect 14274 5624 14280 5636
rect 11204 5596 12204 5624
rect 11204 5584 11210 5596
rect 12176 5568 12204 5596
rect 13547 5596 14280 5624
rect 7650 5556 7656 5568
rect 7156 5528 7512 5556
rect 7611 5528 7656 5556
rect 7156 5516 7162 5528
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 8205 5559 8263 5565
rect 8205 5525 8217 5559
rect 8251 5556 8263 5559
rect 8846 5556 8852 5568
rect 8251 5528 8852 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 8846 5516 8852 5528
rect 8904 5516 8910 5568
rect 9769 5559 9827 5565
rect 9769 5525 9781 5559
rect 9815 5556 9827 5559
rect 11054 5556 11060 5568
rect 9815 5528 11060 5556
rect 9815 5525 9827 5528
rect 9769 5519 9827 5525
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 11238 5556 11244 5568
rect 11199 5528 11244 5556
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 13547 5556 13575 5596
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 14568 5624 14596 5652
rect 15289 5627 15347 5633
rect 15289 5624 15301 5627
rect 14568 5596 15301 5624
rect 15289 5593 15301 5596
rect 15335 5593 15347 5627
rect 18414 5624 18420 5636
rect 18375 5596 18420 5624
rect 15289 5587 15347 5593
rect 18414 5584 18420 5596
rect 18472 5584 18478 5636
rect 12216 5528 13575 5556
rect 12216 5516 12222 5528
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 13872 5528 14105 5556
rect 13872 5516 13878 5528
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 14093 5519 14151 5525
rect 17862 5516 17868 5568
rect 17920 5556 17926 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 17920 5528 18061 5556
rect 17920 5516 17926 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3234 5352 3240 5364
rect 3099 5324 3240 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 3973 5355 4031 5361
rect 3973 5352 3985 5355
rect 3568 5324 3985 5352
rect 3568 5312 3574 5324
rect 3973 5321 3985 5324
rect 4019 5321 4031 5355
rect 3973 5315 4031 5321
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 7282 5352 7288 5364
rect 5951 5324 7288 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 9214 5352 9220 5364
rect 8312 5324 9067 5352
rect 9175 5324 9220 5352
rect 8312 5293 8340 5324
rect 4801 5287 4859 5293
rect 4801 5284 4813 5287
rect 3620 5256 4813 5284
rect 3620 5225 3648 5256
rect 4801 5253 4813 5256
rect 4847 5253 4859 5287
rect 4801 5247 4859 5253
rect 8297 5287 8355 5293
rect 8297 5253 8309 5287
rect 8343 5253 8355 5287
rect 8297 5247 8355 5253
rect 8389 5287 8447 5293
rect 8389 5253 8401 5287
rect 8435 5284 8447 5287
rect 8435 5256 8524 5284
rect 8435 5253 8447 5256
rect 8389 5247 8447 5253
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5185 3755 5219
rect 4614 5216 4620 5228
rect 4575 5188 4620 5216
rect 3697 5179 3755 5185
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5148 1547 5151
rect 1578 5148 1584 5160
rect 1535 5120 1584 5148
rect 1535 5117 1547 5120
rect 1489 5111 1547 5117
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 1756 5151 1814 5157
rect 1756 5117 1768 5151
rect 1802 5148 1814 5151
rect 2866 5148 2872 5160
rect 1802 5120 2872 5148
rect 1802 5117 1814 5120
rect 1756 5111 1814 5117
rect 2866 5108 2872 5120
rect 2924 5148 2930 5160
rect 3712 5148 3740 5179
rect 4614 5176 4620 5188
rect 4672 5216 4678 5228
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 4672 5188 5365 5216
rect 4672 5176 4678 5188
rect 5353 5185 5365 5188
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 5684 5188 6469 5216
rect 5684 5176 5690 5188
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 5166 5148 5172 5160
rect 2924 5120 3740 5148
rect 5127 5120 5172 5148
rect 2924 5108 2930 5120
rect 5166 5108 5172 5120
rect 5224 5108 5230 5160
rect 6472 5080 6500 5179
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 8312 5148 8340 5247
rect 6972 5120 7017 5148
rect 7116 5120 8340 5148
rect 6972 5108 6978 5120
rect 7116 5080 7144 5120
rect 6472 5052 7144 5080
rect 7184 5083 7242 5089
rect 7184 5049 7196 5083
rect 7230 5049 7242 5083
rect 8496 5080 8524 5256
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8812 5188 8953 5216
rect 8812 5176 8818 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 9039 5216 9067 5324
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 10594 5352 10600 5364
rect 9456 5324 10600 5352
rect 9456 5312 9462 5324
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10836 5324 10885 5352
rect 10836 5312 10842 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 12768 5324 13829 5352
rect 12768 5312 12774 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 13817 5315 13875 5321
rect 14016 5324 18061 5352
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 9732 5256 10548 5284
rect 9732 5244 9738 5256
rect 10520 5225 10548 5256
rect 13538 5244 13544 5296
rect 13596 5284 13602 5296
rect 14016 5284 14044 5324
rect 18049 5321 18061 5324
rect 18095 5352 18107 5355
rect 18230 5352 18236 5364
rect 18095 5324 18236 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 13596 5256 14044 5284
rect 13596 5244 13602 5256
rect 9769 5219 9827 5225
rect 9769 5216 9781 5219
rect 9039 5188 9781 5216
rect 8941 5179 8999 5185
rect 9769 5185 9781 5188
rect 9815 5185 9827 5219
rect 9769 5179 9827 5185
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5185 10563 5219
rect 10686 5216 10692 5228
rect 10647 5188 10692 5216
rect 10505 5179 10563 5185
rect 10686 5176 10692 5188
rect 10744 5216 10750 5228
rect 11425 5219 11483 5225
rect 11425 5216 11437 5219
rect 10744 5188 11437 5216
rect 10744 5176 10750 5188
rect 11425 5185 11437 5188
rect 11471 5185 11483 5219
rect 11425 5179 11483 5185
rect 11593 5188 12572 5216
rect 8846 5108 8852 5160
rect 8904 5148 8910 5160
rect 9585 5151 9643 5157
rect 9585 5148 9597 5151
rect 8904 5120 9597 5148
rect 8904 5108 8910 5120
rect 9585 5117 9597 5120
rect 9631 5117 9643 5151
rect 9585 5111 9643 5117
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5148 10471 5151
rect 11054 5148 11060 5160
rect 10459 5120 11060 5148
rect 10459 5117 10471 5120
rect 10413 5111 10471 5117
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 11330 5148 11336 5160
rect 11291 5120 11336 5148
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 9677 5083 9735 5089
rect 9677 5080 9689 5083
rect 8496 5052 9689 5080
rect 7184 5043 7242 5049
rect 9677 5049 9689 5052
rect 9723 5049 9735 5083
rect 11241 5083 11299 5089
rect 9677 5043 9735 5049
rect 9784 5052 11192 5080
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2869 5015 2927 5021
rect 2869 5012 2881 5015
rect 2372 4984 2881 5012
rect 2372 4972 2378 4984
rect 2869 4981 2881 4984
rect 2915 4981 2927 5015
rect 3142 5012 3148 5024
rect 3103 4984 3148 5012
rect 2869 4975 2927 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 3510 5012 3516 5024
rect 3471 4984 3516 5012
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 3602 4972 3608 5024
rect 3660 5012 3666 5024
rect 4341 5015 4399 5021
rect 4341 5012 4353 5015
rect 3660 4984 4353 5012
rect 3660 4972 3666 4984
rect 4341 4981 4353 4984
rect 4387 4981 4399 5015
rect 4341 4975 4399 4981
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 5261 5015 5319 5021
rect 4488 4984 4533 5012
rect 4488 4972 4494 4984
rect 5261 4981 5273 5015
rect 5307 5012 5319 5015
rect 5442 5012 5448 5024
rect 5307 4984 5448 5012
rect 5307 4981 5319 4984
rect 5261 4975 5319 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 5626 5012 5632 5024
rect 5587 4984 5632 5012
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 7199 5012 7227 5043
rect 7374 5012 7380 5024
rect 6420 4984 6465 5012
rect 7199 4984 7380 5012
rect 6420 4972 6426 4984
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 8662 4972 8668 5024
rect 8720 5012 8726 5024
rect 8757 5015 8815 5021
rect 8757 5012 8769 5015
rect 8720 4984 8769 5012
rect 8720 4972 8726 4984
rect 8757 4981 8769 4984
rect 8803 4981 8815 5015
rect 8757 4975 8815 4981
rect 8849 5015 8907 5021
rect 8849 4981 8861 5015
rect 8895 5012 8907 5015
rect 9122 5012 9128 5024
rect 8895 4984 9128 5012
rect 8895 4981 8907 4984
rect 8849 4975 8907 4981
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9214 4972 9220 5024
rect 9272 5012 9278 5024
rect 9784 5012 9812 5052
rect 9272 4984 9812 5012
rect 9272 4972 9278 4984
rect 9858 4972 9864 5024
rect 9916 5012 9922 5024
rect 10045 5015 10103 5021
rect 10045 5012 10057 5015
rect 9916 4984 10057 5012
rect 9916 4972 9922 4984
rect 10045 4981 10057 4984
rect 10091 4981 10103 5015
rect 11164 5012 11192 5052
rect 11241 5049 11253 5083
rect 11287 5080 11299 5083
rect 11422 5080 11428 5092
rect 11287 5052 11428 5080
rect 11287 5049 11299 5052
rect 11241 5043 11299 5049
rect 11422 5040 11428 5052
rect 11480 5040 11486 5092
rect 11593 5012 11621 5188
rect 12066 5108 12072 5160
rect 12124 5148 12130 5160
rect 12253 5151 12311 5157
rect 12253 5148 12265 5151
rect 12124 5120 12265 5148
rect 12124 5108 12130 5120
rect 12253 5117 12265 5120
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12544 5148 12572 5188
rect 13630 5176 13636 5228
rect 13688 5216 13694 5228
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13688 5188 14013 5216
rect 13688 5176 13694 5188
rect 14001 5185 14013 5188
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 15010 5176 15016 5228
rect 15068 5216 15074 5228
rect 16025 5219 16083 5225
rect 16025 5216 16037 5219
rect 15068 5188 16037 5216
rect 15068 5176 15074 5188
rect 16025 5185 16037 5188
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 13906 5148 13912 5160
rect 12544 5120 13912 5148
rect 12437 5111 12495 5117
rect 12452 5024 12480 5111
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 14274 5157 14280 5160
rect 14268 5148 14280 5157
rect 14187 5120 14280 5148
rect 14268 5111 14280 5120
rect 14332 5148 14338 5160
rect 15028 5148 15056 5176
rect 15930 5148 15936 5160
rect 14332 5120 15056 5148
rect 15891 5120 15936 5148
rect 14274 5108 14280 5111
rect 14332 5108 14338 5120
rect 15930 5108 15936 5120
rect 15988 5148 15994 5160
rect 16206 5148 16212 5160
rect 15988 5120 16212 5148
rect 15988 5108 15994 5120
rect 16206 5108 16212 5120
rect 16264 5148 16270 5160
rect 16301 5151 16359 5157
rect 16301 5148 16313 5151
rect 16264 5120 16313 5148
rect 16264 5108 16270 5120
rect 16301 5117 16313 5120
rect 16347 5117 16359 5151
rect 16301 5111 16359 5117
rect 12704 5083 12762 5089
rect 12704 5049 12716 5083
rect 12750 5080 12762 5083
rect 12750 5052 13584 5080
rect 12750 5049 12762 5052
rect 12704 5043 12762 5049
rect 13556 5024 13584 5052
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 13688 5052 15516 5080
rect 13688 5040 13694 5052
rect 11698 5012 11704 5024
rect 11164 4984 11621 5012
rect 11659 4984 11704 5012
rect 10045 4975 10103 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12069 5015 12127 5021
rect 12069 4981 12081 5015
rect 12115 5012 12127 5015
rect 12434 5012 12440 5024
rect 12115 4984 12440 5012
rect 12115 4981 12127 4984
rect 12069 4975 12127 4981
rect 12434 4972 12440 4984
rect 12492 5012 12498 5024
rect 13262 5012 13268 5024
rect 12492 4984 13268 5012
rect 12492 4972 12498 4984
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 15488 5021 15516 5052
rect 15381 5015 15439 5021
rect 15381 5012 15393 5015
rect 13596 4984 15393 5012
rect 13596 4972 13602 4984
rect 15381 4981 15393 4984
rect 15427 4981 15439 5015
rect 15381 4975 15439 4981
rect 15473 5015 15531 5021
rect 15473 4981 15485 5015
rect 15519 4981 15531 5015
rect 15838 5012 15844 5024
rect 15799 4984 15844 5012
rect 15473 4975 15531 4981
rect 15838 4972 15844 4984
rect 15896 4972 15902 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 1854 4808 1860 4820
rect 1627 4780 1860 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 3142 4808 3148 4820
rect 2087 4780 3148 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 4065 4811 4123 4817
rect 4065 4808 4077 4811
rect 3568 4780 4077 4808
rect 3568 4768 3574 4780
rect 4065 4777 4077 4780
rect 4111 4777 4123 4811
rect 4522 4808 4528 4820
rect 4483 4780 4528 4808
rect 4065 4771 4123 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 5077 4811 5135 4817
rect 5077 4777 5089 4811
rect 5123 4808 5135 4811
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 5123 4780 6285 4808
rect 5123 4777 5135 4780
rect 5077 4771 5135 4777
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 6730 4808 6736 4820
rect 6691 4780 6736 4808
rect 6273 4771 6331 4777
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4808 7435 4811
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 7423 4780 8677 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 8665 4777 8677 4780
rect 8711 4777 8723 4811
rect 8665 4771 8723 4777
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 10318 4808 10324 4820
rect 8904 4780 10324 4808
rect 8904 4768 8910 4780
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 11517 4811 11575 4817
rect 11517 4777 11529 4811
rect 11563 4808 11575 4811
rect 11606 4808 11612 4820
rect 11563 4780 11612 4808
rect 11563 4777 11575 4780
rect 11517 4771 11575 4777
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 12529 4811 12587 4817
rect 12529 4777 12541 4811
rect 12575 4808 12587 4811
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 12575 4780 12909 4808
rect 12575 4777 12587 4780
rect 12529 4771 12587 4777
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 12897 4771 12955 4777
rect 13265 4811 13323 4817
rect 13265 4777 13277 4811
rect 13311 4808 13323 4811
rect 13725 4811 13783 4817
rect 13725 4808 13737 4811
rect 13311 4780 13737 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 13725 4777 13737 4780
rect 13771 4777 13783 4811
rect 13725 4771 13783 4777
rect 13998 4768 14004 4820
rect 14056 4808 14062 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 14056 4780 14105 4808
rect 14056 4768 14062 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14093 4771 14151 4777
rect 14553 4811 14611 4817
rect 14553 4777 14565 4811
rect 14599 4808 14611 4811
rect 15838 4808 15844 4820
rect 14599 4780 15844 4808
rect 14599 4777 14611 4780
rect 14553 4771 14611 4777
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 2133 4743 2191 4749
rect 2133 4709 2145 4743
rect 2179 4740 2191 4743
rect 3050 4740 3056 4752
rect 2179 4712 3056 4740
rect 2179 4709 2191 4712
rect 2133 4703 2191 4709
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 4433 4743 4491 4749
rect 4433 4709 4445 4743
rect 4479 4740 4491 4743
rect 5626 4740 5632 4752
rect 4479 4712 5632 4740
rect 4479 4709 4491 4712
rect 4433 4703 4491 4709
rect 5626 4700 5632 4712
rect 5684 4700 5690 4752
rect 7285 4743 7343 4749
rect 7285 4709 7297 4743
rect 7331 4740 7343 4743
rect 7558 4740 7564 4752
rect 7331 4712 7564 4740
rect 7331 4709 7343 4712
rect 7285 4703 7343 4709
rect 7558 4700 7564 4712
rect 7616 4700 7622 4752
rect 7742 4740 7748 4752
rect 7703 4712 7748 4740
rect 7742 4700 7748 4712
rect 7800 4700 7806 4752
rect 9309 4743 9367 4749
rect 9309 4709 9321 4743
rect 9355 4740 9367 4743
rect 9582 4740 9588 4752
rect 9355 4712 9588 4740
rect 9355 4709 9367 4712
rect 9309 4703 9367 4709
rect 2768 4675 2826 4681
rect 2768 4641 2780 4675
rect 2814 4672 2826 4675
rect 3602 4672 3608 4684
rect 2814 4644 3608 4672
rect 2814 4641 2826 4644
rect 2768 4635 2826 4641
rect 3602 4632 3608 4644
rect 3660 4632 3666 4684
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4672 5043 4675
rect 5166 4672 5172 4684
rect 5031 4644 5172 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5445 4675 5503 4681
rect 5445 4641 5457 4675
rect 5491 4672 5503 4675
rect 6178 4672 6184 4684
rect 5491 4644 6184 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 6288 4644 6377 4672
rect 2314 4604 2320 4616
rect 2275 4576 2320 4604
rect 2314 4564 2320 4576
rect 2372 4564 2378 4616
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4573 2559 4607
rect 4614 4604 4620 4616
rect 4575 4576 4620 4604
rect 2501 4567 2559 4573
rect 1578 4496 1584 4548
rect 1636 4536 1642 4548
rect 2130 4536 2136 4548
rect 1636 4508 2136 4536
rect 1636 4496 1642 4508
rect 2130 4496 2136 4508
rect 2188 4536 2194 4548
rect 2516 4536 2544 4567
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5276 4576 5549 4604
rect 2188 4508 2544 4536
rect 2188 4496 2194 4508
rect 3786 4496 3792 4548
rect 3844 4536 3850 4548
rect 5074 4536 5080 4548
rect 3844 4508 5080 4536
rect 3844 4496 3850 4508
rect 5074 4496 5080 4508
rect 5132 4496 5138 4548
rect 1673 4471 1731 4477
rect 1673 4437 1685 4471
rect 1719 4468 1731 4471
rect 2682 4468 2688 4480
rect 1719 4440 2688 4468
rect 1719 4437 1731 4440
rect 1673 4431 1731 4437
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4246 4468 4252 4480
rect 3927 4440 4252 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 5276 4468 5304 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 5684 4576 5729 4604
rect 5684 4564 5690 4576
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 6288 4536 6316 4644
rect 6365 4641 6377 4644
rect 6411 4641 6423 4675
rect 6914 4672 6920 4684
rect 6875 4644 6920 4672
rect 6365 4635 6423 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7576 4672 7604 4700
rect 7837 4675 7895 4681
rect 7837 4672 7849 4675
rect 7576 4644 7849 4672
rect 7837 4641 7849 4644
rect 7883 4641 7895 4675
rect 8478 4672 8484 4684
rect 7837 4635 7895 4641
rect 7944 4644 8484 4672
rect 6454 4604 6460 4616
rect 6415 4576 6460 4604
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 6932 4604 6960 4632
rect 7944 4604 7972 4644
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 9324 4672 9352 4703
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 9944 4743 10002 4749
rect 9944 4709 9956 4743
rect 9990 4740 10002 4743
rect 11238 4740 11244 4752
rect 9990 4712 11244 4740
rect 9990 4709 10002 4712
rect 9944 4703 10002 4709
rect 11238 4700 11244 4712
rect 11296 4700 11302 4752
rect 12434 4700 12440 4752
rect 12492 4740 12498 4752
rect 12492 4712 12537 4740
rect 12492 4700 12498 4712
rect 12618 4700 12624 4752
rect 12676 4740 12682 4752
rect 17402 4740 17408 4752
rect 12676 4712 17408 4740
rect 12676 4700 12682 4712
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 8619 4644 9352 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 13357 4675 13415 4681
rect 9548 4644 11744 4672
rect 9548 4632 9554 4644
rect 6932 4576 7972 4604
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 8294 4604 8300 4616
rect 8067 4576 8300 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8754 4604 8760 4616
rect 8588 4576 8760 4604
rect 8205 4539 8263 4545
rect 8205 4536 8217 4539
rect 5408 4508 6316 4536
rect 7300 4508 8217 4536
rect 5408 4496 5414 4508
rect 5718 4468 5724 4480
rect 5276 4440 5724 4468
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 5902 4468 5908 4480
rect 5863 4440 5908 4468
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 6270 4428 6276 4480
rect 6328 4468 6334 4480
rect 7300 4468 7328 4508
rect 8205 4505 8217 4508
rect 8251 4505 8263 4539
rect 8205 4499 8263 4505
rect 6328 4440 7328 4468
rect 6328 4428 6334 4440
rect 7374 4428 7380 4480
rect 7432 4468 7438 4480
rect 8588 4468 8616 4576
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 9398 4604 9404 4616
rect 9359 4576 9404 4604
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 9732 4576 9777 4604
rect 9732 4564 9738 4576
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 11716 4613 11744 4644
rect 13357 4641 13369 4675
rect 13403 4672 13415 4675
rect 13998 4672 14004 4684
rect 13403 4644 14004 4672
rect 13403 4641 13415 4644
rect 13357 4635 13415 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 14090 4632 14096 4684
rect 14148 4672 14154 4684
rect 14829 4675 14887 4681
rect 14829 4672 14841 4675
rect 14148 4644 14841 4672
rect 14148 4632 14154 4644
rect 14829 4641 14841 4644
rect 14875 4641 14887 4675
rect 14829 4635 14887 4641
rect 17589 4675 17647 4681
rect 17589 4641 17601 4675
rect 17635 4672 17647 4675
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17635 4644 17877 4672
rect 17635 4641 17647 4644
rect 17589 4635 17647 4641
rect 17865 4641 17877 4644
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 10744 4576 11621 4604
rect 10744 4564 10750 4576
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 12710 4604 12716 4616
rect 12671 4576 12716 4604
rect 11701 4567 11759 4573
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 13964 4576 14197 4604
rect 13964 4564 13970 4576
rect 8662 4496 8668 4548
rect 8720 4536 8726 4548
rect 9033 4539 9091 4545
rect 9033 4536 9045 4539
rect 8720 4508 9045 4536
rect 8720 4496 8726 4508
rect 9033 4505 9045 4508
rect 9079 4536 9091 4539
rect 9214 4536 9220 4548
rect 9079 4508 9220 4536
rect 9079 4505 9091 4508
rect 9033 4499 9091 4505
rect 9214 4496 9220 4508
rect 9272 4496 9278 4548
rect 12250 4536 12256 4548
rect 10888 4508 12256 4536
rect 7432 4440 8616 4468
rect 7432 4428 7438 4440
rect 9582 4428 9588 4480
rect 9640 4468 9646 4480
rect 10888 4468 10916 4508
rect 12250 4496 12256 4508
rect 12308 4496 12314 4548
rect 13354 4496 13360 4548
rect 13412 4536 13418 4548
rect 13556 4536 13584 4564
rect 13412 4508 13584 4536
rect 14108 4536 14136 4576
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 14274 4564 14280 4616
rect 14332 4604 14338 4616
rect 14844 4604 14872 4635
rect 18414 4604 18420 4616
rect 14332 4576 14377 4604
rect 14844 4576 18420 4604
rect 14332 4564 14338 4576
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 15013 4539 15071 4545
rect 15013 4536 15025 4539
rect 14108 4508 15025 4536
rect 13412 4496 13418 4508
rect 15013 4505 15025 4508
rect 15059 4505 15071 4539
rect 15013 4499 15071 4505
rect 11054 4468 11060 4480
rect 9640 4440 10916 4468
rect 11015 4440 11060 4468
rect 9640 4428 9646 4440
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11146 4428 11152 4480
rect 11204 4468 11210 4480
rect 12069 4471 12127 4477
rect 11204 4440 11249 4468
rect 11204 4428 11210 4440
rect 12069 4437 12081 4471
rect 12115 4468 12127 4471
rect 12434 4468 12440 4480
rect 12115 4440 12440 4468
rect 12115 4437 12127 4440
rect 12069 4431 12127 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 13538 4428 13544 4480
rect 13596 4468 13602 4480
rect 13814 4468 13820 4480
rect 13596 4440 13820 4468
rect 13596 4428 13602 4440
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 14642 4428 14648 4480
rect 14700 4468 14706 4480
rect 17589 4471 17647 4477
rect 17589 4468 17601 4471
rect 14700 4440 17601 4468
rect 14700 4428 14706 4440
rect 17589 4437 17601 4440
rect 17635 4468 17647 4471
rect 17681 4471 17739 4477
rect 17681 4468 17693 4471
rect 17635 4440 17693 4468
rect 17635 4437 17647 4440
rect 17589 4431 17647 4437
rect 17681 4437 17693 4440
rect 17727 4437 17739 4471
rect 18046 4468 18052 4480
rect 18007 4440 18052 4468
rect 17681 4431 17739 4437
rect 18046 4428 18052 4440
rect 18104 4428 18110 4480
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 3602 4264 3608 4276
rect 3563 4236 3608 4264
rect 3602 4224 3608 4236
rect 3660 4224 3666 4276
rect 5350 4264 5356 4276
rect 5311 4236 5356 4264
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 6420 4236 6837 4264
rect 6420 4224 6426 4236
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 6825 4227 6883 4233
rect 8754 4224 8760 4276
rect 8812 4264 8818 4276
rect 9033 4267 9091 4273
rect 9033 4264 9045 4267
rect 8812 4236 9045 4264
rect 8812 4224 8818 4236
rect 9033 4233 9045 4236
rect 9079 4233 9091 4267
rect 9033 4227 9091 4233
rect 9214 4224 9220 4276
rect 9272 4264 9278 4276
rect 9766 4264 9772 4276
rect 9272 4236 9772 4264
rect 9272 4224 9278 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 10229 4267 10287 4273
rect 10229 4233 10241 4267
rect 10275 4264 10287 4267
rect 10318 4264 10324 4276
rect 10275 4236 10324 4264
rect 10275 4233 10287 4236
rect 10229 4227 10287 4233
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 11974 4264 11980 4276
rect 11931 4236 11980 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12066 4224 12072 4276
rect 12124 4264 12130 4276
rect 12124 4236 12169 4264
rect 12124 4224 12130 4236
rect 12342 4224 12348 4276
rect 12400 4264 12406 4276
rect 12713 4267 12771 4273
rect 12713 4264 12725 4267
rect 12400 4236 12725 4264
rect 12400 4224 12406 4236
rect 12713 4233 12725 4236
rect 12759 4233 12771 4267
rect 12713 4227 12771 4233
rect 12802 4224 12808 4276
rect 12860 4264 12866 4276
rect 12860 4236 13952 4264
rect 12860 4224 12866 4236
rect 4890 4156 4896 4208
rect 4948 4196 4954 4208
rect 5261 4199 5319 4205
rect 5261 4196 5273 4199
rect 4948 4168 5273 4196
rect 4948 4156 4954 4168
rect 5261 4165 5273 4168
rect 5307 4196 5319 4199
rect 5442 4196 5448 4208
rect 5307 4168 5448 4196
rect 5307 4165 5319 4168
rect 5261 4159 5319 4165
rect 5442 4156 5448 4168
rect 5500 4196 5506 4208
rect 6454 4196 6460 4208
rect 5500 4168 6460 4196
rect 5500 4156 5506 4168
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 9125 4199 9183 4205
rect 9125 4165 9137 4199
rect 9171 4196 9183 4199
rect 9398 4196 9404 4208
rect 9171 4168 9404 4196
rect 9171 4165 9183 4168
rect 9125 4159 9183 4165
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 9508 4168 9720 4196
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 5626 4128 5632 4140
rect 5408 4100 5632 4128
rect 5408 4088 5414 4100
rect 5626 4088 5632 4100
rect 5684 4128 5690 4140
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5684 4100 5917 4128
rect 5684 4088 5690 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 6178 4128 6184 4140
rect 6139 4100 6184 4128
rect 5905 4091 5963 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 7374 4128 7380 4140
rect 7335 4100 7380 4128
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7484 4100 7788 4128
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4029 1731 4063
rect 1673 4023 1731 4029
rect 1486 3952 1492 4004
rect 1544 3992 1550 4004
rect 1688 3992 1716 4023
rect 2130 4020 2136 4072
rect 2188 4060 2194 4072
rect 2225 4063 2283 4069
rect 2225 4060 2237 4063
rect 2188 4032 2237 4060
rect 2188 4020 2194 4032
rect 2225 4029 2237 4032
rect 2271 4029 2283 4063
rect 2225 4023 2283 4029
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 2481 4063 2539 4069
rect 2481 4060 2493 4063
rect 2372 4032 2493 4060
rect 2372 4020 2378 4032
rect 2481 4029 2493 4032
rect 2527 4029 2539 4063
rect 3786 4060 3792 4072
rect 3747 4032 3792 4060
rect 2481 4023 2539 4029
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 3878 4020 3884 4072
rect 3936 4060 3942 4072
rect 5166 4060 5172 4072
rect 3936 4032 5172 4060
rect 3936 4020 3942 4032
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 5810 4060 5816 4072
rect 5723 4032 5816 4060
rect 5810 4020 5816 4032
rect 5868 4060 5874 4072
rect 7484 4060 7512 4100
rect 7650 4060 7656 4072
rect 5868 4032 7512 4060
rect 7611 4032 7656 4060
rect 5868 4020 5874 4032
rect 7650 4020 7656 4032
rect 7708 4020 7714 4072
rect 7760 4060 7788 4100
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9508 4128 9536 4168
rect 9692 4137 9720 4168
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 13078 4196 13084 4208
rect 11664 4168 13084 4196
rect 11664 4156 11670 4168
rect 13078 4156 13084 4168
rect 13136 4156 13142 4208
rect 13541 4199 13599 4205
rect 13541 4165 13553 4199
rect 13587 4196 13599 4199
rect 13924 4196 13952 4236
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14369 4267 14427 4273
rect 14369 4264 14381 4267
rect 14056 4236 14381 4264
rect 14056 4224 14062 4236
rect 14369 4233 14381 4236
rect 14415 4233 14427 4267
rect 14369 4227 14427 4233
rect 14458 4224 14464 4276
rect 14516 4264 14522 4276
rect 17954 4264 17960 4276
rect 14516 4236 17960 4264
rect 14516 4224 14522 4236
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 18414 4264 18420 4276
rect 18375 4236 18420 4264
rect 18414 4224 18420 4236
rect 18472 4224 18478 4276
rect 13587 4168 13768 4196
rect 13924 4168 17816 4196
rect 13587 4165 13599 4168
rect 13541 4159 13599 4165
rect 8996 4100 9536 4128
rect 9677 4131 9735 4137
rect 8996 4088 9002 4100
rect 9677 4097 9689 4131
rect 9723 4097 9735 4131
rect 13354 4128 13360 4140
rect 9677 4091 9735 4097
rect 9876 4100 10640 4128
rect 13315 4100 13360 4128
rect 9306 4060 9312 4072
rect 7760 4032 9312 4060
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9585 4063 9643 4069
rect 9456 4032 9536 4060
rect 9456 4020 9462 4032
rect 4148 3995 4206 4001
rect 1544 3964 2176 3992
rect 1544 3952 1550 3964
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 2038 3924 2044 3936
rect 1999 3896 2044 3924
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 2148 3924 2176 3964
rect 4148 3961 4160 3995
rect 4194 3992 4206 3995
rect 4246 3992 4252 4004
rect 4194 3964 4252 3992
rect 4194 3961 4206 3964
rect 4148 3955 4206 3961
rect 4246 3952 4252 3964
rect 4304 3992 4310 4004
rect 5350 3992 5356 4004
rect 4304 3964 5356 3992
rect 4304 3952 4310 3964
rect 5350 3952 5356 3964
rect 5408 3952 5414 4004
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 7742 3992 7748 4004
rect 7239 3964 7748 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 7742 3952 7748 3964
rect 7800 3952 7806 4004
rect 7920 3995 7978 4001
rect 7920 3961 7932 3995
rect 7966 3961 7978 3995
rect 7920 3955 7978 3961
rect 4338 3924 4344 3936
rect 2148 3896 4344 3924
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 5721 3927 5779 3933
rect 5721 3893 5733 3927
rect 5767 3924 5779 3927
rect 6086 3924 6092 3936
rect 5767 3896 6092 3924
rect 5767 3893 5779 3896
rect 5721 3887 5779 3893
rect 6086 3884 6092 3896
rect 6144 3924 6150 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 6144 3896 6561 3924
rect 6144 3884 6150 3896
rect 6549 3893 6561 3896
rect 6595 3924 6607 3927
rect 6730 3924 6736 3936
rect 6595 3896 6736 3924
rect 6595 3893 6607 3896
rect 6549 3887 6607 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7285 3927 7343 3933
rect 7285 3893 7297 3927
rect 7331 3924 7343 3927
rect 7374 3924 7380 3936
rect 7331 3896 7380 3924
rect 7331 3893 7343 3896
rect 7285 3887 7343 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7935 3924 7963 3955
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 9508 3992 9536 4032
rect 9585 4029 9597 4063
rect 9631 4060 9643 4063
rect 9876 4060 9904 4100
rect 9631 4032 9904 4060
rect 9631 4029 9643 4032
rect 9585 4023 9643 4029
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 10008 4032 10517 4060
rect 10008 4020 10014 4032
rect 10505 4029 10517 4032
rect 10551 4029 10563 4063
rect 10612 4060 10640 4100
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 10772 4063 10830 4069
rect 10612 4032 10732 4060
rect 10505 4023 10563 4029
rect 10594 3992 10600 4004
rect 9272 3964 9444 3992
rect 9508 3964 10600 3992
rect 9272 3952 9278 3964
rect 8294 3924 8300 3936
rect 7935 3896 8300 3924
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 9416 3924 9444 3964
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 10704 3992 10732 4032
rect 10772 4029 10784 4063
rect 10818 4060 10830 4063
rect 11054 4060 11060 4072
rect 10818 4032 11060 4060
rect 10818 4029 10830 4032
rect 10772 4023 10830 4029
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11882 4020 11888 4072
rect 11940 4020 11946 4072
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4060 13139 4063
rect 13630 4060 13636 4072
rect 13127 4032 13636 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 11900 3992 11928 4020
rect 10704 3964 11928 3992
rect 13173 3995 13231 4001
rect 13173 3961 13185 3995
rect 13219 3992 13231 3995
rect 13538 3992 13544 4004
rect 13219 3964 13544 3992
rect 13219 3961 13231 3964
rect 13173 3955 13231 3961
rect 13538 3952 13544 3964
rect 13596 3952 13602 4004
rect 13740 3992 13768 4168
rect 14090 4128 14096 4140
rect 14051 4100 14096 4128
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 15010 4128 15016 4140
rect 14971 4100 15016 4128
rect 15010 4088 15016 4100
rect 15068 4088 15074 4140
rect 17788 4137 17816 4168
rect 17773 4131 17831 4137
rect 17773 4097 17785 4131
rect 17819 4128 17831 4131
rect 17819 4100 18092 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 13906 4060 13912 4072
rect 13867 4032 13912 4060
rect 13906 4020 13912 4032
rect 13964 4020 13970 4072
rect 13998 4020 14004 4072
rect 14056 4060 14062 4072
rect 17954 4060 17960 4072
rect 14056 4032 17960 4060
rect 14056 4020 14062 4032
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 18064 4069 18092 4100
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 14829 3995 14887 4001
rect 14829 3992 14841 3995
rect 13740 3964 14841 3992
rect 14829 3961 14841 3964
rect 14875 3961 14887 3995
rect 14829 3955 14887 3961
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 9416 3896 9505 3924
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 9582 3884 9588 3936
rect 9640 3924 9646 3936
rect 9953 3927 10011 3933
rect 9953 3924 9965 3927
rect 9640 3896 9965 3924
rect 9640 3884 9646 3896
rect 9953 3893 9965 3896
rect 9999 3893 10011 3927
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 9953 3887 10011 3893
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 12618 3924 12624 3936
rect 12531 3896 12624 3924
rect 12618 3884 12624 3896
rect 12676 3924 12682 3936
rect 13998 3924 14004 3936
rect 12676 3896 14004 3924
rect 12676 3884 12682 3896
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3924 14795 3927
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 14783 3896 15301 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 15289 3893 15301 3896
rect 15335 3924 15347 3927
rect 15378 3924 15384 3936
rect 15335 3896 15384 3924
rect 15335 3893 15347 3896
rect 15289 3887 15347 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2961 3723 3019 3729
rect 2004 3692 2452 3720
rect 2004 3680 2010 3692
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 1673 3587 1731 3593
rect 1673 3584 1685 3587
rect 1627 3556 1685 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 1673 3553 1685 3556
rect 1719 3553 1731 3587
rect 1673 3547 1731 3553
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3584 2099 3587
rect 2314 3584 2320 3596
rect 2087 3556 2320 3584
rect 2087 3553 2099 3556
rect 2041 3547 2099 3553
rect 1688 3516 1716 3547
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 2424 3593 2452 3692
rect 2961 3689 2973 3723
rect 3007 3720 3019 3723
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 3007 3692 4537 3720
rect 3007 3689 3019 3692
rect 2961 3683 3019 3689
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 4525 3683 4583 3689
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 6089 3723 6147 3729
rect 6089 3720 6101 3723
rect 5960 3692 6101 3720
rect 5960 3680 5966 3692
rect 6089 3689 6101 3692
rect 6135 3689 6147 3723
rect 6089 3683 6147 3689
rect 6638 3680 6644 3732
rect 6696 3720 6702 3732
rect 6733 3723 6791 3729
rect 6733 3720 6745 3723
rect 6696 3692 6745 3720
rect 6696 3680 6702 3692
rect 6733 3689 6745 3692
rect 6779 3689 6791 3723
rect 7374 3720 7380 3732
rect 7335 3692 7380 3720
rect 6733 3683 6791 3689
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 8386 3720 8392 3732
rect 7760 3692 8392 3720
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 3418 3652 3424 3664
rect 2915 3624 3424 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 3418 3612 3424 3624
rect 3476 3652 3482 3664
rect 3476 3624 3556 3652
rect 3476 3612 3482 3624
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3553 2467 3587
rect 3326 3584 3332 3596
rect 3287 3556 3332 3584
rect 2409 3547 2467 3553
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3528 3584 3556 3624
rect 3694 3612 3700 3664
rect 3752 3652 3758 3664
rect 5261 3655 5319 3661
rect 5261 3652 5273 3655
rect 3752 3624 5273 3652
rect 3752 3612 3758 3624
rect 5261 3621 5273 3624
rect 5307 3652 5319 3655
rect 7009 3655 7067 3661
rect 7009 3652 7021 3655
rect 5307 3624 7021 3652
rect 5307 3621 5319 3624
rect 5261 3615 5319 3621
rect 7009 3621 7021 3624
rect 7055 3652 7067 3655
rect 7282 3652 7288 3664
rect 7055 3624 7288 3652
rect 7055 3621 7067 3624
rect 7009 3615 7067 3621
rect 7282 3612 7288 3624
rect 7340 3612 7346 3664
rect 3786 3584 3792 3596
rect 3528 3556 3792 3584
rect 3786 3544 3792 3556
rect 3844 3544 3850 3596
rect 4430 3584 4436 3596
rect 4391 3556 4436 3584
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7760 3593 7788 3692
rect 8386 3680 8392 3692
rect 8444 3720 8450 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8444 3692 9045 3720
rect 8444 3680 8450 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9033 3683 9091 3689
rect 9122 3680 9128 3732
rect 9180 3720 9186 3732
rect 10318 3720 10324 3732
rect 9180 3692 10324 3720
rect 9180 3680 9186 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 10413 3723 10471 3729
rect 10413 3689 10425 3723
rect 10459 3720 10471 3723
rect 10965 3723 11023 3729
rect 10965 3720 10977 3723
rect 10459 3692 10977 3720
rect 10459 3689 10471 3692
rect 10413 3683 10471 3689
rect 10965 3689 10977 3692
rect 11011 3689 11023 3723
rect 10965 3683 11023 3689
rect 11333 3723 11391 3729
rect 11333 3689 11345 3723
rect 11379 3720 11391 3723
rect 11379 3692 12204 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 12176 3664 12204 3692
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 14737 3723 14795 3729
rect 14737 3720 14749 3723
rect 14700 3692 14749 3720
rect 14700 3680 14706 3692
rect 14737 3689 14749 3692
rect 14783 3689 14795 3723
rect 17678 3720 17684 3732
rect 17639 3692 17684 3720
rect 14737 3683 14795 3689
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 8665 3655 8723 3661
rect 8665 3621 8677 3655
rect 8711 3652 8723 3655
rect 8938 3652 8944 3664
rect 8711 3624 8944 3652
rect 8711 3621 8723 3624
rect 8665 3615 8723 3621
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 9306 3612 9312 3664
rect 9364 3652 9370 3664
rect 9401 3655 9459 3661
rect 9401 3652 9413 3655
rect 9364 3624 9413 3652
rect 9364 3612 9370 3624
rect 9401 3621 9413 3624
rect 9447 3621 9459 3655
rect 9401 3615 9459 3621
rect 9674 3612 9680 3664
rect 9732 3652 9738 3664
rect 11974 3652 11980 3664
rect 9732 3624 11980 3652
rect 9732 3612 9738 3624
rect 11974 3612 11980 3624
rect 12032 3661 12038 3664
rect 12032 3655 12096 3661
rect 12032 3621 12050 3655
rect 12084 3621 12096 3655
rect 12032 3615 12096 3621
rect 12032 3612 12038 3615
rect 12158 3612 12164 3664
rect 12216 3612 12222 3664
rect 13532 3655 13590 3661
rect 13532 3621 13544 3655
rect 13578 3652 13590 3655
rect 14090 3652 14096 3664
rect 13578 3624 14096 3652
rect 13578 3621 13590 3624
rect 13532 3615 13590 3621
rect 7745 3587 7803 3593
rect 7745 3584 7757 3587
rect 7524 3556 7757 3584
rect 7524 3544 7530 3556
rect 7745 3553 7757 3556
rect 7791 3553 7803 3587
rect 8110 3584 8116 3596
rect 7745 3547 7803 3553
rect 7852 3556 8116 3584
rect 1688 3488 3004 3516
rect 2593 3451 2651 3457
rect 2593 3417 2605 3451
rect 2639 3448 2651 3451
rect 2866 3448 2872 3460
rect 2639 3420 2872 3448
rect 2639 3417 2651 3420
rect 2593 3411 2651 3417
rect 2866 3408 2872 3420
rect 2924 3408 2930 3460
rect 2976 3448 3004 3488
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 3108 3488 3433 3516
rect 3108 3476 3114 3488
rect 3421 3485 3433 3488
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 4154 3516 4160 3528
rect 3651 3488 4160 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3516 4767 3519
rect 4890 3516 4896 3528
rect 4755 3488 4896 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5258 3516 5264 3528
rect 5132 3488 5264 3516
rect 5132 3476 5138 3488
rect 5258 3476 5264 3488
rect 5316 3516 5322 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5316 3488 5365 3516
rect 5316 3476 5322 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3516 5595 3519
rect 5810 3516 5816 3528
rect 5583 3488 5816 3516
rect 5583 3485 5595 3488
rect 5537 3479 5595 3485
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3516 6423 3519
rect 6546 3516 6552 3528
rect 6411 3488 6552 3516
rect 6411 3485 6423 3488
rect 6365 3479 6423 3485
rect 3694 3448 3700 3460
rect 2976 3420 3700 3448
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 3878 3448 3884 3460
rect 3839 3420 3884 3448
rect 3878 3408 3884 3420
rect 3936 3408 3942 3460
rect 4065 3451 4123 3457
rect 4065 3417 4077 3451
rect 4111 3448 4123 3451
rect 6196 3448 6224 3479
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 7852 3525 7880 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 8573 3587 8631 3593
rect 8573 3584 8585 3587
rect 8536 3556 8585 3584
rect 8536 3544 8542 3556
rect 8573 3553 8585 3556
rect 8619 3584 8631 3587
rect 9217 3587 9275 3593
rect 9217 3584 9229 3587
rect 8619 3556 9229 3584
rect 8619 3553 8631 3556
rect 8573 3547 8631 3553
rect 9217 3553 9229 3556
rect 9263 3584 9275 3587
rect 10226 3584 10232 3596
rect 9263 3556 10232 3584
rect 9263 3553 9275 3556
rect 9217 3547 9275 3553
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 10410 3584 10416 3596
rect 10367 3556 10416 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 11425 3587 11483 3593
rect 11425 3584 11437 3587
rect 10919 3556 11437 3584
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3516 7343 3519
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 7331 3488 7849 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 7837 3485 7849 3488
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3516 8079 3519
rect 8294 3516 8300 3528
rect 8067 3488 8300 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 8294 3476 8300 3488
rect 8352 3516 8358 3528
rect 8757 3519 8815 3525
rect 8757 3516 8769 3519
rect 8352 3488 8769 3516
rect 8352 3476 8358 3488
rect 8757 3485 8769 3488
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 10502 3516 10508 3528
rect 8996 3488 10508 3516
rect 8996 3476 9002 3488
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3516 10655 3519
rect 11238 3516 11244 3528
rect 10643 3488 11244 3516
rect 10643 3485 10655 3488
rect 10597 3479 10655 3485
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 4111 3420 4292 3448
rect 4111 3417 4123 3420
rect 4065 3411 4123 3417
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 2222 3380 2228 3392
rect 2183 3352 2228 3380
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 4264 3380 4292 3420
rect 4448 3420 6224 3448
rect 4448 3380 4476 3420
rect 7742 3408 7748 3460
rect 7800 3448 7806 3460
rect 8205 3451 8263 3457
rect 8205 3448 8217 3451
rect 7800 3420 8217 3448
rect 7800 3408 7806 3420
rect 8205 3417 8217 3420
rect 8251 3417 8263 3451
rect 11348 3448 11376 3556
rect 11425 3553 11437 3556
rect 11471 3584 11483 3587
rect 12894 3584 12900 3596
rect 11471 3556 12900 3584
rect 11471 3553 11483 3556
rect 11425 3547 11483 3553
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 13547 3584 13575 3615
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 17497 3587 17555 3593
rect 17497 3584 17509 3587
rect 13096 3556 13575 3584
rect 17144 3556 17509 3584
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11793 3519 11851 3525
rect 11572 3488 11617 3516
rect 11572 3476 11578 3488
rect 11793 3485 11805 3519
rect 11839 3485 11851 3519
rect 11793 3479 11851 3485
rect 8205 3411 8263 3417
rect 9600 3420 11376 3448
rect 4890 3380 4896 3392
rect 4264 3352 4476 3380
rect 4851 3352 4896 3380
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5721 3383 5779 3389
rect 5721 3380 5733 3383
rect 5040 3352 5733 3380
rect 5040 3340 5046 3352
rect 5721 3349 5733 3352
rect 5767 3349 5779 3383
rect 5721 3343 5779 3349
rect 6362 3340 6368 3392
rect 6420 3380 6426 3392
rect 6549 3383 6607 3389
rect 6549 3380 6561 3383
rect 6420 3352 6561 3380
rect 6420 3340 6426 3352
rect 6549 3349 6561 3352
rect 6595 3349 6607 3383
rect 6549 3343 6607 3349
rect 6638 3340 6644 3392
rect 6696 3380 6702 3392
rect 9600 3380 9628 3420
rect 9766 3380 9772 3392
rect 6696 3352 9628 3380
rect 9727 3352 9772 3380
rect 6696 3340 6702 3352
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 9953 3383 10011 3389
rect 9953 3349 9965 3383
rect 9999 3380 10011 3383
rect 10318 3380 10324 3392
rect 9999 3352 10324 3380
rect 9999 3349 10011 3352
rect 9953 3343 10011 3349
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 11808 3380 11836 3479
rect 13096 3448 13124 3556
rect 17144 3528 17172 3556
rect 17497 3553 17509 3556
rect 17543 3553 17555 3587
rect 17497 3547 17555 3553
rect 17865 3587 17923 3593
rect 17865 3553 17877 3587
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 18414 3584 18420 3596
rect 18279 3556 18420 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 13262 3516 13268 3528
rect 13223 3488 13268 3516
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 17126 3516 17132 3528
rect 17087 3488 17132 3516
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 17880 3516 17908 3547
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 17328 3488 17908 3516
rect 13173 3451 13231 3457
rect 13173 3448 13185 3451
rect 13096 3420 13185 3448
rect 13173 3417 13185 3420
rect 13219 3417 13231 3451
rect 13173 3411 13231 3417
rect 13280 3380 13308 3476
rect 14645 3451 14703 3457
rect 14645 3417 14657 3451
rect 14691 3448 14703 3451
rect 15010 3448 15016 3460
rect 14691 3420 15016 3448
rect 14691 3417 14703 3420
rect 14645 3411 14703 3417
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 11808 3352 13308 3380
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 17328 3389 17356 3488
rect 17313 3383 17371 3389
rect 17313 3380 17325 3383
rect 13688 3352 17325 3380
rect 13688 3340 13694 3352
rect 17313 3349 17325 3352
rect 17359 3349 17371 3383
rect 17313 3343 17371 3349
rect 17862 3340 17868 3392
rect 17920 3380 17926 3392
rect 18049 3383 18107 3389
rect 18049 3380 18061 3383
rect 17920 3352 18061 3380
rect 17920 3340 17926 3352
rect 18049 3349 18061 3352
rect 18095 3349 18107 3383
rect 18414 3380 18420 3392
rect 18375 3352 18420 3380
rect 18049 3343 18107 3349
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 2590 3176 2596 3188
rect 2551 3148 2596 3176
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 3050 3176 3056 3188
rect 3011 3148 3056 3176
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3881 3179 3939 3185
rect 3881 3176 3893 3179
rect 3384 3148 3893 3176
rect 3384 3136 3390 3148
rect 3881 3145 3893 3148
rect 3927 3145 3939 3179
rect 5810 3176 5816 3188
rect 3881 3139 3939 3145
rect 4264 3148 5816 3176
rect 2317 3111 2375 3117
rect 2317 3077 2329 3111
rect 2363 3108 2375 3111
rect 2774 3108 2780 3120
rect 2363 3080 2780 3108
rect 2363 3077 2375 3080
rect 2317 3071 2375 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 2869 3111 2927 3117
rect 2869 3077 2881 3111
rect 2915 3108 2927 3111
rect 3142 3108 3148 3120
rect 2915 3080 3148 3108
rect 2915 3077 2927 3080
rect 2869 3071 2927 3077
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 3602 3040 3608 3052
rect 3563 3012 3608 3040
rect 3602 3000 3608 3012
rect 3660 3040 3666 3052
rect 4264 3040 4292 3148
rect 4338 3068 4344 3120
rect 4396 3068 4402 3120
rect 3660 3012 4292 3040
rect 3660 3000 3666 3012
rect 1394 2932 1400 2984
rect 1452 2972 1458 2984
rect 1452 2944 1532 2972
rect 1452 2932 1458 2944
rect 1504 2904 1532 2944
rect 1578 2932 1584 2984
rect 1636 2972 1642 2984
rect 1636 2944 1681 2972
rect 1636 2932 1642 2944
rect 2038 2932 2044 2984
rect 2096 2972 2102 2984
rect 2133 2975 2191 2981
rect 2133 2972 2145 2975
rect 2096 2944 2145 2972
rect 2096 2932 2102 2944
rect 2133 2941 2145 2944
rect 2179 2941 2191 2975
rect 2133 2935 2191 2941
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2941 2743 2975
rect 3418 2972 3424 2984
rect 3379 2944 3424 2972
rect 2685 2935 2743 2941
rect 1857 2907 1915 2913
rect 1857 2904 1869 2907
rect 1504 2876 1869 2904
rect 1857 2873 1869 2876
rect 1903 2873 1915 2907
rect 2700 2904 2728 2935
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 4356 2981 4384 3068
rect 4448 3049 4476 3148
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 6546 3176 6552 3188
rect 6507 3148 6552 3176
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 8205 3179 8263 3185
rect 6788 3148 7788 3176
rect 6788 3136 6794 3148
rect 4709 3111 4767 3117
rect 4709 3077 4721 3111
rect 4755 3108 4767 3111
rect 5074 3108 5080 3120
rect 4755 3080 5080 3108
rect 4755 3077 4767 3080
rect 4709 3071 4767 3077
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3009 4491 3043
rect 5166 3040 5172 3052
rect 5127 3012 5172 3040
rect 4433 3003 4491 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 6564 3040 6592 3136
rect 7760 3108 7788 3148
rect 8205 3145 8217 3179
rect 8251 3176 8263 3179
rect 8294 3176 8300 3188
rect 8251 3148 8300 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 8938 3176 8944 3188
rect 8435 3148 8944 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 10410 3136 10416 3188
rect 10468 3176 10474 3188
rect 13998 3176 14004 3188
rect 10468 3148 14004 3176
rect 10468 3136 10474 3148
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 17402 3176 17408 3188
rect 17363 3148 17408 3176
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 10870 3108 10876 3120
rect 7760 3080 10876 3108
rect 10870 3068 10876 3080
rect 10928 3068 10934 3120
rect 12250 3108 12256 3120
rect 11164 3080 12256 3108
rect 8757 3043 8815 3049
rect 6564 3012 6960 3040
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2972 5043 2975
rect 5074 2972 5080 2984
rect 5031 2944 5080 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 5074 2932 5080 2944
rect 5132 2972 5138 2984
rect 5994 2972 6000 2984
rect 5132 2944 6000 2972
rect 5132 2932 5138 2944
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2941 6883 2975
rect 6932 2972 6960 3012
rect 8757 3009 8769 3043
rect 8803 3040 8815 3043
rect 9398 3040 9404 3052
rect 8803 3012 9404 3040
rect 8803 3009 8815 3012
rect 8757 3003 8815 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 9674 3040 9680 3052
rect 9635 3012 9680 3040
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 10318 3040 10324 3052
rect 10279 3012 10324 3040
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 11054 3040 11060 3052
rect 10551 3012 11060 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 7081 2975 7139 2981
rect 7081 2972 7093 2975
rect 6932 2944 7093 2972
rect 6825 2935 6883 2941
rect 7081 2941 7093 2944
rect 7127 2941 7139 2975
rect 7081 2935 7139 2941
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 8527 2944 9076 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 5442 2913 5448 2916
rect 5436 2904 5448 2913
rect 1857 2867 1915 2873
rect 2516 2876 3648 2904
rect 5403 2876 5448 2904
rect 1489 2839 1547 2845
rect 1489 2805 1501 2839
rect 1535 2836 1547 2839
rect 2516 2836 2544 2876
rect 1535 2808 2544 2836
rect 1535 2805 1547 2808
rect 1489 2799 1547 2805
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 3513 2839 3571 2845
rect 3513 2836 3525 2839
rect 2648 2808 3525 2836
rect 2648 2796 2654 2808
rect 3513 2805 3525 2808
rect 3559 2805 3571 2839
rect 3620 2836 3648 2876
rect 5436 2867 5448 2876
rect 5442 2864 5448 2867
rect 5500 2864 5506 2916
rect 6840 2904 6868 2935
rect 7650 2904 7656 2916
rect 6840 2876 7656 2904
rect 7650 2864 7656 2876
rect 7708 2864 7714 2916
rect 4249 2839 4307 2845
rect 4249 2836 4261 2839
rect 3620 2808 4261 2836
rect 3513 2799 3571 2805
rect 4249 2805 4261 2808
rect 4295 2836 4307 2839
rect 4706 2836 4712 2848
rect 4295 2808 4712 2836
rect 4295 2805 4307 2808
rect 4249 2799 4307 2805
rect 4706 2796 4712 2808
rect 4764 2836 4770 2848
rect 6362 2836 6368 2848
rect 4764 2808 6368 2836
rect 4764 2796 4770 2808
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 9048 2845 9076 2944
rect 10410 2932 10416 2984
rect 10468 2972 10474 2984
rect 11164 2981 11192 3080
rect 12250 3068 12256 3080
rect 12308 3108 12314 3120
rect 12989 3111 13047 3117
rect 12989 3108 13001 3111
rect 12308 3080 13001 3108
rect 12308 3068 12314 3080
rect 12989 3077 13001 3080
rect 13035 3108 13047 3111
rect 13449 3111 13507 3117
rect 13035 3080 13400 3108
rect 13035 3077 13047 3080
rect 12989 3071 13047 3077
rect 11425 3043 11483 3049
rect 11425 3009 11437 3043
rect 11471 3009 11483 3043
rect 11882 3040 11888 3052
rect 11843 3012 11888 3040
rect 11425 3003 11483 3009
rect 11149 2975 11207 2981
rect 10468 2944 10916 2972
rect 10468 2932 10474 2944
rect 9401 2907 9459 2913
rect 9401 2873 9413 2907
rect 9447 2904 9459 2907
rect 9950 2904 9956 2916
rect 9447 2876 9956 2904
rect 9447 2873 9459 2876
rect 9401 2867 9459 2873
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 10229 2907 10287 2913
rect 10229 2873 10241 2907
rect 10275 2904 10287 2907
rect 10888 2904 10916 2944
rect 11149 2941 11161 2975
rect 11195 2941 11207 2975
rect 11440 2972 11468 3003
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 12526 3000 12532 3052
rect 12584 3040 12590 3052
rect 13173 3043 13231 3049
rect 13173 3040 13185 3043
rect 12584 3012 13185 3040
rect 12584 3000 12590 3012
rect 13173 3009 13185 3012
rect 13219 3009 13231 3043
rect 13372 3040 13400 3080
rect 13449 3077 13461 3111
rect 13495 3108 13507 3111
rect 14366 3108 14372 3120
rect 13495 3080 14372 3108
rect 13495 3077 13507 3080
rect 13449 3071 13507 3077
rect 13630 3040 13636 3052
rect 13372 3012 13636 3040
rect 13173 3003 13231 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 11514 2972 11520 2984
rect 11440 2944 11520 2972
rect 11149 2935 11207 2941
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2972 11759 2975
rect 11790 2972 11796 2984
rect 11747 2944 11796 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12400 2944 12449 2972
rect 12400 2932 12406 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12713 2907 12771 2913
rect 12713 2904 12725 2907
rect 10275 2876 10824 2904
rect 10888 2876 12725 2904
rect 10275 2873 10287 2876
rect 10229 2867 10287 2873
rect 10796 2845 10824 2876
rect 12713 2873 12725 2876
rect 12759 2873 12771 2907
rect 12713 2867 12771 2873
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2805 9091 2839
rect 9033 2799 9091 2805
rect 9493 2839 9551 2845
rect 9493 2805 9505 2839
rect 9539 2836 9551 2839
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 9539 2808 9873 2836
rect 9539 2805 9551 2808
rect 9493 2799 9551 2805
rect 9861 2805 9873 2808
rect 9907 2805 9919 2839
rect 9861 2799 9919 2805
rect 10781 2839 10839 2845
rect 10781 2805 10793 2839
rect 10827 2805 10839 2839
rect 10781 2799 10839 2805
rect 11241 2839 11299 2845
rect 11241 2805 11253 2839
rect 11287 2836 11299 2839
rect 13740 2836 13768 3080
rect 14366 3068 14372 3080
rect 14424 3068 14430 3120
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 15378 2932 15384 2984
rect 15436 2972 15442 2984
rect 16761 2975 16819 2981
rect 16761 2972 16773 2975
rect 15436 2944 16773 2972
rect 15436 2932 15442 2944
rect 16761 2941 16773 2944
rect 16807 2972 16819 2975
rect 16853 2975 16911 2981
rect 16853 2972 16865 2975
rect 16807 2944 16865 2972
rect 16807 2941 16819 2944
rect 16761 2935 16819 2941
rect 16853 2941 16865 2944
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 17589 2975 17647 2981
rect 17589 2972 17601 2975
rect 17460 2944 17601 2972
rect 17460 2932 17466 2944
rect 17589 2941 17601 2944
rect 17635 2941 17647 2975
rect 17589 2935 17647 2941
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 18012 2944 18061 2972
rect 18012 2932 18018 2944
rect 18049 2941 18061 2944
rect 18095 2972 18107 2975
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 18095 2944 18429 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 14461 2907 14519 2913
rect 14461 2873 14473 2907
rect 14507 2904 14519 2907
rect 14826 2904 14832 2916
rect 14507 2876 14832 2904
rect 14507 2873 14519 2876
rect 14461 2867 14519 2873
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 14918 2864 14924 2916
rect 14976 2904 14982 2916
rect 19426 2904 19432 2916
rect 14976 2876 19432 2904
rect 14976 2864 14982 2876
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 17034 2836 17040 2848
rect 11287 2808 13768 2836
rect 16995 2808 17040 2836
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 17770 2836 17776 2848
rect 17731 2808 17776 2836
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18230 2836 18236 2848
rect 18191 2808 18236 2836
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 1486 2632 1492 2644
rect 1447 2604 1492 2632
rect 1486 2592 1492 2604
rect 1544 2592 1550 2644
rect 4430 2592 4436 2644
rect 4488 2632 4494 2644
rect 4709 2635 4767 2641
rect 4709 2632 4721 2635
rect 4488 2604 4721 2632
rect 4488 2592 4494 2604
rect 4709 2601 4721 2604
rect 4755 2601 4767 2635
rect 5074 2632 5080 2644
rect 5035 2604 5080 2632
rect 4709 2595 4767 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 8202 2632 8208 2644
rect 6104 2604 8208 2632
rect 4890 2524 4896 2576
rect 4948 2564 4954 2576
rect 5169 2567 5227 2573
rect 5169 2564 5181 2567
rect 4948 2536 5181 2564
rect 4948 2524 4954 2536
rect 5169 2533 5181 2536
rect 5215 2533 5227 2567
rect 5169 2527 5227 2533
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2496 1639 2499
rect 1670 2496 1676 2508
rect 1627 2468 1676 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 2130 2496 2136 2508
rect 2091 2468 2136 2496
rect 2130 2456 2136 2468
rect 2188 2456 2194 2508
rect 2682 2496 2688 2508
rect 2643 2468 2688 2496
rect 2682 2456 2688 2468
rect 2740 2456 2746 2508
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 3418 2496 3424 2508
rect 3283 2468 3424 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 3605 2499 3663 2505
rect 3605 2465 3617 2499
rect 3651 2465 3663 2499
rect 3605 2459 3663 2465
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4982 2496 4988 2508
rect 4111 2468 4988 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 1210 2388 1216 2440
rect 1268 2428 1274 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1268 2400 1777 2428
rect 1268 2388 1274 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 1765 2391 1823 2397
rect 2148 2400 2329 2428
rect 2148 2372 2176 2400
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 3050 2428 3056 2440
rect 3007 2400 3056 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 2130 2320 2136 2372
rect 2188 2320 2194 2372
rect 3620 2360 3648 2459
rect 4982 2456 4988 2468
rect 5040 2456 5046 2508
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 6104 2505 6132 2604
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 9950 2632 9956 2644
rect 9911 2604 9956 2632
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 10459 2604 10793 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 10781 2595 10839 2601
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11422 2632 11428 2644
rect 11287 2604 11428 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 11609 2635 11667 2641
rect 11609 2601 11621 2635
rect 11655 2601 11667 2635
rect 11609 2595 11667 2601
rect 6730 2524 6736 2576
rect 6788 2564 6794 2576
rect 8297 2567 8355 2573
rect 8297 2564 8309 2567
rect 6788 2536 8309 2564
rect 6788 2524 6794 2536
rect 8297 2533 8309 2536
rect 8343 2533 8355 2567
rect 9030 2564 9036 2576
rect 8297 2527 8355 2533
rect 8404 2536 9036 2564
rect 6089 2499 6147 2505
rect 6089 2465 6101 2499
rect 6135 2465 6147 2499
rect 6914 2496 6920 2508
rect 6875 2468 6920 2496
rect 6089 2459 6147 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7834 2456 7840 2508
rect 7892 2496 7898 2508
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7892 2468 8033 2496
rect 7892 2456 7898 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 8404 2496 8432 2536
rect 9030 2524 9036 2536
rect 9088 2524 9094 2576
rect 10321 2567 10379 2573
rect 10321 2533 10333 2567
rect 10367 2564 10379 2567
rect 11624 2564 11652 2595
rect 11698 2592 11704 2644
rect 11756 2632 11762 2644
rect 11977 2635 12035 2641
rect 11977 2632 11989 2635
rect 11756 2604 11989 2632
rect 11756 2592 11762 2604
rect 11977 2601 11989 2604
rect 12023 2601 12035 2635
rect 11977 2595 12035 2601
rect 12069 2635 12127 2641
rect 12069 2601 12081 2635
rect 12115 2632 12127 2635
rect 12526 2632 12532 2644
rect 12115 2604 12532 2632
rect 12115 2601 12127 2604
rect 12069 2595 12127 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 13998 2632 14004 2644
rect 13959 2604 14004 2632
rect 13998 2592 14004 2604
rect 14056 2632 14062 2644
rect 14918 2632 14924 2644
rect 14056 2604 14924 2632
rect 14056 2592 14062 2604
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 16758 2632 16764 2644
rect 16719 2604 16764 2632
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 13446 2564 13452 2576
rect 10367 2536 11652 2564
rect 12636 2536 13452 2564
rect 10367 2533 10379 2536
rect 10321 2527 10379 2533
rect 8570 2496 8576 2508
rect 8021 2459 8079 2465
rect 8312 2468 8432 2496
rect 8531 2468 8576 2496
rect 4246 2428 4252 2440
rect 4207 2400 4252 2428
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 5350 2428 5356 2440
rect 5311 2400 5356 2428
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 4798 2360 4804 2372
rect 3620 2332 4804 2360
rect 4798 2320 4804 2332
rect 4856 2320 4862 2372
rect 4890 2320 4896 2372
rect 4948 2360 4954 2372
rect 5736 2360 5764 2391
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6273 2431 6331 2437
rect 6273 2428 6285 2431
rect 5868 2400 6285 2428
rect 5868 2388 5874 2400
rect 6273 2397 6285 2400
rect 6319 2397 6331 2431
rect 6273 2391 6331 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 8312 2428 8340 2468
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 9125 2499 9183 2505
rect 9125 2465 9137 2499
rect 9171 2496 9183 2499
rect 9171 2468 10548 2496
rect 9171 2465 9183 2468
rect 9125 2459 9183 2465
rect 8757 2431 8815 2437
rect 8757 2428 8769 2431
rect 7791 2400 8340 2428
rect 8404 2400 8769 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 4948 2332 5764 2360
rect 4948 2320 4954 2332
rect 7558 2320 7564 2372
rect 7616 2360 7622 2372
rect 8404 2360 8432 2400
rect 8757 2397 8769 2400
rect 8803 2397 8815 2431
rect 8757 2391 8815 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 7616 2332 8432 2360
rect 7616 2320 7622 2332
rect 8478 2320 8484 2372
rect 8536 2360 8542 2372
rect 9324 2360 9352 2391
rect 8536 2332 9352 2360
rect 10520 2360 10548 2468
rect 10870 2456 10876 2508
rect 10928 2496 10934 2508
rect 12636 2505 12664 2536
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 10928 2468 11161 2496
rect 10928 2456 10934 2468
rect 11149 2465 11161 2468
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2465 12679 2499
rect 13170 2496 13176 2508
rect 13131 2468 13176 2496
rect 12621 2459 12679 2465
rect 13170 2456 13176 2468
rect 13228 2456 13234 2508
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 15286 2496 15292 2508
rect 14415 2468 15292 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 16117 2499 16175 2505
rect 16117 2465 16129 2499
rect 16163 2465 16175 2499
rect 16776 2496 16804 2592
rect 16942 2524 16948 2576
rect 17000 2564 17006 2576
rect 17000 2536 17908 2564
rect 17000 2524 17006 2536
rect 17880 2505 17908 2536
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16776 2468 17141 2496
rect 16117 2459 16175 2465
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 17497 2499 17555 2505
rect 17497 2465 17509 2499
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 17865 2499 17923 2505
rect 17865 2465 17877 2499
rect 17911 2496 17923 2499
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 17911 2468 18337 2496
rect 17911 2465 17923 2468
rect 17865 2459 17923 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 11054 2428 11060 2440
rect 10643 2400 11060 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11330 2388 11336 2440
rect 11388 2428 11394 2440
rect 11425 2431 11483 2437
rect 11425 2428 11437 2431
rect 11388 2400 11437 2428
rect 11388 2388 11394 2400
rect 11425 2397 11437 2400
rect 11471 2428 11483 2431
rect 12161 2431 12219 2437
rect 12161 2428 12173 2431
rect 11471 2400 12173 2428
rect 11471 2397 11483 2400
rect 11425 2391 11483 2397
rect 12161 2397 12173 2400
rect 12207 2397 12219 2431
rect 12161 2391 12219 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12308 2400 12817 2428
rect 12308 2388 12314 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 13136 2400 13369 2428
rect 13136 2388 13142 2400
rect 13357 2397 13369 2400
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 13964 2400 14565 2428
rect 13964 2388 13970 2400
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 16132 2428 16160 2459
rect 16666 2428 16672 2440
rect 16132 2400 16672 2428
rect 14553 2391 14611 2397
rect 16666 2388 16672 2400
rect 16724 2428 16730 2440
rect 16850 2428 16856 2440
rect 16724 2400 16856 2428
rect 16724 2388 16730 2400
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 17218 2428 17224 2440
rect 17083 2400 17224 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 17218 2388 17224 2400
rect 17276 2428 17282 2440
rect 17512 2428 17540 2459
rect 17276 2400 17540 2428
rect 17276 2388 17282 2400
rect 11146 2360 11152 2372
rect 10520 2332 11152 2360
rect 8536 2320 8542 2332
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 3418 2292 3424 2304
rect 3379 2264 3424 2292
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 3786 2292 3792 2304
rect 3747 2264 3792 2292
rect 3786 2252 3792 2264
rect 3844 2252 3850 2304
rect 4816 2292 4844 2320
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 4816 2264 6653 2292
rect 6641 2261 6653 2264
rect 6687 2292 6699 2295
rect 7466 2292 7472 2304
rect 6687 2264 7472 2292
rect 6687 2261 6699 2264
rect 6641 2255 6699 2261
rect 7466 2252 7472 2264
rect 7524 2252 7530 2304
rect 9861 2295 9919 2301
rect 9861 2261 9873 2295
rect 9907 2292 9919 2295
rect 10870 2292 10876 2304
rect 9907 2264 10876 2292
rect 9907 2261 9919 2264
rect 9861 2255 9919 2261
rect 10870 2252 10876 2264
rect 10928 2252 10934 2304
rect 11422 2252 11428 2304
rect 11480 2292 11486 2304
rect 13725 2295 13783 2301
rect 13725 2292 13737 2295
rect 11480 2264 13737 2292
rect 11480 2252 11486 2264
rect 13725 2261 13737 2264
rect 13771 2261 13783 2295
rect 16298 2292 16304 2304
rect 16259 2264 16304 2292
rect 13725 2255 13783 2261
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 17310 2292 17316 2304
rect 17271 2264 17316 2292
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 17678 2292 17684 2304
rect 17639 2264 17684 2292
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 18049 2295 18107 2301
rect 18049 2292 18061 2295
rect 17920 2264 18061 2292
rect 17920 2252 17926 2264
rect 18049 2261 18061 2264
rect 18095 2261 18107 2295
rect 18049 2255 18107 2261
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 382 2048 388 2100
rect 440 2088 446 2100
rect 16298 2088 16304 2100
rect 440 2060 16304 2088
rect 440 2048 446 2060
rect 16298 2048 16304 2060
rect 16356 2048 16362 2100
<< via1 >>
rect 3424 15716 3476 15768
rect 6644 15716 6696 15768
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 13268 14560 13320 14612
rect 18052 14560 18104 14612
rect 12164 14492 12216 14544
rect 14372 14492 14424 14544
rect 18788 14492 18840 14544
rect 5908 14424 5960 14476
rect 4068 14356 4120 14408
rect 11428 14424 11480 14476
rect 15292 14356 15344 14408
rect 3792 14288 3844 14340
rect 8944 14288 8996 14340
rect 3332 14220 3384 14272
rect 13268 14220 13320 14272
rect 13360 14220 13412 14272
rect 16212 14220 16264 14272
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 5908 14059 5960 14068
rect 5908 14025 5917 14059
rect 5917 14025 5951 14059
rect 5951 14025 5960 14059
rect 5908 14016 5960 14025
rect 6736 14016 6788 14068
rect 16580 14016 16632 14068
rect 8208 13948 8260 14000
rect 14740 13948 14792 14000
rect 16028 13948 16080 14000
rect 6000 13880 6052 13932
rect 14372 13880 14424 13932
rect 16856 13923 16908 13932
rect 7196 13812 7248 13864
rect 7748 13812 7800 13864
rect 12716 13812 12768 13864
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 5540 13744 5592 13796
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 18052 13855 18104 13864
rect 16028 13787 16080 13796
rect 16028 13753 16037 13787
rect 16037 13753 16071 13787
rect 16071 13753 16080 13787
rect 16028 13744 16080 13753
rect 6092 13676 6144 13728
rect 6368 13719 6420 13728
rect 6368 13685 6377 13719
rect 6377 13685 6411 13719
rect 6411 13685 6420 13719
rect 6368 13676 6420 13685
rect 8392 13676 8444 13728
rect 10232 13676 10284 13728
rect 13636 13676 13688 13728
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 17592 13719 17644 13728
rect 17592 13685 17601 13719
rect 17601 13685 17635 13719
rect 17635 13685 17644 13719
rect 17592 13676 17644 13685
rect 18512 13676 18564 13728
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 8208 13515 8260 13524
rect 8208 13481 8217 13515
rect 8217 13481 8251 13515
rect 8251 13481 8260 13515
rect 8208 13472 8260 13481
rect 11704 13472 11756 13524
rect 13636 13472 13688 13524
rect 5724 13336 5776 13388
rect 4344 13268 4396 13320
rect 6828 13336 6880 13388
rect 8668 13404 8720 13456
rect 13084 13404 13136 13456
rect 13176 13404 13228 13456
rect 16948 13404 17000 13456
rect 8116 13379 8168 13388
rect 8116 13345 8125 13379
rect 8125 13345 8159 13379
rect 8159 13345 8168 13379
rect 8116 13336 8168 13345
rect 10784 13336 10836 13388
rect 13820 13336 13872 13388
rect 6736 13268 6788 13320
rect 8576 13268 8628 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 14556 13311 14608 13320
rect 1124 13132 1176 13184
rect 12716 13200 12768 13252
rect 6000 13175 6052 13184
rect 6000 13141 6009 13175
rect 6009 13141 6043 13175
rect 6043 13141 6052 13175
rect 6000 13132 6052 13141
rect 6828 13132 6880 13184
rect 9312 13132 9364 13184
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 14464 13132 14516 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 3700 12928 3752 12980
rect 5540 12928 5592 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 6368 12928 6420 12980
rect 13360 12928 13412 12980
rect 13728 12928 13780 12980
rect 13912 12860 13964 12912
rect 3792 12724 3844 12776
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 4344 12724 4396 12733
rect 6184 12656 6236 12708
rect 6736 12656 6788 12708
rect 7288 12724 7340 12776
rect 7564 12724 7616 12776
rect 7380 12656 7432 12708
rect 6000 12588 6052 12640
rect 7472 12588 7524 12640
rect 7656 12631 7708 12640
rect 7656 12597 7665 12631
rect 7665 12597 7699 12631
rect 7699 12597 7708 12631
rect 7656 12588 7708 12597
rect 13820 12792 13872 12844
rect 14188 12792 14240 12844
rect 16948 12971 17000 12980
rect 16948 12937 16957 12971
rect 16957 12937 16991 12971
rect 16991 12937 17000 12971
rect 16948 12928 17000 12937
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 8392 12724 8444 12776
rect 14372 12724 14424 12776
rect 15016 12724 15068 12776
rect 14924 12656 14976 12708
rect 17684 12835 17736 12844
rect 17684 12801 17693 12835
rect 17693 12801 17727 12835
rect 17727 12801 17736 12835
rect 17684 12792 17736 12801
rect 16304 12656 16356 12708
rect 14004 12631 14056 12640
rect 14004 12597 14013 12631
rect 14013 12597 14047 12631
rect 14047 12597 14056 12631
rect 14004 12588 14056 12597
rect 14096 12631 14148 12640
rect 14096 12597 14105 12631
rect 14105 12597 14139 12631
rect 14139 12597 14148 12631
rect 15936 12631 15988 12640
rect 14096 12588 14148 12597
rect 15936 12597 15945 12631
rect 15945 12597 15979 12631
rect 15979 12597 15988 12631
rect 15936 12588 15988 12597
rect 16120 12631 16172 12640
rect 16120 12597 16129 12631
rect 16129 12597 16163 12631
rect 16163 12597 16172 12631
rect 16120 12588 16172 12597
rect 17132 12631 17184 12640
rect 17132 12597 17141 12631
rect 17141 12597 17175 12631
rect 17175 12597 17184 12631
rect 17132 12588 17184 12597
rect 17408 12588 17460 12640
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 6000 12384 6052 12436
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 3976 12316 4028 12368
rect 5908 12316 5960 12368
rect 6000 12248 6052 12300
rect 6460 12316 6512 12368
rect 9680 12384 9732 12436
rect 13176 12384 13228 12436
rect 14096 12384 14148 12436
rect 14372 12384 14424 12436
rect 16120 12384 16172 12436
rect 16212 12384 16264 12436
rect 16764 12384 16816 12436
rect 8208 12359 8260 12368
rect 8208 12325 8217 12359
rect 8217 12325 8251 12359
rect 8251 12325 8260 12359
rect 8208 12316 8260 12325
rect 1492 12180 1544 12232
rect 2780 12180 2832 12232
rect 3792 12180 3844 12232
rect 5540 12180 5592 12232
rect 5908 12180 5960 12232
rect 6736 12248 6788 12300
rect 6920 12291 6972 12300
rect 6920 12257 6929 12291
rect 6929 12257 6963 12291
rect 6963 12257 6972 12291
rect 6920 12248 6972 12257
rect 6184 12180 6236 12232
rect 9036 12248 9088 12300
rect 9312 12316 9364 12368
rect 12348 12316 12400 12368
rect 14188 12316 14240 12368
rect 10600 12291 10652 12300
rect 10600 12257 10609 12291
rect 10609 12257 10643 12291
rect 10643 12257 10652 12291
rect 10600 12248 10652 12257
rect 7380 12180 7432 12232
rect 7656 12180 7708 12232
rect 8392 12180 8444 12232
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 9588 12180 9640 12232
rect 9680 12180 9732 12232
rect 10968 12180 11020 12232
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12716 12180 12768 12189
rect 14372 12248 14424 12300
rect 15016 12248 15068 12300
rect 2136 12044 2188 12096
rect 4252 12044 4304 12096
rect 4712 12044 4764 12096
rect 5448 12087 5500 12096
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 9036 12044 9088 12096
rect 10232 12087 10284 12096
rect 10232 12053 10241 12087
rect 10241 12053 10275 12087
rect 10275 12053 10284 12087
rect 10232 12044 10284 12053
rect 10600 12044 10652 12096
rect 12256 12044 12308 12096
rect 13820 12112 13872 12164
rect 14464 12044 14516 12096
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 15200 12180 15252 12232
rect 16672 12316 16724 12368
rect 17684 12248 17736 12300
rect 18144 12291 18196 12300
rect 18144 12257 18153 12291
rect 18153 12257 18187 12291
rect 18187 12257 18196 12291
rect 18144 12248 18196 12257
rect 17776 12180 17828 12232
rect 15384 12155 15436 12164
rect 15384 12121 15393 12155
rect 15393 12121 15427 12155
rect 15427 12121 15436 12155
rect 15384 12112 15436 12121
rect 17684 12112 17736 12164
rect 14832 12044 14884 12096
rect 16120 12044 16172 12096
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 3608 11883 3660 11892
rect 3608 11849 3617 11883
rect 3617 11849 3651 11883
rect 3651 11849 3660 11883
rect 3608 11840 3660 11849
rect 6736 11840 6788 11892
rect 9220 11840 9272 11892
rect 9312 11840 9364 11892
rect 12532 11840 12584 11892
rect 5356 11772 5408 11824
rect 7564 11772 7616 11824
rect 10324 11815 10376 11824
rect 2412 11704 2464 11756
rect 2688 11636 2740 11688
rect 3884 11636 3936 11688
rect 4620 11636 4672 11688
rect 5448 11636 5500 11688
rect 5540 11636 5592 11688
rect 1584 11568 1636 11620
rect 1400 11543 1452 11552
rect 1400 11509 1409 11543
rect 1409 11509 1443 11543
rect 1443 11509 1452 11543
rect 1400 11500 1452 11509
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 1768 11500 1820 11509
rect 2780 11568 2832 11620
rect 5816 11568 5868 11620
rect 6920 11568 6972 11620
rect 7564 11568 7616 11620
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 3792 11500 3844 11552
rect 5632 11500 5684 11552
rect 6460 11500 6512 11552
rect 7472 11500 7524 11552
rect 10324 11781 10333 11815
rect 10333 11781 10367 11815
rect 10367 11781 10376 11815
rect 10324 11772 10376 11781
rect 10692 11772 10744 11824
rect 14004 11840 14056 11892
rect 15200 11883 15252 11892
rect 15200 11849 15209 11883
rect 15209 11849 15243 11883
rect 15243 11849 15252 11883
rect 15200 11840 15252 11849
rect 16304 11840 16356 11892
rect 8392 11704 8444 11756
rect 7932 11636 7984 11688
rect 10600 11704 10652 11756
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 11060 11704 11112 11756
rect 10232 11636 10284 11688
rect 14372 11772 14424 11824
rect 17132 11840 17184 11892
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 18144 11840 18196 11892
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 13176 11704 13228 11756
rect 14740 11747 14792 11756
rect 14740 11713 14749 11747
rect 14749 11713 14783 11747
rect 14783 11713 14792 11747
rect 14740 11704 14792 11713
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 16212 11704 16264 11756
rect 13544 11636 13596 11688
rect 14556 11636 14608 11688
rect 16120 11636 16172 11688
rect 9220 11611 9272 11620
rect 9220 11577 9254 11611
rect 9254 11577 9272 11611
rect 9220 11568 9272 11577
rect 10140 11500 10192 11552
rect 14004 11568 14056 11620
rect 10600 11500 10652 11552
rect 11060 11500 11112 11552
rect 11244 11500 11296 11552
rect 13268 11500 13320 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 16580 11772 16632 11824
rect 16672 11747 16724 11756
rect 16672 11713 16681 11747
rect 16681 11713 16715 11747
rect 16715 11713 16724 11747
rect 16672 11704 16724 11713
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 16948 11568 17000 11620
rect 16764 11500 16816 11552
rect 17224 11543 17276 11552
rect 17224 11509 17233 11543
rect 17233 11509 17267 11543
rect 17267 11509 17276 11543
rect 17224 11500 17276 11509
rect 17316 11543 17368 11552
rect 17316 11509 17325 11543
rect 17325 11509 17359 11543
rect 17359 11509 17368 11543
rect 17316 11500 17368 11509
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 2688 11296 2740 11348
rect 2412 11271 2464 11280
rect 2412 11237 2446 11271
rect 2446 11237 2464 11271
rect 2412 11228 2464 11237
rect 3608 11228 3660 11280
rect 1952 11160 2004 11212
rect 2964 11160 3016 11212
rect 5540 11160 5592 11212
rect 5724 11203 5776 11212
rect 5724 11169 5758 11203
rect 5758 11169 5776 11203
rect 5724 11160 5776 11169
rect 6184 11160 6236 11212
rect 9220 11296 9272 11348
rect 9312 11296 9364 11348
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 11152 11339 11204 11348
rect 11152 11305 11161 11339
rect 11161 11305 11195 11339
rect 11195 11305 11204 11339
rect 13268 11339 13320 11348
rect 11152 11296 11204 11305
rect 13268 11305 13277 11339
rect 13277 11305 13311 11339
rect 13311 11305 13320 11339
rect 13268 11296 13320 11305
rect 13820 11296 13872 11348
rect 14004 11296 14056 11348
rect 14648 11296 14700 11348
rect 15016 11296 15068 11348
rect 16672 11296 16724 11348
rect 17224 11296 17276 11348
rect 18420 11339 18472 11348
rect 18420 11305 18429 11339
rect 18429 11305 18463 11339
rect 18463 11305 18472 11339
rect 18420 11296 18472 11305
rect 8208 11228 8260 11280
rect 10692 11228 10744 11280
rect 10968 11228 11020 11280
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 7840 11160 7892 11212
rect 8300 11160 8352 11212
rect 10508 11203 10560 11212
rect 1492 11092 1544 11144
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 3608 11092 3660 11144
rect 4344 11092 4396 11144
rect 5356 11092 5408 11144
rect 7012 11092 7064 11144
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 8760 11092 8812 11144
rect 9588 11092 9640 11144
rect 3884 11024 3936 11076
rect 5264 11067 5316 11076
rect 5264 11033 5273 11067
rect 5273 11033 5307 11067
rect 5307 11033 5316 11067
rect 5264 11024 5316 11033
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 9404 11024 9456 11076
rect 10508 11169 10517 11203
rect 10517 11169 10551 11203
rect 10551 11169 10560 11203
rect 10508 11160 10560 11169
rect 11152 11160 11204 11212
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 12808 11228 12860 11280
rect 12900 11228 12952 11280
rect 11336 11092 11388 11144
rect 12808 11092 12860 11144
rect 13176 11024 13228 11076
rect 3700 10956 3752 11008
rect 4436 10956 4488 11008
rect 4528 10999 4580 11008
rect 4528 10965 4537 10999
rect 4537 10965 4571 10999
rect 4571 10965 4580 10999
rect 4896 10999 4948 11008
rect 4528 10956 4580 10965
rect 4896 10965 4905 10999
rect 4905 10965 4939 10999
rect 4939 10965 4948 10999
rect 4896 10956 4948 10965
rect 5080 10956 5132 11008
rect 13268 10956 13320 11008
rect 13912 11160 13964 11212
rect 15108 11203 15160 11212
rect 15108 11169 15117 11203
rect 15117 11169 15151 11203
rect 15151 11169 15160 11203
rect 15108 11160 15160 11169
rect 15568 11160 15620 11212
rect 16948 11203 17000 11212
rect 16948 11169 16957 11203
rect 16957 11169 16991 11203
rect 16991 11169 17000 11203
rect 16948 11160 17000 11169
rect 17868 11203 17920 11212
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 14004 11092 14056 11144
rect 15016 11092 15068 11144
rect 17776 11092 17828 11144
rect 14832 11024 14884 11076
rect 13820 10956 13872 11008
rect 16764 10956 16816 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 1768 10752 1820 10804
rect 3424 10752 3476 10804
rect 5080 10752 5132 10804
rect 5540 10752 5592 10804
rect 6184 10795 6236 10804
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2964 10684 3016 10736
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 7012 10752 7064 10804
rect 7472 10752 7524 10804
rect 8852 10795 8904 10804
rect 8852 10761 8861 10795
rect 8861 10761 8895 10795
rect 8895 10761 8904 10795
rect 8852 10752 8904 10761
rect 9128 10752 9180 10804
rect 17500 10795 17552 10804
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 4620 10659 4672 10668
rect 4620 10625 4629 10659
rect 4629 10625 4663 10659
rect 4663 10625 4672 10659
rect 4620 10616 4672 10625
rect 5816 10616 5868 10668
rect 11336 10684 11388 10736
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 7564 10616 7616 10668
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 9404 10659 9456 10668
rect 9404 10625 9413 10659
rect 9413 10625 9447 10659
rect 9447 10625 9456 10659
rect 9404 10616 9456 10625
rect 1400 10548 1452 10600
rect 3056 10548 3108 10600
rect 4712 10548 4764 10600
rect 6460 10591 6512 10600
rect 2964 10480 3016 10532
rect 1676 10412 1728 10464
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 3424 10412 3476 10464
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 4804 10412 4856 10464
rect 6460 10557 6469 10591
rect 6469 10557 6503 10591
rect 6503 10557 6512 10591
rect 6460 10548 6512 10557
rect 6920 10548 6972 10600
rect 8852 10548 8904 10600
rect 5080 10523 5132 10532
rect 5080 10489 5114 10523
rect 5114 10489 5132 10523
rect 5080 10480 5132 10489
rect 5172 10480 5224 10532
rect 9772 10591 9824 10600
rect 9772 10557 9781 10591
rect 9781 10557 9815 10591
rect 9815 10557 9824 10591
rect 9772 10548 9824 10557
rect 9680 10480 9732 10532
rect 10324 10480 10376 10532
rect 10600 10480 10652 10532
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 7380 10412 7432 10464
rect 7840 10412 7892 10464
rect 9312 10412 9364 10464
rect 9496 10412 9548 10464
rect 11336 10548 11388 10600
rect 11612 10548 11664 10600
rect 11888 10591 11940 10600
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 17684 10684 17736 10736
rect 18972 10684 19024 10736
rect 13912 10659 13964 10668
rect 11888 10548 11940 10557
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 12164 10480 12216 10532
rect 13176 10548 13228 10600
rect 14280 10548 14332 10600
rect 15016 10548 15068 10600
rect 12624 10480 12676 10532
rect 12440 10412 12492 10464
rect 13728 10480 13780 10532
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 15568 10412 15620 10464
rect 16028 10455 16080 10464
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 16580 10480 16632 10532
rect 16672 10412 16724 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 2044 10208 2096 10260
rect 4436 10208 4488 10260
rect 5172 10208 5224 10260
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 7288 10208 7340 10260
rect 7472 10208 7524 10260
rect 10324 10251 10376 10260
rect 2688 10140 2740 10192
rect 4344 10140 4396 10192
rect 2596 10072 2648 10124
rect 3424 10072 3476 10124
rect 6184 10140 6236 10192
rect 7380 10140 7432 10192
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 4160 10004 4212 10056
rect 4436 9936 4488 9988
rect 3424 9868 3476 9920
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 5540 10047 5592 10056
rect 4712 10004 4764 10013
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 6920 10072 6972 10124
rect 7656 10072 7708 10124
rect 7932 10115 7984 10124
rect 7932 10081 7941 10115
rect 7941 10081 7975 10115
rect 7975 10081 7984 10115
rect 7932 10072 7984 10081
rect 9496 10140 9548 10192
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 11520 10208 11572 10260
rect 12072 10208 12124 10260
rect 15108 10208 15160 10260
rect 10876 10140 10928 10192
rect 9404 10115 9456 10124
rect 7380 10047 7432 10056
rect 5080 9936 5132 9988
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 7012 9936 7064 9988
rect 9404 10081 9413 10115
rect 9413 10081 9447 10115
rect 9447 10081 9456 10115
rect 9404 10072 9456 10081
rect 9220 10004 9272 10056
rect 10416 10072 10468 10124
rect 10232 10004 10284 10056
rect 10692 9936 10744 9988
rect 13820 10140 13872 10192
rect 13912 10140 13964 10192
rect 16028 10140 16080 10192
rect 17316 10251 17368 10260
rect 17316 10217 17325 10251
rect 17325 10217 17359 10251
rect 17359 10217 17368 10251
rect 17316 10208 17368 10217
rect 17684 10208 17736 10260
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 11244 10004 11296 10056
rect 12072 10004 12124 10056
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 12808 10072 12860 10124
rect 14556 10072 14608 10124
rect 15660 10072 15712 10124
rect 12992 10004 13044 10056
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 16672 10140 16724 10192
rect 17500 10140 17552 10192
rect 17868 10208 17920 10260
rect 17132 10072 17184 10124
rect 17684 10115 17736 10124
rect 17684 10081 17693 10115
rect 17693 10081 17727 10115
rect 17727 10081 17736 10115
rect 17684 10072 17736 10081
rect 16672 10047 16724 10056
rect 11888 9936 11940 9988
rect 12900 9936 12952 9988
rect 16672 10013 16681 10047
rect 16681 10013 16715 10047
rect 16715 10013 16724 10047
rect 16672 10004 16724 10013
rect 5356 9868 5408 9920
rect 6092 9868 6144 9920
rect 6920 9868 6972 9920
rect 7472 9868 7524 9920
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 9404 9868 9456 9920
rect 10416 9868 10468 9920
rect 12256 9868 12308 9920
rect 15016 9936 15068 9988
rect 16580 9936 16632 9988
rect 17776 10004 17828 10056
rect 17132 9979 17184 9988
rect 17132 9945 17141 9979
rect 17141 9945 17175 9979
rect 17175 9945 17184 9979
rect 17132 9936 17184 9945
rect 14740 9911 14792 9920
rect 14740 9877 14749 9911
rect 14749 9877 14783 9911
rect 14783 9877 14792 9911
rect 14740 9868 14792 9877
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 16304 9868 16356 9920
rect 18052 9868 18104 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 4344 9664 4396 9716
rect 4436 9596 4488 9648
rect 5540 9596 5592 9648
rect 1400 9528 1452 9580
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 4712 9528 4764 9580
rect 6184 9528 6236 9580
rect 7012 9528 7064 9580
rect 8116 9664 8168 9716
rect 8852 9664 8904 9716
rect 11336 9664 11388 9716
rect 12256 9664 12308 9716
rect 2044 9460 2096 9512
rect 4436 9460 4488 9512
rect 4804 9460 4856 9512
rect 3700 9435 3752 9444
rect 3056 9324 3108 9376
rect 3700 9401 3712 9435
rect 3712 9401 3752 9435
rect 3700 9392 3752 9401
rect 5080 9392 5132 9444
rect 7380 9392 7432 9444
rect 7748 9392 7800 9444
rect 8208 9596 8260 9648
rect 8484 9596 8536 9648
rect 11428 9639 11480 9648
rect 8024 9571 8076 9580
rect 8024 9537 8033 9571
rect 8033 9537 8067 9571
rect 8067 9537 8076 9571
rect 8024 9528 8076 9537
rect 9496 9528 9548 9580
rect 9680 9528 9732 9580
rect 11428 9605 11437 9639
rect 11437 9605 11471 9639
rect 11471 9605 11480 9639
rect 11428 9596 11480 9605
rect 11980 9596 12032 9648
rect 14004 9596 14056 9648
rect 14188 9596 14240 9648
rect 15660 9664 15712 9716
rect 16672 9707 16724 9716
rect 16672 9673 16681 9707
rect 16681 9673 16715 9707
rect 16715 9673 16724 9707
rect 16672 9664 16724 9673
rect 15752 9596 15804 9648
rect 12072 9571 12124 9580
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 9772 9460 9824 9512
rect 12072 9537 12081 9571
rect 12081 9537 12115 9571
rect 12115 9537 12124 9571
rect 12072 9528 12124 9537
rect 16580 9528 16632 9580
rect 17224 9571 17276 9580
rect 17224 9537 17233 9571
rect 17233 9537 17267 9571
rect 17267 9537 17276 9571
rect 17224 9528 17276 9537
rect 9680 9392 9732 9444
rect 4160 9324 4212 9376
rect 4620 9324 4672 9376
rect 6092 9324 6144 9376
rect 6276 9367 6328 9376
rect 6276 9333 6285 9367
rect 6285 9333 6319 9367
rect 6319 9333 6328 9367
rect 6276 9324 6328 9333
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 9220 9324 9272 9376
rect 9772 9324 9824 9376
rect 11612 9460 11664 9512
rect 10876 9392 10928 9444
rect 10968 9392 11020 9444
rect 12164 9460 12216 9512
rect 12716 9503 12768 9512
rect 12716 9469 12750 9503
rect 12750 9469 12768 9503
rect 11888 9435 11940 9444
rect 11888 9401 11897 9435
rect 11897 9401 11931 9435
rect 11931 9401 11940 9435
rect 11888 9392 11940 9401
rect 12716 9460 12768 9469
rect 14280 9460 14332 9512
rect 14740 9460 14792 9512
rect 15200 9460 15252 9512
rect 18144 9460 18196 9512
rect 12900 9392 12952 9444
rect 10048 9324 10100 9376
rect 10324 9324 10376 9376
rect 10600 9324 10652 9376
rect 10692 9324 10744 9376
rect 11980 9367 12032 9376
rect 11980 9333 11989 9367
rect 11989 9333 12023 9367
rect 12023 9333 12032 9367
rect 11980 9324 12032 9333
rect 12348 9324 12400 9376
rect 15108 9324 15160 9376
rect 15752 9367 15804 9376
rect 15752 9333 15761 9367
rect 15761 9333 15795 9367
rect 15795 9333 15804 9367
rect 15752 9324 15804 9333
rect 16672 9324 16724 9376
rect 17132 9367 17184 9376
rect 17132 9333 17141 9367
rect 17141 9333 17175 9367
rect 17175 9333 17184 9367
rect 17132 9324 17184 9333
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 2596 9163 2648 9172
rect 2596 9129 2605 9163
rect 2605 9129 2639 9163
rect 2639 9129 2648 9163
rect 2596 9120 2648 9129
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 3148 9120 3200 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 4160 9163 4212 9172
rect 3424 9120 3476 9129
rect 4160 9129 4169 9163
rect 4169 9129 4203 9163
rect 4203 9129 4212 9163
rect 4160 9120 4212 9129
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 4896 9163 4948 9172
rect 1952 8984 2004 9036
rect 2688 9052 2740 9104
rect 2872 8984 2924 9036
rect 3424 8984 3476 9036
rect 2780 8916 2832 8968
rect 4896 9129 4905 9163
rect 4905 9129 4939 9163
rect 4939 9129 4948 9163
rect 4896 9120 4948 9129
rect 5172 9120 5224 9172
rect 4804 9052 4856 9104
rect 6000 8984 6052 9036
rect 7380 9052 7432 9104
rect 8208 9120 8260 9172
rect 9036 9163 9088 9172
rect 9036 9129 9045 9163
rect 9045 9129 9079 9163
rect 9079 9129 9088 9163
rect 9036 9120 9088 9129
rect 11796 9120 11848 9172
rect 11980 9163 12032 9172
rect 11980 9129 11989 9163
rect 11989 9129 12023 9163
rect 12023 9129 12032 9163
rect 11980 9120 12032 9129
rect 12348 9163 12400 9172
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 9312 9052 9364 9104
rect 10048 9052 10100 9104
rect 12532 9052 12584 9104
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 2136 8823 2188 8832
rect 2136 8789 2145 8823
rect 2145 8789 2179 8823
rect 2179 8789 2188 8823
rect 2136 8780 2188 8789
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 7472 8984 7524 9036
rect 7932 8984 7984 9036
rect 8392 8984 8444 9036
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 9312 8916 9364 8968
rect 11152 8984 11204 9036
rect 7196 8780 7248 8832
rect 7564 8780 7616 8832
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 11060 8916 11112 8968
rect 10692 8848 10744 8900
rect 12532 8916 12584 8968
rect 13728 9052 13780 9104
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 13636 8984 13688 9036
rect 15200 9120 15252 9172
rect 15384 9120 15436 9172
rect 16028 9120 16080 9172
rect 16396 9120 16448 9172
rect 17868 9120 17920 9172
rect 14280 9052 14332 9104
rect 14648 8984 14700 9036
rect 16120 9052 16172 9104
rect 17224 9052 17276 9104
rect 12716 8916 12768 8968
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 16396 8984 16448 9036
rect 16672 8984 16724 9036
rect 14464 8848 14516 8900
rect 14740 8848 14792 8900
rect 15476 8916 15528 8968
rect 15568 8916 15620 8968
rect 15384 8848 15436 8900
rect 10600 8780 10652 8832
rect 10876 8780 10928 8832
rect 11796 8780 11848 8832
rect 11888 8780 11940 8832
rect 13360 8780 13412 8832
rect 13636 8823 13688 8832
rect 13636 8789 13645 8823
rect 13645 8789 13679 8823
rect 13679 8789 13688 8823
rect 13636 8780 13688 8789
rect 13820 8780 13872 8832
rect 14188 8780 14240 8832
rect 14556 8780 14608 8832
rect 15292 8823 15344 8832
rect 15292 8789 15301 8823
rect 15301 8789 15335 8823
rect 15335 8789 15344 8823
rect 15292 8780 15344 8789
rect 15476 8780 15528 8832
rect 16580 8780 16632 8832
rect 18328 8780 18380 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 2596 8576 2648 8628
rect 2964 8619 3016 8628
rect 2964 8585 2973 8619
rect 2973 8585 3007 8619
rect 3007 8585 3016 8619
rect 2964 8576 3016 8585
rect 4436 8576 4488 8628
rect 5356 8576 5408 8628
rect 6276 8576 6328 8628
rect 3424 8508 3476 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 5724 8508 5776 8560
rect 6460 8551 6512 8560
rect 6460 8517 6469 8551
rect 6469 8517 6503 8551
rect 6503 8517 6512 8551
rect 6460 8508 6512 8517
rect 5632 8440 5684 8492
rect 2780 8372 2832 8424
rect 2964 8372 3016 8424
rect 3976 8415 4028 8424
rect 3424 8304 3476 8356
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 5816 8372 5868 8424
rect 6460 8304 6512 8356
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 7472 8440 7524 8492
rect 8760 8440 8812 8492
rect 10140 8440 10192 8492
rect 7196 8372 7248 8424
rect 12624 8576 12676 8628
rect 17224 8619 17276 8628
rect 17224 8585 17233 8619
rect 17233 8585 17267 8619
rect 17267 8585 17276 8619
rect 17224 8576 17276 8585
rect 11796 8508 11848 8560
rect 13176 8508 13228 8560
rect 10508 8440 10560 8492
rect 11060 8440 11112 8492
rect 11520 8440 11572 8492
rect 11980 8440 12032 8492
rect 12256 8440 12308 8492
rect 14188 8508 14240 8560
rect 13912 8483 13964 8492
rect 6736 8304 6788 8356
rect 7472 8347 7524 8356
rect 7472 8313 7481 8347
rect 7481 8313 7515 8347
rect 7515 8313 7524 8347
rect 7472 8304 7524 8313
rect 8668 8304 8720 8356
rect 9036 8347 9088 8356
rect 9036 8313 9045 8347
rect 9045 8313 9079 8347
rect 9079 8313 9088 8347
rect 9036 8304 9088 8313
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 15660 8508 15712 8560
rect 17868 8508 17920 8560
rect 15108 8440 15160 8492
rect 15568 8440 15620 8492
rect 10692 8304 10744 8356
rect 2872 8236 2924 8288
rect 3148 8279 3200 8288
rect 3148 8245 3157 8279
rect 3157 8245 3191 8279
rect 3191 8245 3200 8279
rect 3148 8236 3200 8245
rect 3700 8236 3752 8288
rect 4252 8236 4304 8288
rect 6000 8279 6052 8288
rect 6000 8245 6009 8279
rect 6009 8245 6043 8279
rect 6043 8245 6052 8279
rect 6000 8236 6052 8245
rect 6276 8279 6328 8288
rect 6276 8245 6285 8279
rect 6285 8245 6319 8279
rect 6319 8245 6328 8279
rect 6276 8236 6328 8245
rect 8392 8236 8444 8288
rect 8944 8279 8996 8288
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 9220 8236 9272 8288
rect 11428 8304 11480 8356
rect 12532 8304 12584 8356
rect 11244 8236 11296 8288
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 14188 8304 14240 8356
rect 14924 8304 14976 8356
rect 15384 8347 15436 8356
rect 15384 8313 15393 8347
rect 15393 8313 15427 8347
rect 15427 8313 15436 8347
rect 16396 8372 16448 8424
rect 17684 8372 17736 8424
rect 15384 8304 15436 8313
rect 16672 8304 16724 8356
rect 14372 8236 14424 8288
rect 14464 8279 14516 8288
rect 14464 8245 14473 8279
rect 14473 8245 14507 8279
rect 14507 8245 14516 8279
rect 14464 8236 14516 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 2136 8032 2188 8084
rect 3148 8032 3200 8084
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 4344 8032 4396 8084
rect 4804 8032 4856 8084
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 9680 8075 9732 8084
rect 9680 8041 9689 8075
rect 9689 8041 9723 8075
rect 9723 8041 9732 8075
rect 9680 8032 9732 8041
rect 10232 8032 10284 8084
rect 10508 8075 10560 8084
rect 10508 8041 10517 8075
rect 10517 8041 10551 8075
rect 10551 8041 10560 8075
rect 10508 8032 10560 8041
rect 10600 8032 10652 8084
rect 11428 8032 11480 8084
rect 12716 8075 12768 8084
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 5632 7964 5684 8016
rect 5816 7964 5868 8016
rect 4344 7896 4396 7948
rect 2872 7828 2924 7880
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 3516 7828 3568 7880
rect 3700 7828 3752 7880
rect 4436 7828 4488 7880
rect 3608 7760 3660 7812
rect 5540 7896 5592 7948
rect 6000 7871 6052 7880
rect 6000 7837 6009 7871
rect 6009 7837 6043 7871
rect 6043 7837 6052 7871
rect 6000 7828 6052 7837
rect 6644 7964 6696 8016
rect 6736 7964 6788 8016
rect 8300 7964 8352 8016
rect 7472 7896 7524 7948
rect 7656 7896 7708 7948
rect 8024 7896 8076 7948
rect 10508 7896 10560 7948
rect 11520 7964 11572 8016
rect 14924 7964 14976 8016
rect 11428 7896 11480 7948
rect 13360 7896 13412 7948
rect 13820 7896 13872 7948
rect 13912 7896 13964 7948
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 10416 7828 10468 7880
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 5264 7760 5316 7812
rect 1768 7735 1820 7744
rect 1768 7701 1777 7735
rect 1777 7701 1811 7735
rect 1811 7701 1820 7735
rect 1768 7692 1820 7701
rect 2136 7692 2188 7744
rect 3332 7692 3384 7744
rect 4804 7692 4856 7744
rect 6184 7692 6236 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 7012 7760 7064 7812
rect 10048 7760 10100 7812
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 8300 7692 8352 7744
rect 9220 7692 9272 7744
rect 9496 7692 9548 7744
rect 10968 7692 11020 7744
rect 11060 7692 11112 7744
rect 12348 7828 12400 7880
rect 16396 7896 16448 7948
rect 12808 7692 12860 7744
rect 14280 7692 14332 7744
rect 14556 7692 14608 7744
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 14924 7735 14976 7744
rect 14924 7701 14933 7735
rect 14933 7701 14967 7735
rect 14967 7701 14976 7735
rect 14924 7692 14976 7701
rect 18052 7803 18104 7812
rect 18052 7769 18061 7803
rect 18061 7769 18095 7803
rect 18095 7769 18104 7803
rect 18052 7760 18104 7769
rect 15568 7692 15620 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 5172 7488 5224 7540
rect 5816 7488 5868 7540
rect 1584 7420 1636 7472
rect 8024 7488 8076 7540
rect 11244 7488 11296 7540
rect 2412 7284 2464 7336
rect 3608 7352 3660 7404
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 6460 7395 6512 7404
rect 6460 7361 6469 7395
rect 6469 7361 6503 7395
rect 6503 7361 6512 7395
rect 6460 7352 6512 7361
rect 6552 7352 6604 7404
rect 11060 7420 11112 7472
rect 14188 7531 14240 7540
rect 14188 7497 14197 7531
rect 14197 7497 14231 7531
rect 14231 7497 14240 7531
rect 14188 7488 14240 7497
rect 14372 7488 14424 7540
rect 16488 7488 16540 7540
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 4252 7284 4304 7336
rect 6276 7284 6328 7336
rect 6368 7284 6420 7336
rect 7012 7284 7064 7336
rect 2872 7216 2924 7268
rect 3424 7216 3476 7268
rect 2780 7148 2832 7200
rect 3240 7191 3292 7200
rect 3240 7157 3249 7191
rect 3249 7157 3283 7191
rect 3283 7157 3292 7191
rect 3240 7148 3292 7157
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 4068 7148 4120 7200
rect 4804 7191 4856 7200
rect 4804 7157 4813 7191
rect 4813 7157 4847 7191
rect 4847 7157 4856 7191
rect 4804 7148 4856 7157
rect 5816 7216 5868 7268
rect 7656 7216 7708 7268
rect 10048 7352 10100 7404
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 12532 7420 12584 7472
rect 13452 7420 13504 7472
rect 13912 7395 13964 7404
rect 8944 7284 8996 7336
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 15016 7420 15068 7472
rect 18236 7463 18288 7472
rect 18236 7429 18245 7463
rect 18245 7429 18279 7463
rect 18279 7429 18288 7463
rect 18236 7420 18288 7429
rect 15108 7352 15160 7404
rect 15660 7352 15712 7404
rect 16396 7395 16448 7404
rect 16396 7361 16405 7395
rect 16405 7361 16439 7395
rect 16439 7361 16448 7395
rect 16396 7352 16448 7361
rect 11336 7284 11388 7336
rect 12808 7327 12860 7336
rect 11152 7216 11204 7268
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 15476 7327 15528 7336
rect 5632 7148 5684 7200
rect 8024 7191 8076 7200
rect 8024 7157 8033 7191
rect 8033 7157 8067 7191
rect 8067 7157 8076 7191
rect 8024 7148 8076 7157
rect 9496 7191 9548 7200
rect 9496 7157 9505 7191
rect 9505 7157 9539 7191
rect 9539 7157 9548 7191
rect 9496 7148 9548 7157
rect 10416 7148 10468 7200
rect 12348 7216 12400 7268
rect 13728 7259 13780 7268
rect 13728 7225 13737 7259
rect 13737 7225 13771 7259
rect 13771 7225 13780 7259
rect 13728 7216 13780 7225
rect 12164 7148 12216 7200
rect 12256 7148 12308 7200
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 13360 7148 13412 7157
rect 13636 7148 13688 7200
rect 15476 7293 15485 7327
rect 15485 7293 15519 7327
rect 15519 7293 15528 7327
rect 15476 7284 15528 7293
rect 16488 7284 16540 7336
rect 17960 7284 18012 7336
rect 14556 7191 14608 7200
rect 14556 7157 14565 7191
rect 14565 7157 14599 7191
rect 14599 7157 14608 7191
rect 14556 7148 14608 7157
rect 15384 7191 15436 7200
rect 15384 7157 15393 7191
rect 15393 7157 15427 7191
rect 15427 7157 15436 7191
rect 15384 7148 15436 7157
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 2872 6944 2924 6996
rect 3608 6944 3660 6996
rect 4620 6944 4672 6996
rect 4804 6944 4856 6996
rect 5908 6944 5960 6996
rect 6000 6944 6052 6996
rect 2136 6919 2188 6928
rect 2136 6885 2145 6919
rect 2145 6885 2179 6919
rect 2179 6885 2188 6919
rect 2136 6876 2188 6885
rect 1860 6808 1912 6860
rect 4344 6876 4396 6928
rect 4712 6876 4764 6928
rect 11244 6944 11296 6996
rect 11520 6987 11572 6996
rect 11520 6953 11529 6987
rect 11529 6953 11563 6987
rect 11563 6953 11572 6987
rect 11520 6944 11572 6953
rect 12072 6987 12124 6996
rect 12072 6953 12081 6987
rect 12081 6953 12115 6987
rect 12115 6953 12124 6987
rect 12072 6944 12124 6953
rect 11152 6876 11204 6928
rect 12164 6876 12216 6928
rect 2780 6851 2832 6860
rect 2780 6817 2814 6851
rect 2814 6817 2832 6851
rect 2780 6808 2832 6817
rect 4804 6808 4856 6860
rect 5080 6808 5132 6860
rect 2412 6740 2464 6792
rect 1768 6672 1820 6724
rect 4344 6672 4396 6724
rect 5540 6672 5592 6724
rect 6368 6808 6420 6860
rect 6828 6808 6880 6860
rect 7196 6851 7248 6860
rect 7196 6817 7230 6851
rect 7230 6817 7248 6851
rect 7196 6808 7248 6817
rect 9128 6851 9180 6860
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 9128 6808 9180 6817
rect 10232 6808 10284 6860
rect 11336 6808 11388 6860
rect 13268 6944 13320 6996
rect 13636 6944 13688 6996
rect 14096 6808 14148 6860
rect 14372 6876 14424 6928
rect 15384 6944 15436 6996
rect 16120 6944 16172 6996
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 6276 6740 6328 6792
rect 5724 6672 5776 6724
rect 2228 6604 2280 6656
rect 4528 6604 4580 6656
rect 5816 6604 5868 6656
rect 7932 6672 7984 6724
rect 10048 6740 10100 6792
rect 11152 6740 11204 6792
rect 9588 6672 9640 6724
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 9680 6604 9732 6656
rect 11520 6604 11572 6656
rect 12072 6604 12124 6656
rect 12164 6604 12216 6656
rect 12808 6604 12860 6656
rect 13084 6740 13136 6792
rect 14280 6740 14332 6792
rect 13820 6672 13872 6724
rect 14648 6740 14700 6792
rect 15016 6740 15068 6792
rect 14832 6715 14884 6724
rect 14832 6681 14841 6715
rect 14841 6681 14875 6715
rect 14875 6681 14884 6715
rect 14832 6672 14884 6681
rect 16948 6672 17000 6724
rect 13912 6604 13964 6656
rect 14280 6604 14332 6656
rect 14648 6604 14700 6656
rect 17500 6604 17552 6656
rect 18420 6715 18472 6724
rect 18420 6681 18429 6715
rect 18429 6681 18463 6715
rect 18463 6681 18472 6715
rect 18420 6672 18472 6681
rect 18052 6647 18104 6656
rect 18052 6613 18061 6647
rect 18061 6613 18095 6647
rect 18095 6613 18104 6647
rect 18052 6604 18104 6613
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 2872 6400 2924 6452
rect 3608 6443 3660 6452
rect 3608 6409 3617 6443
rect 3617 6409 3651 6443
rect 3651 6409 3660 6443
rect 3608 6400 3660 6409
rect 2964 6332 3016 6384
rect 6276 6400 6328 6452
rect 1768 6196 1820 6248
rect 1952 6196 2004 6248
rect 2780 6264 2832 6316
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 5080 6264 5132 6316
rect 2504 6196 2556 6248
rect 3516 6196 3568 6248
rect 3332 6128 3384 6180
rect 3424 6128 3476 6180
rect 4344 6196 4396 6248
rect 5632 6196 5684 6248
rect 1400 6060 1452 6112
rect 2780 6060 2832 6112
rect 4896 6128 4948 6180
rect 5908 6196 5960 6248
rect 6460 6264 6512 6316
rect 7196 6400 7248 6452
rect 9128 6400 9180 6452
rect 10508 6443 10560 6452
rect 10508 6409 10517 6443
rect 10517 6409 10551 6443
rect 10551 6409 10560 6443
rect 10508 6400 10560 6409
rect 9956 6332 10008 6384
rect 11520 6400 11572 6452
rect 12440 6400 12492 6452
rect 13084 6400 13136 6452
rect 13728 6400 13780 6452
rect 13912 6400 13964 6452
rect 15016 6332 15068 6384
rect 6644 6264 6696 6316
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 6736 6196 6788 6248
rect 7472 6196 7524 6248
rect 7656 6196 7708 6248
rect 10048 6264 10100 6316
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 4620 6060 4672 6112
rect 6920 6128 6972 6180
rect 9864 6196 9916 6248
rect 10232 6196 10284 6248
rect 10968 6196 11020 6248
rect 11152 6239 11204 6248
rect 11152 6205 11186 6239
rect 11186 6205 11204 6239
rect 11152 6196 11204 6205
rect 12624 6239 12676 6248
rect 12624 6205 12633 6239
rect 12633 6205 12667 6239
rect 12667 6205 12676 6239
rect 12624 6196 12676 6205
rect 13452 6196 13504 6248
rect 13728 6196 13780 6248
rect 17960 6196 18012 6248
rect 9496 6128 9548 6180
rect 5816 6060 5868 6112
rect 6736 6060 6788 6112
rect 8024 6060 8076 6112
rect 10600 6128 10652 6180
rect 11060 6128 11112 6180
rect 11980 6128 12032 6180
rect 12072 6128 12124 6180
rect 10140 6103 10192 6112
rect 10140 6069 10149 6103
rect 10149 6069 10183 6103
rect 10183 6069 10192 6103
rect 10140 6060 10192 6069
rect 10232 6060 10284 6112
rect 11336 6060 11388 6112
rect 12348 6060 12400 6112
rect 12808 6128 12860 6180
rect 14372 6128 14424 6180
rect 15016 6128 15068 6180
rect 12624 6060 12676 6112
rect 14464 6060 14516 6112
rect 17224 6060 17276 6112
rect 18236 6103 18288 6112
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 2412 5856 2464 5908
rect 3424 5856 3476 5908
rect 4528 5899 4580 5908
rect 4528 5865 4537 5899
rect 4537 5865 4571 5899
rect 4571 5865 4580 5899
rect 4528 5856 4580 5865
rect 1584 5720 1636 5772
rect 3516 5763 3568 5772
rect 3516 5729 3525 5763
rect 3525 5729 3559 5763
rect 3559 5729 3568 5763
rect 3516 5720 3568 5729
rect 6644 5856 6696 5908
rect 9864 5856 9916 5908
rect 10048 5856 10100 5908
rect 11152 5856 11204 5908
rect 11244 5856 11296 5908
rect 11612 5856 11664 5908
rect 12164 5899 12216 5908
rect 12164 5865 12173 5899
rect 12173 5865 12207 5899
rect 12207 5865 12216 5899
rect 12164 5856 12216 5865
rect 13360 5856 13412 5908
rect 13820 5856 13872 5908
rect 14096 5856 14148 5908
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 7104 5788 7156 5840
rect 9220 5788 9272 5840
rect 5632 5763 5684 5772
rect 5632 5729 5666 5763
rect 5666 5729 5684 5763
rect 5632 5720 5684 5729
rect 5908 5720 5960 5772
rect 12072 5788 12124 5840
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 10140 5763 10192 5772
rect 10140 5729 10174 5763
rect 10174 5729 10192 5763
rect 10140 5720 10192 5729
rect 11520 5720 11572 5772
rect 12440 5720 12492 5772
rect 12716 5720 12768 5772
rect 13636 5720 13688 5772
rect 13912 5720 13964 5772
rect 17500 5720 17552 5772
rect 18236 5763 18288 5772
rect 18236 5729 18245 5763
rect 18245 5729 18279 5763
rect 18279 5729 18288 5763
rect 18236 5720 18288 5729
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 5356 5584 5408 5636
rect 7472 5652 7524 5704
rect 8484 5652 8536 5704
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 10876 5652 10928 5704
rect 11336 5652 11388 5704
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 15016 5652 15068 5704
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 3056 5516 3108 5568
rect 3700 5516 3752 5568
rect 5540 5516 5592 5568
rect 7104 5516 7156 5568
rect 9864 5584 9916 5636
rect 11152 5584 11204 5636
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 8852 5516 8904 5568
rect 11060 5516 11112 5568
rect 11244 5559 11296 5568
rect 11244 5525 11253 5559
rect 11253 5525 11287 5559
rect 11287 5525 11296 5559
rect 11244 5516 11296 5525
rect 12164 5516 12216 5568
rect 14280 5584 14332 5636
rect 18420 5627 18472 5636
rect 18420 5593 18429 5627
rect 18429 5593 18463 5627
rect 18463 5593 18472 5627
rect 18420 5584 18472 5593
rect 13820 5516 13872 5568
rect 17868 5516 17920 5568
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 3240 5312 3292 5364
rect 3516 5312 3568 5364
rect 7288 5312 7340 5364
rect 9220 5355 9272 5364
rect 4620 5219 4672 5228
rect 1584 5108 1636 5160
rect 2872 5108 2924 5160
rect 4620 5185 4629 5219
rect 4629 5185 4663 5219
rect 4663 5185 4672 5219
rect 4620 5176 4672 5185
rect 5632 5176 5684 5228
rect 5172 5151 5224 5160
rect 5172 5117 5181 5151
rect 5181 5117 5215 5151
rect 5215 5117 5224 5151
rect 5172 5108 5224 5117
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 8760 5176 8812 5228
rect 9220 5321 9229 5355
rect 9229 5321 9263 5355
rect 9263 5321 9272 5355
rect 9220 5312 9272 5321
rect 9404 5312 9456 5364
rect 10600 5312 10652 5364
rect 10784 5312 10836 5364
rect 12716 5312 12768 5364
rect 9680 5244 9732 5296
rect 13544 5244 13596 5296
rect 18236 5312 18288 5364
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 8852 5108 8904 5160
rect 11060 5108 11112 5160
rect 11336 5151 11388 5160
rect 11336 5117 11345 5151
rect 11345 5117 11379 5151
rect 11379 5117 11388 5151
rect 11336 5108 11388 5117
rect 2320 4972 2372 5024
rect 3148 5015 3200 5024
rect 3148 4981 3157 5015
rect 3157 4981 3191 5015
rect 3191 4981 3200 5015
rect 3148 4972 3200 4981
rect 3516 5015 3568 5024
rect 3516 4981 3525 5015
rect 3525 4981 3559 5015
rect 3559 4981 3568 5015
rect 3516 4972 3568 4981
rect 3608 4972 3660 5024
rect 4436 5015 4488 5024
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 5448 4972 5500 5024
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 7380 4972 7432 5024
rect 8668 4972 8720 5024
rect 9128 4972 9180 5024
rect 9220 4972 9272 5024
rect 9864 4972 9916 5024
rect 11428 5040 11480 5092
rect 12072 5108 12124 5160
rect 13636 5176 13688 5228
rect 15016 5176 15068 5228
rect 13912 5108 13964 5160
rect 14280 5151 14332 5160
rect 14280 5117 14314 5151
rect 14314 5117 14332 5151
rect 15936 5151 15988 5160
rect 14280 5108 14332 5117
rect 15936 5117 15945 5151
rect 15945 5117 15979 5151
rect 15979 5117 15988 5151
rect 15936 5108 15988 5117
rect 16212 5108 16264 5160
rect 13636 5040 13688 5092
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 12440 4972 12492 5024
rect 13268 4972 13320 5024
rect 13544 4972 13596 5024
rect 15844 5015 15896 5024
rect 15844 4981 15853 5015
rect 15853 4981 15887 5015
rect 15887 4981 15896 5015
rect 15844 4972 15896 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 1860 4768 1912 4820
rect 3148 4768 3200 4820
rect 3516 4768 3568 4820
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 8852 4768 8904 4820
rect 10324 4768 10376 4820
rect 11612 4768 11664 4820
rect 14004 4768 14056 4820
rect 15844 4768 15896 4820
rect 3056 4700 3108 4752
rect 5632 4700 5684 4752
rect 7564 4700 7616 4752
rect 7748 4743 7800 4752
rect 7748 4709 7757 4743
rect 7757 4709 7791 4743
rect 7791 4709 7800 4743
rect 7748 4700 7800 4709
rect 3608 4632 3660 4684
rect 5172 4632 5224 4684
rect 6184 4632 6236 4684
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 4620 4607 4672 4616
rect 1584 4496 1636 4548
rect 2136 4496 2188 4548
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 3792 4496 3844 4548
rect 5080 4496 5132 4548
rect 2688 4428 2740 4480
rect 4252 4428 4304 4480
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 5356 4496 5408 4548
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 8484 4632 8536 4684
rect 9588 4700 9640 4752
rect 11244 4700 11296 4752
rect 12440 4743 12492 4752
rect 12440 4709 12449 4743
rect 12449 4709 12483 4743
rect 12483 4709 12492 4743
rect 12440 4700 12492 4709
rect 12624 4700 12676 4752
rect 17408 4700 17460 4752
rect 9496 4632 9548 4684
rect 8300 4564 8352 4616
rect 8760 4607 8812 4616
rect 5724 4428 5776 4480
rect 5908 4471 5960 4480
rect 5908 4437 5917 4471
rect 5917 4437 5951 4471
rect 5951 4437 5960 4471
rect 5908 4428 5960 4437
rect 6276 4428 6328 4480
rect 7380 4428 7432 4480
rect 8760 4573 8769 4607
rect 8769 4573 8803 4607
rect 8803 4573 8812 4607
rect 8760 4564 8812 4573
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 10692 4564 10744 4616
rect 14004 4632 14056 4684
rect 14096 4632 14148 4684
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 13912 4564 13964 4616
rect 8668 4496 8720 4548
rect 9220 4496 9272 4548
rect 9588 4428 9640 4480
rect 12256 4496 12308 4548
rect 13360 4496 13412 4548
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 18420 4564 18472 4616
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 11152 4471 11204 4480
rect 11152 4437 11161 4471
rect 11161 4437 11195 4471
rect 11195 4437 11204 4471
rect 11152 4428 11204 4437
rect 12440 4428 12492 4480
rect 13544 4428 13596 4480
rect 13820 4428 13872 4480
rect 14648 4428 14700 4480
rect 18052 4471 18104 4480
rect 18052 4437 18061 4471
rect 18061 4437 18095 4471
rect 18095 4437 18104 4471
rect 18052 4428 18104 4437
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 3608 4267 3660 4276
rect 3608 4233 3617 4267
rect 3617 4233 3651 4267
rect 3651 4233 3660 4267
rect 3608 4224 3660 4233
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 6368 4224 6420 4276
rect 8760 4224 8812 4276
rect 9220 4224 9272 4276
rect 9772 4224 9824 4276
rect 10324 4224 10376 4276
rect 11980 4224 12032 4276
rect 12072 4267 12124 4276
rect 12072 4233 12081 4267
rect 12081 4233 12115 4267
rect 12115 4233 12124 4267
rect 12072 4224 12124 4233
rect 12348 4224 12400 4276
rect 12808 4224 12860 4276
rect 4896 4156 4948 4208
rect 5448 4156 5500 4208
rect 6460 4156 6512 4208
rect 9404 4156 9456 4208
rect 5356 4088 5408 4140
rect 5632 4088 5684 4140
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 1492 3952 1544 4004
rect 2136 4020 2188 4072
rect 2320 4020 2372 4072
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 3884 4063 3936 4072
rect 3884 4029 3893 4063
rect 3893 4029 3927 4063
rect 3927 4029 3936 4063
rect 3884 4020 3936 4029
rect 5172 4020 5224 4072
rect 5816 4063 5868 4072
rect 5816 4029 5825 4063
rect 5825 4029 5859 4063
rect 5859 4029 5868 4063
rect 7656 4063 7708 4072
rect 5816 4020 5868 4029
rect 7656 4029 7665 4063
rect 7665 4029 7699 4063
rect 7699 4029 7708 4063
rect 7656 4020 7708 4029
rect 8944 4088 8996 4140
rect 11612 4156 11664 4208
rect 13084 4156 13136 4208
rect 14004 4224 14056 4276
rect 14464 4224 14516 4276
rect 17960 4224 18012 4276
rect 18420 4267 18472 4276
rect 18420 4233 18429 4267
rect 18429 4233 18463 4267
rect 18463 4233 18472 4267
rect 18420 4224 18472 4233
rect 13360 4131 13412 4140
rect 9312 4020 9364 4072
rect 9404 4020 9456 4072
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2044 3884 2096 3893
rect 4252 3952 4304 4004
rect 5356 3952 5408 4004
rect 7748 3952 7800 4004
rect 4344 3884 4396 3936
rect 6092 3884 6144 3936
rect 6736 3884 6788 3936
rect 7380 3884 7432 3936
rect 9220 3952 9272 4004
rect 9956 4020 10008 4072
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 8300 3884 8352 3936
rect 10600 3952 10652 4004
rect 11060 4020 11112 4072
rect 11888 4020 11940 4072
rect 13636 4020 13688 4072
rect 13544 3952 13596 4004
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 15016 4131 15068 4140
rect 15016 4097 15025 4131
rect 15025 4097 15059 4131
rect 15059 4097 15068 4131
rect 15016 4088 15068 4097
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 17960 4020 18012 4072
rect 9588 3884 9640 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12624 3884 12676 3893
rect 14004 3884 14056 3936
rect 15384 3884 15436 3936
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 1952 3680 2004 3732
rect 2320 3544 2372 3596
rect 5908 3680 5960 3732
rect 6644 3680 6696 3732
rect 7380 3723 7432 3732
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 3424 3612 3476 3664
rect 3332 3587 3384 3596
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 3700 3612 3752 3664
rect 7288 3612 7340 3664
rect 3792 3544 3844 3596
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 7472 3544 7524 3596
rect 8392 3680 8444 3732
rect 9128 3680 9180 3732
rect 10324 3680 10376 3732
rect 14648 3680 14700 3732
rect 17684 3723 17736 3732
rect 17684 3689 17693 3723
rect 17693 3689 17727 3723
rect 17727 3689 17736 3723
rect 17684 3680 17736 3689
rect 8944 3612 8996 3664
rect 9312 3612 9364 3664
rect 9680 3612 9732 3664
rect 11980 3612 12032 3664
rect 12164 3612 12216 3664
rect 2872 3408 2924 3460
rect 3056 3476 3108 3528
rect 4160 3476 4212 3528
rect 4896 3476 4948 3528
rect 5080 3476 5132 3528
rect 5264 3476 5316 3528
rect 5816 3476 5868 3528
rect 3700 3408 3752 3460
rect 3884 3451 3936 3460
rect 3884 3417 3893 3451
rect 3893 3417 3927 3451
rect 3927 3417 3936 3451
rect 3884 3408 3936 3417
rect 6552 3476 6604 3528
rect 8116 3544 8168 3596
rect 8484 3544 8536 3596
rect 10232 3544 10284 3596
rect 10416 3544 10468 3596
rect 8300 3476 8352 3528
rect 8944 3476 8996 3528
rect 10508 3476 10560 3528
rect 11244 3476 11296 3528
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 7748 3408 7800 3460
rect 12900 3544 12952 3596
rect 14096 3612 14148 3664
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 4896 3383 4948 3392
rect 4896 3349 4905 3383
rect 4905 3349 4939 3383
rect 4939 3349 4948 3383
rect 4896 3340 4948 3349
rect 4988 3340 5040 3392
rect 6368 3340 6420 3392
rect 6644 3340 6696 3392
rect 9772 3383 9824 3392
rect 9772 3349 9781 3383
rect 9781 3349 9815 3383
rect 9815 3349 9824 3383
rect 9772 3340 9824 3349
rect 10324 3340 10376 3392
rect 13268 3519 13320 3528
rect 13268 3485 13277 3519
rect 13277 3485 13311 3519
rect 13311 3485 13320 3519
rect 13268 3476 13320 3485
rect 17132 3519 17184 3528
rect 17132 3485 17141 3519
rect 17141 3485 17175 3519
rect 17175 3485 17184 3519
rect 17132 3476 17184 3485
rect 18420 3544 18472 3596
rect 15016 3408 15068 3460
rect 13636 3340 13688 3392
rect 17868 3340 17920 3392
rect 18420 3383 18472 3392
rect 18420 3349 18429 3383
rect 18429 3349 18463 3383
rect 18463 3349 18472 3383
rect 18420 3340 18472 3349
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 2596 3179 2648 3188
rect 2596 3145 2605 3179
rect 2605 3145 2639 3179
rect 2639 3145 2648 3179
rect 2596 3136 2648 3145
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 3056 3136 3108 3145
rect 3332 3136 3384 3188
rect 2780 3068 2832 3120
rect 3148 3068 3200 3120
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 4344 3068 4396 3120
rect 3608 3000 3660 3009
rect 1400 2932 1452 2984
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 2044 2932 2096 2984
rect 3424 2975 3476 2984
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 5816 3136 5868 3188
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 6736 3136 6788 3188
rect 5080 3068 5132 3120
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 8300 3136 8352 3188
rect 8944 3136 8996 3188
rect 10416 3136 10468 3188
rect 14004 3136 14056 3188
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 10876 3068 10928 3120
rect 5080 2932 5132 2984
rect 6000 2932 6052 2984
rect 9404 3000 9456 3052
rect 9680 3043 9732 3052
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 11060 3000 11112 3052
rect 5448 2907 5500 2916
rect 2596 2796 2648 2848
rect 5448 2873 5482 2907
rect 5482 2873 5500 2907
rect 5448 2864 5500 2873
rect 7656 2864 7708 2916
rect 4712 2796 4764 2848
rect 6368 2796 6420 2848
rect 10416 2932 10468 2984
rect 12256 3068 12308 3120
rect 11888 3043 11940 3052
rect 9956 2864 10008 2916
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 12532 3000 12584 3052
rect 13636 3000 13688 3052
rect 11520 2932 11572 2984
rect 11796 2932 11848 2984
rect 12348 2932 12400 2984
rect 14372 3068 14424 3120
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 15384 2932 15436 2984
rect 17408 2932 17460 2984
rect 17960 2932 18012 2984
rect 14832 2864 14884 2916
rect 14924 2864 14976 2916
rect 19432 2864 19484 2916
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 17776 2839 17828 2848
rect 17776 2805 17785 2839
rect 17785 2805 17819 2839
rect 17819 2805 17828 2839
rect 17776 2796 17828 2805
rect 18236 2839 18288 2848
rect 18236 2805 18245 2839
rect 18245 2805 18279 2839
rect 18279 2805 18288 2839
rect 18236 2796 18288 2805
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 1492 2635 1544 2644
rect 1492 2601 1501 2635
rect 1501 2601 1535 2635
rect 1535 2601 1544 2635
rect 1492 2592 1544 2601
rect 4436 2592 4488 2644
rect 5080 2635 5132 2644
rect 5080 2601 5089 2635
rect 5089 2601 5123 2635
rect 5123 2601 5132 2635
rect 5080 2592 5132 2601
rect 4896 2524 4948 2576
rect 1676 2456 1728 2508
rect 2136 2499 2188 2508
rect 2136 2465 2145 2499
rect 2145 2465 2179 2499
rect 2179 2465 2188 2499
rect 2136 2456 2188 2465
rect 2688 2499 2740 2508
rect 2688 2465 2697 2499
rect 2697 2465 2731 2499
rect 2731 2465 2740 2499
rect 2688 2456 2740 2465
rect 3424 2456 3476 2508
rect 1216 2388 1268 2440
rect 3056 2388 3108 2440
rect 2136 2320 2188 2372
rect 4988 2456 5040 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 8208 2592 8260 2644
rect 9956 2635 10008 2644
rect 9956 2601 9965 2635
rect 9965 2601 9999 2635
rect 9999 2601 10008 2635
rect 9956 2592 10008 2601
rect 11428 2592 11480 2644
rect 6736 2524 6788 2576
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 7840 2456 7892 2508
rect 9036 2524 9088 2576
rect 11704 2592 11756 2644
rect 12532 2592 12584 2644
rect 14004 2635 14056 2644
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 14924 2592 14976 2644
rect 16764 2635 16816 2644
rect 16764 2601 16773 2635
rect 16773 2601 16807 2635
rect 16807 2601 16816 2635
rect 16764 2592 16816 2601
rect 8576 2499 8628 2508
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 4804 2320 4856 2372
rect 4896 2320 4948 2372
rect 5816 2388 5868 2440
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 7564 2320 7616 2372
rect 8484 2320 8536 2372
rect 10876 2456 10928 2508
rect 13452 2524 13504 2576
rect 13176 2499 13228 2508
rect 13176 2465 13185 2499
rect 13185 2465 13219 2499
rect 13219 2465 13228 2499
rect 13176 2456 13228 2465
rect 15292 2456 15344 2508
rect 16948 2524 17000 2576
rect 11060 2388 11112 2440
rect 11336 2388 11388 2440
rect 12256 2388 12308 2440
rect 13084 2388 13136 2440
rect 13912 2388 13964 2440
rect 16672 2388 16724 2440
rect 16856 2388 16908 2440
rect 17224 2388 17276 2440
rect 11152 2320 11204 2372
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 3792 2295 3844 2304
rect 3792 2261 3801 2295
rect 3801 2261 3835 2295
rect 3835 2261 3844 2295
rect 3792 2252 3844 2261
rect 7472 2252 7524 2304
rect 10876 2252 10928 2304
rect 11428 2252 11480 2304
rect 16304 2295 16356 2304
rect 16304 2261 16313 2295
rect 16313 2261 16347 2295
rect 16347 2261 16356 2295
rect 16304 2252 16356 2261
rect 17316 2295 17368 2304
rect 17316 2261 17325 2295
rect 17325 2261 17359 2295
rect 17359 2261 17368 2295
rect 17316 2252 17368 2261
rect 17684 2295 17736 2304
rect 17684 2261 17693 2295
rect 17693 2261 17727 2295
rect 17727 2261 17736 2295
rect 17684 2252 17736 2261
rect 17868 2252 17920 2304
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 388 2048 440 2100
rect 16304 2048 16356 2100
<< metal2 >>
rect 1122 16400 1178 17200
rect 3238 16824 3294 16833
rect 3238 16759 3294 16768
rect 1136 13190 1164 16400
rect 1490 16008 1546 16017
rect 1490 15943 1546 15952
rect 1124 13184 1176 13190
rect 1124 13126 1176 13132
rect 1504 12238 1532 15943
rect 2134 14784 2190 14793
rect 2134 14719 2190 14728
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 2148 12102 2176 14719
rect 2594 13560 2650 13569
rect 2594 13495 2650 13504
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 1584 11620 1636 11626
rect 1584 11562 1636 11568
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 10606 1440 11494
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1400 10056 1452 10062
rect 1504 10044 1532 11086
rect 1452 10016 1532 10044
rect 1400 9998 1452 10004
rect 1412 9586 1440 9998
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 8498 1440 9522
rect 1596 9518 1624 11562
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1780 10810 1808 11494
rect 2424 11286 2452 11698
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1596 7478 1624 7890
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1596 7041 1624 7414
rect 1582 7032 1638 7041
rect 1582 6967 1638 6976
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 3913 1440 6054
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1596 5166 1624 5714
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1596 4554 1624 5102
rect 1584 4548 1636 4554
rect 1584 4490 1636 4496
rect 1492 4004 1544 4010
rect 1492 3946 1544 3952
rect 1398 3904 1454 3913
rect 1398 3839 1454 3848
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1216 2440 1268 2446
rect 1216 2382 1268 2388
rect 388 2100 440 2106
rect 388 2042 440 2048
rect 400 800 428 2042
rect 1228 800 1256 2382
rect 386 0 442 800
rect 1214 0 1270 800
rect 1412 241 1440 2926
rect 1504 2650 1532 3946
rect 1584 3936 1636 3942
rect 1582 3904 1584 3913
rect 1636 3904 1638 3913
rect 1582 3839 1638 3848
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1596 2553 1624 2926
rect 1582 2544 1638 2553
rect 1688 2514 1716 10406
rect 1872 8922 1900 11018
rect 1964 9042 1992 11154
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2056 10266 2084 10610
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2056 9518 2084 10202
rect 2608 10130 2636 13495
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2700 11354 2728 11630
rect 2792 11626 2820 12174
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2700 10198 2728 11290
rect 2792 11257 2820 11562
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2870 11384 2926 11393
rect 2870 11319 2926 11328
rect 2778 11248 2834 11257
rect 2778 11183 2834 11192
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2594 9616 2650 9625
rect 2594 9551 2650 9560
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2608 9178 2636 9551
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2700 9110 2728 10134
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2884 9042 2912 11319
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2976 10742 3004 11154
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 3068 10606 3096 11494
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2976 9178 3004 10474
rect 3148 10464 3200 10470
rect 3252 10441 3280 16759
rect 3330 16400 3386 17200
rect 3422 16416 3478 16425
rect 3344 14278 3372 16400
rect 5538 16400 5594 17200
rect 7746 16400 7802 17200
rect 9954 16400 10010 17200
rect 12162 16400 12218 17200
rect 14370 16400 14426 17200
rect 16486 16416 16542 16425
rect 3422 16351 3478 16360
rect 3436 15774 3464 16351
rect 3424 15768 3476 15774
rect 3424 15710 3476 15716
rect 4986 15192 5042 15201
rect 4986 15127 5042 15136
rect 4068 14408 4120 14414
rect 4066 14376 4068 14385
rect 4120 14376 4122 14385
rect 3792 14340 3844 14346
rect 4066 14311 4122 14320
rect 3792 14282 3844 14288
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3804 13977 3832 14282
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 3790 13968 3846 13977
rect 3790 13903 3846 13912
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 3698 13152 3754 13161
rect 3698 13087 3754 13096
rect 3712 12986 3740 13087
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 4356 12782 4384 13262
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 3804 12238 3832 12718
rect 3976 12368 4028 12374
rect 3974 12336 3976 12345
rect 4028 12336 4030 12345
rect 3974 12271 4030 12280
rect 3792 12232 3844 12238
rect 3606 12200 3662 12209
rect 3792 12174 3844 12180
rect 3606 12135 3662 12144
rect 3422 11928 3478 11937
rect 3620 11898 3648 12135
rect 3422 11863 3478 11872
rect 3608 11892 3660 11898
rect 3436 10810 3464 11863
rect 3608 11834 3660 11840
rect 3620 11286 3648 11834
rect 3804 11676 3832 12174
rect 4252 12096 4304 12102
rect 4712 12096 4764 12102
rect 4252 12038 4304 12044
rect 4540 12056 4712 12084
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3884 11688 3936 11694
rect 3804 11648 3884 11676
rect 3884 11630 3936 11636
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3608 11144 3660 11150
rect 3514 11112 3570 11121
rect 3608 11086 3660 11092
rect 3514 11047 3570 11056
rect 3424 10804 3476 10810
rect 3344 10764 3424 10792
rect 3148 10406 3200 10412
rect 3238 10432 3294 10441
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2780 8968 2832 8974
rect 1872 8894 1992 8922
rect 2780 8910 2832 8916
rect 2962 8936 3018 8945
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1768 7744 1820 7750
rect 1872 7721 1900 8774
rect 1768 7686 1820 7692
rect 1858 7712 1914 7721
rect 1780 6905 1808 7686
rect 1858 7647 1914 7656
rect 1964 6905 1992 8894
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2148 8090 2176 8774
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2502 7848 2558 7857
rect 2502 7783 2558 7792
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2148 6934 2176 7686
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2136 6928 2188 6934
rect 1766 6896 1822 6905
rect 1950 6896 2006 6905
rect 1766 6831 1822 6840
rect 1860 6860 1912 6866
rect 2136 6870 2188 6876
rect 1950 6831 2006 6840
rect 1860 6802 1912 6808
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1780 6254 1808 6666
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1780 4185 1808 6190
rect 1872 4826 1900 6802
rect 1964 6254 1992 6831
rect 2424 6798 2452 7278
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 2042 4992 2098 5001
rect 2042 4927 2098 4936
rect 1860 4820 1912 4826
rect 1912 4780 1992 4808
rect 1860 4762 1912 4768
rect 1766 4176 1822 4185
rect 1766 4111 1822 4120
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1872 3505 1900 3878
rect 1964 3738 1992 4780
rect 2056 3942 2084 4927
rect 2136 4548 2188 4554
rect 2136 4490 2188 4496
rect 2148 4078 2176 4490
rect 2136 4072 2188 4078
rect 2134 4040 2136 4049
rect 2188 4040 2190 4049
rect 2134 3975 2190 3984
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1582 2479 1638 2488
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1872 2281 1900 3334
rect 2056 2990 2084 3878
rect 2240 3618 2268 6598
rect 2424 5914 2452 6734
rect 2516 6254 2544 7783
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2332 4622 2360 4966
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2332 4078 2360 4558
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2318 3904 2374 3913
rect 2318 3839 2374 3848
rect 2148 3590 2268 3618
rect 2332 3602 2360 3839
rect 2320 3596 2372 3602
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2148 2514 2176 3590
rect 2320 3538 2372 3544
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 2689 2268 3334
rect 2608 3194 2636 8570
rect 2792 8430 2820 8910
rect 2962 8871 3018 8880
rect 2976 8634 3004 8871
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2976 8430 3004 8570
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2884 7886 2912 8230
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2884 7274 2912 7822
rect 2872 7268 2924 7274
rect 2872 7210 2924 7216
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6866 2820 7142
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2778 6488 2834 6497
rect 2884 6458 2912 6938
rect 2778 6423 2834 6432
rect 2872 6452 2924 6458
rect 2792 6322 2820 6423
rect 2872 6394 2924 6400
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 4729 2820 6054
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5166 2912 5510
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2778 4720 2834 4729
rect 2778 4655 2834 4664
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2608 2854 2636 3130
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2226 2680 2282 2689
rect 2226 2615 2282 2624
rect 2700 2514 2728 4422
rect 2976 4321 3004 6326
rect 3068 5658 3096 9318
rect 3160 9178 3188 10406
rect 3238 10367 3294 10376
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 8090 3188 8230
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3344 7834 3372 10764
rect 3424 10746 3476 10752
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10130 3464 10406
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 9178 3464 9862
rect 3528 9761 3556 11047
rect 3620 10169 3648 11086
rect 3700 11008 3752 11014
rect 3698 10976 3700 10985
rect 3752 10976 3754 10985
rect 3698 10911 3754 10920
rect 3804 10674 3832 11494
rect 3896 11082 3924 11630
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3606 10160 3662 10169
rect 3606 10095 3662 10104
rect 3804 10062 3832 10610
rect 4158 10160 4214 10169
rect 4158 10095 4214 10104
rect 4172 10062 4200 10095
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3514 9752 3570 9761
rect 3921 9744 4217 9764
rect 3514 9687 3570 9696
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3436 8945 3464 8978
rect 3422 8936 3478 8945
rect 3422 8871 3478 8880
rect 3424 8560 3476 8566
rect 3422 8528 3424 8537
rect 3476 8528 3478 8537
rect 3422 8463 3478 8472
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3436 7886 3464 8298
rect 3528 7886 3556 9687
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3712 8498 3740 9386
rect 4172 9382 4200 9413
rect 4160 9376 4212 9382
rect 4158 9344 4160 9353
rect 4212 9344 4214 9353
rect 4158 9279 4214 9288
rect 4172 9178 4200 9279
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3700 8288 3752 8294
rect 3804 8276 3832 8774
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3976 8424 4028 8430
rect 3974 8392 3976 8401
rect 4028 8392 4030 8401
rect 4264 8378 4292 12038
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4356 10305 4384 11086
rect 4540 11014 4568 12056
rect 4712 12038 4764 12044
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4448 10470 4476 10950
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4342 10296 4398 10305
rect 4448 10266 4476 10406
rect 4342 10231 4398 10240
rect 4436 10260 4488 10266
rect 4356 10198 4384 10231
rect 4436 10202 4488 10208
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4356 8514 4384 9658
rect 4448 9654 4476 9930
rect 4436 9648 4488 9654
rect 4540 9625 4568 10950
rect 4632 10674 4660 11630
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4632 10044 4660 10610
rect 4712 10600 4764 10606
rect 4908 10588 4936 10950
rect 4764 10577 4936 10588
rect 4764 10568 4950 10577
rect 4764 10560 4894 10568
rect 4712 10542 4764 10548
rect 4894 10503 4950 10512
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4894 10432 4950 10441
rect 4712 10056 4764 10062
rect 4632 10016 4712 10044
rect 4712 9998 4764 10004
rect 4436 9590 4488 9596
rect 4526 9616 4582 9625
rect 4582 9574 4660 9602
rect 4724 9586 4752 9998
rect 4526 9551 4582 9560
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4526 9480 4582 9489
rect 4448 8634 4476 9454
rect 4632 9466 4660 9574
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4816 9518 4844 10406
rect 4894 10367 4950 10376
rect 4804 9512 4856 9518
rect 4632 9438 4752 9466
rect 4804 9454 4856 9460
rect 4526 9415 4582 9424
rect 4540 9178 4568 9415
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4356 8486 4476 8514
rect 4264 8350 4384 8378
rect 3974 8327 4030 8336
rect 3752 8248 3832 8276
rect 4252 8288 4304 8294
rect 3700 8230 3752 8236
rect 4252 8230 4304 8236
rect 3712 7970 3740 8230
rect 3790 8120 3846 8129
rect 3790 8055 3792 8064
rect 3844 8055 3846 8064
rect 3792 8026 3844 8032
rect 3712 7942 3832 7970
rect 3160 7806 3372 7834
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3608 7812 3660 7818
rect 3160 5760 3188 7806
rect 3608 7754 3660 7760
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3252 6089 3280 7142
rect 3344 6186 3372 7686
rect 3620 7410 3648 7754
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3436 6322 3464 7210
rect 3516 7200 3568 7206
rect 3712 7177 3740 7822
rect 3516 7142 3568 7148
rect 3698 7168 3754 7177
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3528 6254 3556 7142
rect 3698 7103 3754 7112
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3620 6458 3648 6938
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3238 6080 3294 6089
rect 3238 6015 3294 6024
rect 3436 5914 3464 6122
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3516 5772 3568 5778
rect 3160 5732 3280 5760
rect 3068 5630 3188 5658
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 4758 3096 5510
rect 3160 5137 3188 5630
rect 3252 5370 3280 5732
rect 3516 5714 3568 5720
rect 3528 5370 3556 5714
rect 3700 5568 3752 5574
rect 3698 5536 3700 5545
rect 3752 5536 3754 5545
rect 3698 5471 3754 5480
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3146 5128 3202 5137
rect 3252 5114 3280 5306
rect 3252 5086 3648 5114
rect 3146 5063 3202 5072
rect 3620 5030 3648 5086
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3160 4826 3188 4966
rect 3528 4826 3556 4966
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 2962 4312 3018 4321
rect 3620 4282 3648 4626
rect 3804 4554 3832 7942
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4264 7342 4292 8230
rect 4356 8090 4384 8350
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4252 7336 4304 7342
rect 4066 7304 4122 7313
rect 4252 7278 4304 7284
rect 4066 7239 4122 7248
rect 4080 7206 4108 7239
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4356 6934 4384 7890
rect 4448 7886 4476 8486
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4434 7032 4490 7041
rect 4632 7002 4660 9318
rect 4434 6967 4490 6976
rect 4620 6996 4672 7002
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 4356 6254 4384 6666
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4448 5658 4476 6967
rect 4620 6938 4672 6944
rect 4724 6934 4752 9438
rect 4816 9110 4844 9454
rect 4908 9178 4936 10367
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4816 7750 4844 8026
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4816 7002 4844 7142
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 5914 4568 6598
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4632 5710 4660 6054
rect 4620 5704 4672 5710
rect 4448 5630 4568 5658
rect 4620 5646 4672 5652
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4436 5024 4488 5030
rect 4434 4992 4436 5001
rect 4488 4992 4490 5001
rect 4434 4927 4490 4936
rect 4540 4826 4568 5630
rect 4632 5234 4660 5646
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4540 4729 4568 4762
rect 4526 4720 4582 4729
rect 4526 4655 4582 4664
rect 4632 4622 4660 5170
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 2962 4247 3018 4256
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2780 3120 2832 3126
rect 2884 3097 2912 3402
rect 3068 3194 3096 3470
rect 3344 3194 3372 3538
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3148 3120 3200 3126
rect 2780 3062 2832 3068
rect 2870 3088 2926 3097
rect 2136 2508 2188 2514
rect 2136 2450 2188 2456
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2136 2372 2188 2378
rect 2136 2314 2188 2320
rect 1858 2272 1914 2281
rect 1858 2207 1914 2216
rect 2148 800 2176 2314
rect 2792 1873 2820 3062
rect 3148 3062 3200 3068
rect 2870 3023 2926 3032
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 2778 1864 2834 1873
rect 2778 1799 2834 1808
rect 3068 800 3096 2382
rect 3160 1465 3188 3062
rect 3436 2990 3464 3606
rect 3620 3058 3648 4218
rect 3804 4078 3832 4490
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4342 4448 4398 4457
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3792 4072 3844 4078
rect 3884 4072 3936 4078
rect 3792 4014 3844 4020
rect 3882 4040 3884 4049
rect 3936 4040 3938 4049
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3712 3466 3740 3606
rect 3804 3602 3832 4014
rect 4264 4010 4292 4422
rect 4342 4383 4398 4392
rect 3882 3975 3938 3984
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4264 3618 4292 3946
rect 4356 3942 4384 4383
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 4172 3590 4292 3618
rect 4436 3596 4488 3602
rect 4172 3534 4200 3590
rect 4436 3538 4488 3544
rect 4160 3528 4212 3534
rect 3882 3496 3938 3505
rect 3700 3460 3752 3466
rect 4160 3470 4212 3476
rect 4342 3496 4398 3505
rect 3882 3431 3884 3440
rect 3700 3402 3752 3408
rect 3936 3431 3938 3440
rect 4342 3431 4398 3440
rect 3884 3402 3936 3408
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4356 3126 4384 3431
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3436 2514 3464 2926
rect 4448 2650 4476 3538
rect 4724 2854 4752 6870
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3146 1456 3202 1465
rect 3146 1391 3202 1400
rect 1398 232 1454 241
rect 1398 167 1454 176
rect 2134 0 2190 800
rect 3054 0 3110 800
rect 3436 649 3464 2246
rect 3804 1057 3832 2246
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 4264 1442 4292 2382
rect 4816 2378 4844 6802
rect 4908 6186 4936 7346
rect 5000 6440 5028 15127
rect 5552 13802 5580 16400
rect 6644 15768 6696 15774
rect 6644 15710 6696 15716
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5920 14074 5948 14418
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5736 12986 5764 13330
rect 6012 13190 6040 13874
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6104 13530 6132 13670
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6000 13184 6052 13190
rect 5920 13144 6000 13172
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5552 12238 5580 12922
rect 5920 12374 5948 13144
rect 6000 13126 6052 13132
rect 6380 12986 6408 13670
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 12442 6040 12582
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5368 11150 5396 11766
rect 5460 11694 5488 12038
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5552 11218 5580 11630
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5092 10810 5120 10950
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5092 9994 5120 10474
rect 5184 10266 5212 10474
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 5092 6866 5120 9386
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5184 8090 5212 9114
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5184 7546 5212 8026
rect 5276 7818 5304 11018
rect 5552 10810 5580 11154
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5446 10704 5502 10713
rect 5644 10690 5672 11494
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5502 10662 5672 10690
rect 5446 10639 5502 10648
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 8634 5396 9862
rect 5552 9654 5580 9998
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5644 9466 5672 10662
rect 5736 10062 5764 11154
rect 5828 10674 5856 11562
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5460 9438 5672 9466
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5000 6412 5212 6440
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 5092 4554 5120 6258
rect 5184 5273 5212 6412
rect 5368 5642 5396 8570
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5460 5522 5488 9438
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5644 8022 5672 8434
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5552 6730 5580 7890
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5644 6254 5672 7142
rect 5736 6730 5764 8502
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5828 8022 5856 8366
rect 5816 8016 5868 8022
rect 5816 7958 5868 7964
rect 5828 7546 5856 7958
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5828 6882 5856 7210
rect 5920 7002 5948 12174
rect 6012 9194 6040 12242
rect 6196 12238 6224 12650
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6472 11558 6500 12310
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 10810 6224 11154
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6366 10296 6422 10305
rect 6366 10231 6368 10240
rect 6420 10231 6422 10240
rect 6368 10202 6420 10208
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6104 9382 6132 9862
rect 6196 9586 6224 10134
rect 6366 10024 6422 10033
rect 6366 9959 6422 9968
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6012 9166 6132 9194
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6012 8294 6040 8978
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 7993 6040 8230
rect 5998 7984 6054 7993
rect 5998 7919 6054 7928
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6012 7002 6040 7822
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5828 6854 5948 6882
rect 5920 6798 5948 6854
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5828 6338 5856 6598
rect 5828 6310 5948 6338
rect 5920 6254 5948 6310
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5276 5494 5488 5522
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5170 5264 5226 5273
rect 5170 5199 5226 5208
rect 5184 5166 5212 5199
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5184 4690 5212 5102
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4548 5132 4554
rect 5080 4490 5132 4496
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4908 3534 4936 4150
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4908 2582 4936 3334
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5000 2514 5028 3334
rect 5092 3126 5120 3470
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 5184 3058 5212 4014
rect 5276 3534 5304 5494
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4282 5396 4490
rect 5460 4457 5488 4966
rect 5446 4448 5502 4457
rect 5446 4383 5502 4392
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5368 4010 5396 4082
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5092 2650 5120 2926
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 5368 2446 5396 3946
rect 5460 2922 5488 4150
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 5552 2514 5580 5510
rect 5644 5234 5672 5714
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4758 5672 4966
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5644 4146 5672 4558
rect 5724 4480 5776 4486
rect 5828 4468 5856 6054
rect 5920 5778 5948 6190
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 6104 4978 6132 9166
rect 6196 8809 6224 9522
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6182 8800 6238 8809
rect 6182 8735 6238 8744
rect 6288 8634 6316 9318
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6288 8537 6316 8570
rect 6274 8528 6330 8537
rect 6274 8463 6330 8472
rect 6276 8288 6328 8294
rect 6380 8276 6408 9959
rect 6472 8566 6500 10542
rect 6552 10464 6604 10470
rect 6550 10432 6552 10441
rect 6604 10432 6606 10441
rect 6550 10367 6606 10376
rect 6656 10010 6684 15710
rect 6734 15600 6790 15609
rect 6734 15535 6790 15544
rect 6748 14074 6776 15535
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6748 13410 6776 14010
rect 7760 13870 7788 16400
rect 9968 14634 9996 16400
rect 9968 14606 10272 14634
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8208 14000 8260 14006
rect 8956 13954 8984 14282
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 8208 13942 8260 13948
rect 7196 13864 7248 13870
rect 7748 13864 7800 13870
rect 7248 13824 7328 13852
rect 7196 13806 7248 13812
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 6748 13394 6868 13410
rect 6748 13388 6880 13394
rect 6748 13382 6828 13388
rect 6828 13330 6880 13336
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 12714 6776 13262
rect 6840 13190 6868 13330
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 7300 12782 7328 13824
rect 7748 13806 7800 13812
rect 8220 13530 8248 13942
rect 8864 13926 8984 13954
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8208 13524 8260 13530
rect 8036 13484 8208 13512
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 7392 12442 7420 12650
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6748 11898 6776 12242
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6932 11626 6960 12242
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6932 10606 6960 11018
rect 7024 10810 7052 11086
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 7300 10266 7328 11154
rect 7392 11121 7420 12174
rect 7484 11558 7512 12582
rect 7576 11830 7604 12718
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7668 12238 7696 12582
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7564 11824 7616 11830
rect 7564 11766 7616 11772
rect 7932 11688 7984 11694
rect 7852 11648 7932 11676
rect 7564 11620 7616 11626
rect 7564 11562 7616 11568
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7472 11144 7524 11150
rect 7378 11112 7434 11121
rect 7576 11121 7604 11562
rect 7852 11218 7880 11648
rect 7932 11630 7984 11636
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7472 11086 7524 11092
rect 7562 11112 7618 11121
rect 7378 11047 7434 11056
rect 7484 10810 7512 11086
rect 7562 11047 7618 11056
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7852 10690 7880 11154
rect 7564 10668 7616 10674
rect 7852 10662 7972 10690
rect 7564 10610 7616 10616
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7392 10198 7420 10406
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6656 9982 6868 10010
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6328 8248 6408 8276
rect 6276 8230 6328 8236
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6012 4950 6132 4978
rect 5776 4440 5856 4468
rect 5908 4480 5960 4486
rect 5724 4422 5776 4428
rect 5908 4422 5960 4428
rect 5814 4176 5870 4185
rect 5632 4140 5684 4146
rect 5814 4111 5870 4120
rect 5632 4082 5684 4088
rect 5828 4078 5856 4111
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5920 3738 5948 4422
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 6012 3641 6040 4950
rect 6196 4842 6224 7686
rect 6288 7342 6316 8230
rect 6472 7410 6500 8298
rect 6656 8022 6684 9982
rect 6840 9625 6868 9982
rect 6932 9926 6960 10066
rect 7380 10056 7432 10062
rect 7300 10016 7380 10044
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6826 9616 6882 9625
rect 7024 9586 7052 9930
rect 6826 9551 6882 9560
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 7300 9081 7328 10016
rect 7484 10044 7512 10202
rect 7576 10062 7604 10610
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7432 10016 7512 10044
rect 7564 10056 7616 10062
rect 7380 9998 7432 10004
rect 7564 9998 7616 10004
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7392 9110 7420 9386
rect 7484 9217 7512 9862
rect 7470 9208 7526 9217
rect 7470 9143 7526 9152
rect 7380 9104 7432 9110
rect 7010 9072 7066 9081
rect 7010 9007 7066 9016
rect 7286 9072 7342 9081
rect 7380 9046 7432 9052
rect 7286 9007 7342 9016
rect 7472 9036 7524 9042
rect 7024 8498 7052 9007
rect 7472 8978 7524 8984
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7024 8401 7052 8434
rect 7208 8430 7236 8774
rect 7378 8664 7434 8673
rect 7378 8599 7434 8608
rect 7196 8424 7248 8430
rect 7010 8392 7066 8401
rect 6736 8356 6788 8362
rect 7196 8366 7248 8372
rect 7010 8327 7066 8336
rect 6736 8298 6788 8304
rect 6748 8022 6776 8298
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7410 6592 7686
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 7177 6408 7278
rect 6366 7168 6422 7177
rect 6366 7103 6422 7112
rect 6380 6866 6408 7103
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6276 6792 6328 6798
rect 6380 6769 6408 6802
rect 6276 6734 6328 6740
rect 6366 6760 6422 6769
rect 6288 6458 6316 6734
rect 6366 6695 6422 6704
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6472 6322 6500 7346
rect 7024 7342 7052 7754
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 6840 6361 6868 6802
rect 7208 6458 7236 6802
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 6826 6352 6882 6361
rect 6460 6316 6512 6322
rect 6644 6316 6696 6322
rect 6512 6276 6592 6304
rect 6460 6258 6512 6264
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6104 4814 6224 4842
rect 6104 3942 6132 4814
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6196 4146 6224 4626
rect 6288 4486 6316 4966
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6380 4282 6408 4966
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6472 4214 6500 4558
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 5998 3632 6054 3641
rect 6564 3618 6592 6276
rect 6826 6287 6828 6296
rect 6644 6258 6696 6264
rect 6880 6287 6882 6296
rect 6828 6258 6880 6264
rect 6656 5914 6684 6258
rect 6736 6248 6788 6254
rect 6788 6196 6868 6202
rect 6736 6190 6868 6196
rect 6748 6174 6868 6190
rect 6840 6168 6868 6174
rect 6920 6180 6972 6186
rect 6840 6140 6920 6168
rect 6920 6122 6972 6128
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6642 4992 6698 5001
rect 6642 4927 6698 4936
rect 6656 4049 6684 4927
rect 6748 4826 6776 6054
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 7116 5574 7144 5782
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7300 5370 7328 5646
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 6920 5160 6972 5166
rect 6918 5128 6920 5137
rect 6972 5128 6974 5137
rect 7392 5114 7420 8599
rect 7484 8498 7512 8978
rect 7576 8838 7604 9998
rect 7668 9382 7696 10066
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7654 9208 7710 9217
rect 7654 9143 7710 9152
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7484 7954 7512 8298
rect 7668 8072 7696 9143
rect 7576 8044 7696 8072
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7484 7857 7512 7890
rect 7470 7848 7526 7857
rect 7470 7783 7526 7792
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 5710 7512 6190
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 6918 5063 6974 5072
rect 7300 5086 7420 5114
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6918 4720 6974 4729
rect 6918 4655 6920 4664
rect 6972 4655 6974 4664
rect 6920 4626 6972 4632
rect 6642 4040 6698 4049
rect 6642 3975 6698 3984
rect 6656 3738 6684 3975
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6564 3590 6684 3618
rect 5998 3567 6054 3576
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5828 3194 5856 3470
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6012 2990 6040 3567
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6380 2854 6408 3334
rect 6564 3194 6592 3470
rect 6656 3398 6684 3590
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6748 3194 6776 3878
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 7300 3670 7328 5086
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4486 7420 4966
rect 7576 4758 7604 8044
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7668 7410 7696 7890
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7668 6361 7696 7210
rect 7654 6352 7710 6361
rect 7654 6287 7710 6296
rect 7668 6254 7696 6287
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 5574 7696 6190
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 5137 7696 5510
rect 7654 5128 7710 5137
rect 7654 5063 7710 5072
rect 7564 4752 7616 4758
rect 7562 4720 7564 4729
rect 7616 4720 7618 4729
rect 7562 4655 7618 4664
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 4146 7420 4422
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7668 4078 7696 5063
rect 7760 4758 7788 9386
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7760 4185 7788 4694
rect 7746 4176 7802 4185
rect 7746 4111 7802 4120
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3738 7420 3878
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 6736 2576 6788 2582
rect 6736 2518 6788 2524
rect 6918 2544 6974 2553
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 3988 1414 4292 1442
rect 3790 1048 3846 1057
rect 3790 983 3846 992
rect 3988 800 4016 1414
rect 4908 800 4936 2314
rect 5828 800 5856 2382
rect 6748 800 6776 2518
rect 6918 2479 6920 2488
rect 6972 2479 6974 2488
rect 6920 2450 6972 2456
rect 7484 2310 7512 3538
rect 7668 2922 7696 4014
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7760 3466 7788 3946
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 7852 2514 7880 10406
rect 7944 10130 7972 10662
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7944 9042 7972 10066
rect 8036 10033 8064 13484
rect 8208 13466 8260 13472
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8128 12322 8156 13330
rect 8404 12782 8432 13670
rect 8668 13456 8720 13462
rect 8668 13398 8720 13404
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8208 12368 8260 12374
rect 8128 12316 8208 12322
rect 8128 12310 8260 12316
rect 8128 12294 8248 12310
rect 8404 12238 8432 12718
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11762 8432 12174
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8298 11248 8354 11257
rect 8220 10674 8248 11222
rect 8298 11183 8300 11192
rect 8352 11183 8354 11192
rect 8300 11154 8352 11160
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8206 10568 8262 10577
rect 8206 10503 8262 10512
rect 8022 10024 8078 10033
rect 8022 9959 8078 9968
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8022 9616 8078 9625
rect 8022 9551 8024 9560
rect 8076 9551 8078 9560
rect 8024 9522 8076 9528
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 6730 7972 7822
rect 8036 7546 8064 7890
rect 8128 7834 8156 9658
rect 8220 9654 8248 10503
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9178 8248 9318
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8022 8340 8910
rect 8404 8294 8432 8978
rect 8496 8809 8524 9590
rect 8588 9489 8616 13262
rect 8574 9480 8630 9489
rect 8574 9415 8630 9424
rect 8576 8832 8628 8838
rect 8482 8800 8538 8809
rect 8576 8774 8628 8780
rect 8482 8735 8538 8744
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8128 7806 8340 7834
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 8036 6118 8064 7142
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8128 3602 8156 7806
rect 8312 7750 8340 7806
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8220 2650 8248 7686
rect 8404 6662 8432 8230
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 3942 8340 4558
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8312 3534 8340 3878
rect 8404 3738 8432 6598
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8496 4690 8524 5646
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8496 4593 8524 4626
rect 8482 4584 8538 4593
rect 8482 4519 8538 4528
rect 8482 4040 8538 4049
rect 8482 3975 8538 3984
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8496 3602 8524 3975
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8312 3194 8340 3470
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8588 2514 8616 8774
rect 8680 8362 8708 13398
rect 8758 12744 8814 12753
rect 8758 12679 8814 12688
rect 8772 11150 8800 12679
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8864 10810 8892 13926
rect 10244 13734 10272 14606
rect 12176 14550 12204 16400
rect 13450 14784 13506 14793
rect 12817 14716 13113 14736
rect 13450 14719 13506 14728
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 10414 13832 10470 13841
rect 10414 13767 10470 13776
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 9128 13320 9180 13326
rect 8956 13280 9128 13308
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8864 10606 8892 10746
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8864 9722 8892 10542
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8758 8528 8814 8537
rect 8758 8463 8760 8472
rect 8812 8463 8814 8472
rect 8760 8434 8812 8440
rect 8956 8412 8984 13280
rect 9128 13262 9180 13268
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12374 9352 13126
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9036 12300 9088 12306
rect 9088 12260 9168 12288
rect 9036 12242 9088 12248
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9048 9178 9076 12038
rect 9140 10810 9168 12260
rect 9692 12238 9720 12378
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9312 12232 9364 12238
rect 9588 12232 9640 12238
rect 9364 12192 9444 12220
rect 9508 12209 9588 12220
rect 9312 12174 9364 12180
rect 9232 12050 9260 12174
rect 9232 12022 9352 12050
rect 9324 11898 9352 12022
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9232 11778 9260 11834
rect 9232 11750 9352 11778
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9232 11354 9260 11562
rect 9324 11354 9352 11750
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9416 11200 9444 12192
rect 9494 12200 9588 12209
rect 9550 12192 9588 12200
rect 9588 12174 9640 12180
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9494 12135 9550 12144
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 10244 11694 10272 12038
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10232 11688 10284 11694
rect 10138 11656 10194 11665
rect 10232 11630 10284 11636
rect 10138 11591 10194 11600
rect 10152 11558 10180 11591
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9324 11172 9444 11200
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9324 10470 9352 11172
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 10674 9444 11018
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10198 9536 10406
rect 9496 10192 9548 10198
rect 9402 10160 9458 10169
rect 9496 10134 9548 10140
rect 9402 10095 9404 10104
rect 9456 10095 9458 10104
rect 9404 10066 9456 10072
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9382 9260 9998
rect 9416 9926 9444 10066
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9324 9110 9352 9862
rect 9508 9586 9536 10134
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9324 8974 9352 9046
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 8864 8384 8984 8412
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8864 8276 8892 8384
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 8944 8288 8996 8294
rect 8864 8248 8944 8276
rect 8944 8230 8996 8236
rect 8758 7984 8814 7993
rect 8758 7919 8814 7928
rect 8772 7886 8800 7919
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8956 7342 8984 8230
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8666 5264 8722 5273
rect 8772 5234 8800 5646
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8666 5199 8722 5208
rect 8760 5228 8812 5234
rect 8680 5030 8708 5199
rect 8760 5170 8812 5176
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8680 4554 8708 4966
rect 8772 4622 8800 5170
rect 8864 5166 8892 5510
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8772 4282 8800 4558
rect 8864 4457 8892 4762
rect 8850 4448 8906 4457
rect 8850 4383 8906 4392
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8956 4146 8984 7278
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8956 3534 8984 3606
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8956 3194 8984 3470
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9048 2582 9076 8298
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7750 9260 8230
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9126 7304 9182 7313
rect 9126 7239 9182 7248
rect 9140 6905 9168 7239
rect 9126 6896 9182 6905
rect 9126 6831 9128 6840
rect 9180 6831 9182 6840
rect 9128 6802 9180 6808
rect 9140 6458 9168 6802
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9140 5030 9168 6394
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9232 5370 9260 5782
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9232 4554 9260 4966
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9232 4010 9260 4218
rect 9324 4078 9352 7919
rect 9416 7732 9444 9454
rect 9496 7744 9548 7750
rect 9416 7704 9496 7732
rect 9496 7686 9548 7692
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 6186 9536 7142
rect 9600 6730 9628 11086
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 9586 9720 10474
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9784 9518 9812 10542
rect 10336 10538 10364 11766
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9692 8090 9720 9386
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9416 4622 9444 5306
rect 9508 4690 9536 6122
rect 9600 4758 9628 6666
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 5302 9720 6598
rect 9784 6372 9812 9318
rect 10060 9110 10088 9318
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 10138 8528 10194 8537
rect 10138 8463 10140 8472
rect 10192 8463 10194 8472
rect 10140 8434 10192 8440
rect 10046 7848 10102 7857
rect 10046 7783 10048 7792
rect 10100 7783 10102 7792
rect 10048 7754 10100 7760
rect 10152 7732 10180 8434
rect 10244 8090 10272 9998
rect 10336 9761 10364 10202
rect 10428 10130 10456 13767
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 12102 10640 12242
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10692 11824 10744 11830
rect 10690 11792 10692 11801
rect 10744 11792 10746 11801
rect 10600 11756 10652 11762
rect 10690 11727 10746 11736
rect 10600 11698 10652 11704
rect 10612 11558 10640 11698
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10336 7886 10364 9318
rect 10428 9081 10456 9862
rect 10414 9072 10470 9081
rect 10414 9007 10470 9016
rect 10520 8616 10548 11154
rect 10704 11150 10732 11222
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10612 9382 10640 10474
rect 10690 10024 10746 10033
rect 10690 9959 10692 9968
rect 10744 9959 10746 9968
rect 10692 9930 10744 9936
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10598 8936 10654 8945
rect 10704 8906 10732 9318
rect 10598 8871 10654 8880
rect 10692 8900 10744 8906
rect 10612 8838 10640 8871
rect 10692 8842 10744 8848
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10428 8588 10548 8616
rect 10428 7993 10456 8588
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10520 8090 10548 8434
rect 10612 8090 10640 8774
rect 10704 8362 10732 8842
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10414 7984 10470 7993
rect 10414 7919 10470 7928
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10152 7704 10364 7732
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 10230 7576 10286 7585
rect 10230 7511 10286 7520
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10060 6798 10088 7346
rect 10244 7342 10272 7511
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10244 7018 10272 7278
rect 10336 7188 10364 7704
rect 10428 7410 10456 7822
rect 10520 7585 10548 7890
rect 10506 7576 10562 7585
rect 10506 7511 10562 7520
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10416 7200 10468 7206
rect 10336 7160 10416 7188
rect 10416 7142 10468 7148
rect 10244 6990 10364 7018
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 9956 6384 10008 6390
rect 9784 6344 9956 6372
rect 9956 6326 10008 6332
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9876 5914 9904 6190
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9876 5778 9904 5850
rect 9864 5772 9916 5778
rect 9784 5732 9864 5760
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9784 5148 9812 5732
rect 9864 5714 9916 5720
rect 9864 5636 9916 5642
rect 9968 5624 9996 6326
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5914 10088 6258
rect 10244 6254 10272 6802
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10232 6112 10284 6118
rect 10336 6100 10364 6990
rect 10428 6338 10456 7142
rect 10520 6458 10548 7511
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10612 6361 10640 8026
rect 10598 6352 10654 6361
rect 10428 6310 10548 6338
rect 10284 6072 10364 6100
rect 10232 6054 10284 6060
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10152 5778 10180 6054
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 9916 5596 9996 5624
rect 9864 5578 9916 5584
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9692 5120 9812 5148
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9404 4616 9456 4622
rect 9402 4584 9404 4593
rect 9456 4584 9458 4593
rect 9402 4519 9458 4528
rect 9600 4486 9628 4694
rect 9692 4622 9720 5120
rect 9864 5024 9916 5030
rect 9784 4984 9864 5012
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9586 4176 9642 4185
rect 9416 4078 9444 4150
rect 9586 4111 9642 4120
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9036 2576 9088 2582
rect 9140 2553 9168 3674
rect 9324 3670 9352 4014
rect 9600 3942 9628 4111
rect 9692 4060 9720 4558
rect 9784 4282 9812 4984
rect 9864 4966 9916 4972
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10244 4321 10272 6054
rect 10322 5672 10378 5681
rect 10322 5607 10378 5616
rect 10336 4826 10364 5607
rect 10414 4856 10470 4865
rect 10324 4820 10376 4826
rect 10414 4791 10470 4800
rect 10324 4762 10376 4768
rect 10230 4312 10286 4321
rect 9772 4276 9824 4282
rect 10336 4282 10364 4762
rect 10230 4247 10286 4256
rect 10324 4276 10376 4282
rect 9772 4218 9824 4224
rect 9956 4072 10008 4078
rect 9692 4032 9956 4060
rect 9956 4014 10008 4020
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9770 3768 9826 3777
rect 9770 3703 9826 3712
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9692 3058 9720 3606
rect 9784 3505 9812 3703
rect 10244 3602 10272 4247
rect 10324 4218 10376 4224
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3738 10364 3878
rect 10428 3777 10456 4791
rect 10414 3768 10470 3777
rect 10324 3732 10376 3738
rect 10414 3703 10470 3712
rect 10324 3674 10376 3680
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 9770 3496 9826 3505
rect 10336 3482 10364 3674
rect 10428 3602 10456 3703
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10520 3534 10548 6310
rect 10598 6287 10654 6296
rect 10598 6216 10654 6225
rect 10598 6151 10600 6160
rect 10652 6151 10654 6160
rect 10600 6122 10652 6128
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10612 5273 10640 5306
rect 10598 5264 10654 5273
rect 10704 5234 10732 8298
rect 10796 5370 10824 13330
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10980 11762 11008 12174
rect 11150 12064 11206 12073
rect 11150 11999 11206 12008
rect 11058 11792 11114 11801
rect 10968 11756 11020 11762
rect 11058 11727 11060 11736
rect 10968 11698 11020 11704
rect 11112 11727 11114 11736
rect 11060 11698 11112 11704
rect 10980 11286 11008 11698
rect 11058 11656 11114 11665
rect 11058 11591 11114 11600
rect 11072 11558 11100 11591
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 11354 11100 11494
rect 11164 11354 11192 11999
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 11164 11218 11192 11290
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 10876 10192 10928 10198
rect 10874 10160 10876 10169
rect 10928 10160 10930 10169
rect 10874 10095 10930 10104
rect 11256 10062 11284 11494
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11348 10742 11376 11086
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11348 10606 11376 10678
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11440 10112 11468 14418
rect 13280 14278 13308 14554
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11520 10464 11572 10470
rect 11624 10441 11652 10542
rect 11520 10406 11572 10412
rect 11610 10432 11666 10441
rect 11532 10266 11560 10406
rect 11610 10367 11666 10376
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11520 10124 11572 10130
rect 11440 10084 11520 10112
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10888 8838 10916 9386
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10888 8401 10916 8774
rect 10874 8392 10930 8401
rect 10874 8327 10930 8336
rect 10980 7834 11008 9386
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8498 11100 8910
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11058 8392 11114 8401
rect 11058 8327 11114 8336
rect 11072 7886 11100 8327
rect 10888 7806 11008 7834
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10888 5710 10916 7806
rect 10968 7744 11020 7750
rect 10966 7712 10968 7721
rect 11060 7744 11112 7750
rect 11020 7712 11022 7721
rect 11060 7686 11112 7692
rect 10966 7647 11022 7656
rect 11072 7562 11100 7686
rect 10980 7534 11100 7562
rect 10980 6254 11008 7534
rect 11060 7472 11112 7478
rect 11164 7460 11192 8978
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 7546 11284 8230
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11112 7432 11192 7460
rect 11348 7449 11376 9658
rect 11440 9654 11468 10084
rect 11520 10066 11572 10072
rect 11428 9648 11480 9654
rect 11428 9590 11480 9596
rect 11610 9616 11666 9625
rect 11610 9551 11666 9560
rect 11624 9518 11652 9551
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11440 8090 11468 8298
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11532 8022 11560 8434
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11334 7440 11390 7449
rect 11060 7414 11112 7420
rect 11334 7375 11390 7384
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11164 6934 11192 7210
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11152 6928 11204 6934
rect 11256 6905 11284 6938
rect 11152 6870 11204 6876
rect 11242 6896 11298 6905
rect 11348 6866 11376 7278
rect 11242 6831 11298 6840
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11164 6254 11192 6734
rect 11242 6352 11298 6361
rect 11242 6287 11298 6296
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 11072 5574 11100 6122
rect 11256 5914 11284 6287
rect 11348 6118 11376 6802
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11164 5642 11192 5850
rect 11256 5817 11284 5850
rect 11242 5808 11298 5817
rect 11242 5743 11298 5752
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10598 5199 10654 5208
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 11072 5166 11100 5510
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11256 4758 11284 5510
rect 11348 5166 11376 5646
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11440 5098 11468 7890
rect 11532 7002 11560 7958
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11532 6458 11560 6598
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11624 5914 11652 8230
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11520 5772 11572 5778
rect 11716 5760 11744 13466
rect 12728 13258 12756 13806
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 13096 12889 13124 13398
rect 13082 12880 13138 12889
rect 13082 12815 13138 12824
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 13188 12442 13216 13398
rect 13372 12986 13400 14214
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 12348 12368 12400 12374
rect 12346 12336 12348 12345
rect 12400 12336 12402 12345
rect 12346 12271 12402 12280
rect 12530 12336 12586 12345
rect 12530 12271 12586 12280
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11794 10296 11850 10305
rect 11794 10231 11850 10240
rect 11808 9178 11836 10231
rect 11900 9994 11928 10542
rect 11992 10538 12204 10554
rect 11992 10532 12216 10538
rect 11992 10526 12164 10532
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11992 9654 12020 10526
rect 12164 10474 12216 10480
rect 12070 10432 12126 10441
rect 12070 10367 12126 10376
rect 12084 10266 12112 10367
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12162 10160 12218 10169
rect 12162 10095 12218 10104
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 12084 9586 12112 9998
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12176 9518 12204 10095
rect 12268 9926 12296 12038
rect 12544 11898 12572 12271
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12622 11792 12678 11801
rect 12544 11736 12622 11744
rect 12544 11716 12624 11736
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10305 12480 10406
rect 12438 10296 12494 10305
rect 12438 10231 12494 10240
rect 12544 10146 12572 11716
rect 12676 11727 12678 11736
rect 12624 11698 12676 11704
rect 12624 10532 12676 10538
rect 12728 10520 12756 12174
rect 13188 11914 13216 12378
rect 13188 11886 13400 11914
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12820 11150 12848 11222
rect 12808 11144 12860 11150
rect 12912 11121 12940 11222
rect 12808 11086 12860 11092
rect 12898 11112 12954 11121
rect 13188 11082 13216 11698
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11354 13308 11494
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 12898 11047 12954 11056
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13188 10606 13216 11018
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 12676 10492 12756 10520
rect 12624 10474 12676 10480
rect 12728 10248 12756 10492
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12728 10220 12940 10248
rect 12360 10130 12572 10146
rect 12348 10124 12572 10130
rect 12400 10118 12572 10124
rect 12808 10124 12860 10130
rect 12348 10066 12400 10072
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11900 8838 11928 9386
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 9178 12020 9318
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11808 8650 11836 8774
rect 11808 8622 11928 8650
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11520 5714 11572 5720
rect 11624 5732 11744 5760
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 10692 4616 10744 4622
rect 10612 4576 10692 4604
rect 10612 4010 10640 4576
rect 10692 4558 10744 4564
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 10874 4176 10930 4185
rect 10874 4111 10930 4120
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10508 3528 10560 3534
rect 10336 3454 10456 3482
rect 10508 3470 10560 3476
rect 9770 3431 9826 3440
rect 9784 3398 9812 3431
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 10336 3058 10364 3334
rect 10428 3194 10456 3454
rect 10520 3369 10548 3470
rect 10506 3360 10562 3369
rect 10506 3295 10562 3304
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10888 3126 10916 4111
rect 11072 4078 11100 4422
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 9036 2518 9088 2524
rect 9126 2544 9182 2553
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 8576 2508 8628 2514
rect 9126 2479 9182 2488
rect 8576 2450 8628 2456
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7576 800 7604 2314
rect 8496 800 8524 2314
rect 9416 800 9444 2994
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9968 2650 9996 2858
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 10428 898 10456 2926
rect 10888 2514 10916 3062
rect 11072 3058 11100 4014
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10888 2310 10916 2450
rect 11072 2446 11100 2994
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11164 2378 11192 4422
rect 11256 3534 11284 4694
rect 11532 3534 11560 5714
rect 11624 4826 11652 5732
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11612 4208 11664 4214
rect 11610 4176 11612 4185
rect 11664 4176 11666 4185
rect 11610 4111 11666 4120
rect 11244 3528 11296 3534
rect 11520 3528 11572 3534
rect 11296 3476 11376 3482
rect 11244 3470 11376 3476
rect 11520 3470 11572 3476
rect 11256 3454 11376 3470
rect 11348 2938 11376 3454
rect 11520 2984 11572 2990
rect 11348 2932 11520 2938
rect 11348 2926 11572 2932
rect 11348 2910 11560 2926
rect 11242 2816 11298 2825
rect 11242 2751 11298 2760
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10336 870 10456 898
rect 10336 800 10364 870
rect 11256 800 11284 2751
rect 11348 2446 11376 2910
rect 11426 2680 11482 2689
rect 11716 2650 11744 4966
rect 11808 2990 11836 8502
rect 11900 4078 11928 8622
rect 12268 8498 12296 9658
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12360 9178 12388 9318
rect 12452 9217 12480 10118
rect 12636 10084 12808 10112
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12438 9208 12494 9217
rect 12348 9172 12400 9178
rect 12438 9143 12494 9152
rect 12348 9114 12400 9120
rect 12360 8945 12388 9114
rect 12544 9110 12572 9998
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12532 8968 12584 8974
rect 12346 8936 12402 8945
rect 12346 8871 12402 8880
rect 12530 8936 12532 8945
rect 12584 8936 12586 8945
rect 12530 8871 12586 8880
rect 12438 8800 12494 8809
rect 12438 8735 12494 8744
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 11992 6186 12020 8434
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12070 7440 12126 7449
rect 12070 7375 12126 7384
rect 12084 7002 12112 7375
rect 12360 7274 12388 7822
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12176 6934 12204 7142
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12268 6746 12296 7142
rect 12084 6718 12296 6746
rect 12084 6662 12112 6718
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 11992 5409 12020 6122
rect 12084 5846 12112 6122
rect 12176 5914 12204 6598
rect 12452 6458 12480 8735
rect 12544 8362 12572 8871
rect 12636 8634 12664 10084
rect 12808 10066 12860 10072
rect 12912 9994 12940 10220
rect 13280 10062 13308 10950
rect 12992 10056 13044 10062
rect 13268 10056 13320 10062
rect 13044 10016 13268 10044
rect 12992 9998 13044 10004
rect 13268 9998 13320 10004
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 8974 12756 9454
rect 12912 9450 12940 9930
rect 13280 9897 13308 9998
rect 13266 9888 13322 9897
rect 13266 9823 13322 9832
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13174 9072 13230 9081
rect 13174 9007 13176 9016
rect 13228 9007 13230 9016
rect 13176 8978 13228 8984
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12440 6452 12492 6458
rect 12268 6412 12440 6440
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 11978 5400 12034 5409
rect 11978 5335 12034 5344
rect 12084 5166 12112 5782
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12176 5012 12204 5510
rect 12084 4984 12204 5012
rect 12084 4282 12112 4984
rect 12268 4672 12296 6412
rect 12440 6394 12492 6400
rect 12544 6225 12572 7414
rect 12636 6254 12664 8570
rect 12728 8090 12756 8910
rect 13372 8838 13400 11886
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7342 12848 7686
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12624 6248 12676 6254
rect 12530 6216 12586 6225
rect 12624 6190 12676 6196
rect 12820 6186 12848 6598
rect 13096 6458 13124 6734
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12530 6151 12586 6160
rect 12808 6180 12860 6186
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12360 5710 12388 6054
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12452 5030 12480 5714
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12176 4644 12296 4672
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11992 3670 12020 4218
rect 11980 3664 12032 3670
rect 12084 3652 12112 4218
rect 12176 3754 12204 4644
rect 12254 4584 12310 4593
rect 12452 4570 12480 4694
rect 12254 4519 12256 4528
rect 12308 4519 12310 4528
rect 12360 4542 12480 4570
rect 12256 4490 12308 4496
rect 12360 4282 12388 4542
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12176 3726 12296 3754
rect 12164 3664 12216 3670
rect 12084 3624 12164 3652
rect 11980 3606 12032 3612
rect 12164 3606 12216 3612
rect 12268 3126 12296 3726
rect 12256 3120 12308 3126
rect 12452 3074 12480 4422
rect 12256 3062 12308 3068
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 12360 3046 12480 3074
rect 12544 3058 12572 6151
rect 12808 6122 12860 6128
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12636 4865 12664 6054
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 5370 12756 5714
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12622 4856 12678 4865
rect 12622 4791 12678 4800
rect 12624 4752 12676 4758
rect 12622 4720 12624 4729
rect 12676 4720 12678 4729
rect 12622 4655 12678 4664
rect 12728 4622 12756 5306
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12806 4584 12862 4593
rect 12806 4519 12862 4528
rect 12622 4448 12678 4457
rect 12622 4383 12678 4392
rect 12636 3942 12664 4383
rect 12820 4282 12848 4519
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13084 4208 13136 4214
rect 13082 4176 13084 4185
rect 13136 4176 13138 4185
rect 13082 4111 13138 4120
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12898 3632 12954 3641
rect 12898 3567 12900 3576
rect 12952 3567 12954 3576
rect 12900 3538 12952 3544
rect 12532 3052 12584 3058
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11900 2825 11928 2994
rect 12360 2990 12388 3046
rect 12532 2994 12584 3000
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 11886 2816 11942 2825
rect 11886 2751 11942 2760
rect 12544 2650 12572 2994
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 11426 2615 11428 2624
rect 11480 2615 11482 2624
rect 11704 2644 11756 2650
rect 11428 2586 11480 2592
rect 11704 2586 11756 2592
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11440 2310 11468 2586
rect 13188 2514 13216 8502
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13266 7848 13322 7857
rect 13266 7783 13322 7792
rect 13280 7002 13308 7783
rect 13372 7290 13400 7890
rect 13464 7478 13492 14719
rect 14384 14550 14412 16400
rect 16578 16400 16634 17200
rect 18418 16824 18474 16833
rect 18418 16759 18474 16768
rect 16486 16351 16542 16360
rect 14646 16008 14702 16017
rect 14646 15943 14702 15952
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14384 13938 14412 14486
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13648 13734 13676 13806
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13530 13676 13670
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13556 10305 13584 11630
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13542 10296 13598 10305
rect 13542 10231 13598 10240
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13372 7262 13492 7290
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13372 5914 13400 7142
rect 13464 6254 13492 7262
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13556 6100 13584 9687
rect 13648 9042 13676 11494
rect 13740 11150 13768 12922
rect 13832 12850 13860 13330
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12170 13860 12786
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13924 11778 13952 12854
rect 14476 12850 14504 13126
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14016 11898 14044 12582
rect 14108 12442 14136 12582
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14200 12374 14228 12786
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14384 12442 14412 12718
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 14384 11830 14412 12242
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14372 11824 14424 11830
rect 13924 11750 14136 11778
rect 14372 11766 14424 11772
rect 14004 11620 14056 11626
rect 14004 11562 14056 11568
rect 14016 11354 14044 11562
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13728 11144 13780 11150
rect 13832 11121 13860 11290
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13728 11086 13780 11092
rect 13818 11112 13874 11121
rect 13740 10538 13768 11086
rect 13818 11047 13874 11056
rect 13832 11014 13860 11047
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13924 10674 13952 11154
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10198 13860 10406
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 13924 10010 13952 10134
rect 13740 9982 13952 10010
rect 13740 9110 13768 9982
rect 13910 9888 13966 9897
rect 13910 9823 13966 9832
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13636 8832 13688 8838
rect 13740 8820 13768 9046
rect 13688 8792 13768 8820
rect 13820 8832 13872 8838
rect 13636 8774 13688 8780
rect 13820 8774 13872 8780
rect 13648 8537 13676 8774
rect 13634 8528 13690 8537
rect 13634 8463 13690 8472
rect 13832 7954 13860 8774
rect 13924 8616 13952 9823
rect 14016 9654 14044 11086
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 13924 8588 14044 8616
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13924 7954 13952 8434
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 7002 13676 7142
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13740 6458 13768 7210
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13832 6322 13860 6666
rect 13924 6662 13952 7346
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13924 6458 13952 6598
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13464 6072 13584 6100
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 3534 13308 4966
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13372 4146 13400 4490
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13464 2582 13492 6072
rect 13740 5896 13768 6190
rect 13832 5914 13860 6258
rect 13648 5868 13768 5896
rect 13820 5908 13872 5914
rect 13648 5778 13676 5868
rect 13820 5850 13872 5856
rect 13726 5808 13782 5817
rect 13636 5772 13688 5778
rect 13726 5743 13782 5752
rect 13912 5772 13964 5778
rect 13636 5714 13688 5720
rect 13542 5400 13598 5409
rect 13542 5335 13598 5344
rect 13556 5302 13584 5335
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 13648 5234 13676 5714
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13556 4622 13584 4966
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13556 4010 13584 4422
rect 13648 4078 13676 5034
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13740 4026 13768 5743
rect 13912 5714 13964 5720
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 4486 13860 5510
rect 13924 5166 13952 5714
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 14016 4826 14044 8588
rect 14108 7426 14136 11750
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14188 9648 14240 9654
rect 14186 9616 14188 9625
rect 14240 9616 14242 9625
rect 14186 9551 14242 9560
rect 14292 9518 14320 10542
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14292 9110 14320 9454
rect 14280 9104 14332 9110
rect 14280 9046 14332 9052
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8566 14228 8774
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14384 8378 14412 11766
rect 14476 11336 14504 12038
rect 14568 11694 14596 13262
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14660 11354 14688 15943
rect 14738 15600 14794 15609
rect 14738 15535 14794 15544
rect 14752 14006 14780 15535
rect 16394 15192 16450 15201
rect 16394 15127 16450 15136
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14752 11762 14780 13942
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14936 12238 14964 12650
rect 15028 12306 15056 12718
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14648 11348 14700 11354
rect 14476 11308 14648 11336
rect 14568 10130 14596 11308
rect 14648 11290 14700 11296
rect 14844 11082 14872 12038
rect 14936 11762 14964 12174
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14922 11656 14978 11665
rect 14922 11591 14978 11600
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14646 10296 14702 10305
rect 14646 10231 14702 10240
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14660 9042 14688 10231
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9518 14780 9862
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14292 8350 14412 8378
rect 14200 7546 14228 8298
rect 14292 7750 14320 8350
rect 14476 8294 14504 8842
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14568 8498 14596 8774
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14292 7426 14320 7686
rect 14384 7546 14412 8230
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14108 7398 14228 7426
rect 14292 7398 14412 7426
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14108 5914 14136 6802
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14004 4820 14056 4826
rect 14056 4780 14136 4808
rect 14004 4762 14056 4768
rect 14108 4690 14136 4780
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13924 4321 13952 4558
rect 13910 4312 13966 4321
rect 14016 4282 14044 4626
rect 13910 4247 13966 4256
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 13912 4072 13964 4078
rect 13910 4040 13912 4049
rect 14004 4072 14056 4078
rect 13964 4040 13966 4049
rect 13544 4004 13596 4010
rect 13740 3998 13910 4026
rect 14004 4014 14056 4020
rect 13910 3975 13966 3984
rect 13544 3946 13596 3952
rect 13924 3915 13952 3975
rect 14016 3942 14044 4014
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14108 3670 14136 4082
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3058 13676 3334
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 14016 2650 14044 3130
rect 14200 2990 14228 7398
rect 14384 6934 14412 7398
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 6662 14320 6734
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14292 5642 14320 6598
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14292 4622 14320 5102
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14384 3126 14412 6122
rect 14476 6118 14504 8230
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7206 14596 7686
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 6905 14596 7142
rect 14554 6896 14610 6905
rect 14554 6831 14610 6840
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14568 5794 14596 6831
rect 14660 6798 14688 8978
rect 14752 8906 14780 9454
rect 14832 8968 14884 8974
rect 14936 8956 14964 11591
rect 15028 11354 15056 12242
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15212 11898 15240 12174
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15028 11150 15056 11290
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15028 10606 15056 11086
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15120 10266 15148 11154
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 15028 9625 15056 9930
rect 15014 9616 15070 9625
rect 15014 9551 15070 9560
rect 14884 8928 14964 8956
rect 14832 8910 14884 8916
rect 14740 8900 14792 8906
rect 14740 8842 14792 8848
rect 14738 8800 14794 8809
rect 14738 8735 14794 8744
rect 14752 7750 14780 8735
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14660 6662 14688 6734
rect 14844 6730 14872 8910
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14936 8022 14964 8298
rect 14924 8016 14976 8022
rect 14924 7958 14976 7964
rect 14936 7750 14964 7958
rect 14924 7744 14976 7750
rect 14922 7712 14924 7721
rect 14976 7712 14978 7721
rect 14922 7647 14978 7656
rect 15028 7478 15056 9551
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15120 8498 15148 9318
rect 15212 9178 15240 9454
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15304 8922 15332 14350
rect 16212 14272 16264 14278
rect 16210 14240 16212 14249
rect 16264 14240 16266 14249
rect 15782 14172 16078 14192
rect 16210 14175 16266 14184
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16040 13802 16068 13942
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15382 12880 15438 12889
rect 15382 12815 15438 12824
rect 15396 12170 15424 12815
rect 16304 12708 16356 12714
rect 16304 12650 16356 12656
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 15948 12345 15976 12582
rect 16132 12442 16160 12582
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 15934 12336 15990 12345
rect 15934 12271 15990 12280
rect 15384 12164 15436 12170
rect 15436 12124 15516 12152
rect 15384 12106 15436 12112
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 9178 15424 9862
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15488 9058 15516 12124
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 16132 11694 16160 12038
rect 16224 11762 16252 12378
rect 16316 11898 16344 12650
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16120 11688 16172 11694
rect 16408 11642 16436 15127
rect 16120 11630 16172 11636
rect 16224 11614 16436 11642
rect 16118 11520 16174 11529
rect 16118 11455 16174 11464
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15580 10470 15608 11154
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15212 8894 15332 8922
rect 15396 9030 15516 9058
rect 15396 8906 15424 9030
rect 15580 8974 15608 10406
rect 16040 10198 16068 10406
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15672 9722 15700 10066
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15764 9382 15792 9590
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15384 8900 15436 8906
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 15028 6798 15056 7414
rect 15120 7410 15148 8434
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 15028 6390 15056 6734
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 15028 6186 15056 6326
rect 15016 6180 15068 6186
rect 15016 6122 15068 6128
rect 14568 5766 14688 5794
rect 14556 5704 14608 5710
rect 14554 5672 14556 5681
rect 14608 5672 14610 5681
rect 14554 5607 14610 5616
rect 14660 4486 14688 5766
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15028 5234 15056 5646
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14476 4185 14504 4218
rect 14462 4176 14518 4185
rect 15028 4146 15056 5170
rect 14462 4111 14518 4120
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 14646 4040 14702 4049
rect 14646 3975 14702 3984
rect 14660 3738 14688 3975
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 15028 3466 15056 4082
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 12268 1306 12296 2382
rect 12176 1278 12296 1306
rect 12176 800 12204 1278
rect 13096 800 13124 2382
rect 13924 800 13952 2382
rect 14844 800 14872 2858
rect 14936 2650 14964 2858
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15212 1442 15240 8894
rect 15384 8842 15436 8848
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15304 2514 15332 8774
rect 15396 8362 15424 8842
rect 15488 8838 15516 8910
rect 15476 8832 15528 8838
rect 16040 8820 16068 9114
rect 16132 9110 16160 11455
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16040 8792 16160 8820
rect 15476 8774 15528 8780
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15580 7750 15608 8434
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15474 7576 15530 7585
rect 15474 7511 15530 7520
rect 15488 7342 15516 7511
rect 15672 7410 15700 8502
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 7002 15424 7142
rect 16132 7002 16160 8792
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 15934 5264 15990 5273
rect 15934 5199 15990 5208
rect 15948 5166 15976 5199
rect 16224 5166 16252 11614
rect 16394 11384 16450 11393
rect 16394 11319 16450 11328
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 7449 16344 9862
rect 16408 9178 16436 11319
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16408 8430 16436 8978
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16302 7440 16358 7449
rect 16408 7410 16436 7890
rect 16500 7546 16528 16351
rect 16592 14074 16620 16400
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16776 12442 16804 12786
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16592 11529 16620 11766
rect 16684 11762 16712 12310
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16578 11520 16634 11529
rect 16578 11455 16634 11464
rect 16684 11354 16712 11698
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16776 11014 16804 11494
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16592 9994 16620 10474
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 10198 16712 10406
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 16592 9586 16620 9930
rect 16684 9722 16712 9998
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 9042 16712 9318
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16580 8832 16632 8838
rect 16578 8800 16580 8809
rect 16632 8800 16634 8809
rect 16578 8735 16634 8744
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16684 8090 16712 8298
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16302 7375 16358 7384
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16500 7342 16528 7482
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15856 4826 15884 4966
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15396 3369 15424 3878
rect 15382 3360 15438 3369
rect 15382 3295 15438 3304
rect 15396 2990 15424 3295
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 16776 2650 16804 10950
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 16868 2446 16896 13874
rect 18064 13870 18092 14554
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 16948 13456 17000 13462
rect 16948 13398 17000 13404
rect 16960 12986 16988 13398
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17144 11898 17172 12582
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 16960 11218 16988 11562
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17236 11354 17264 11494
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16960 10441 16988 11154
rect 16946 10432 17002 10441
rect 16946 10367 17002 10376
rect 17328 10266 17356 11494
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17144 10033 17172 10066
rect 17130 10024 17186 10033
rect 17130 9959 17132 9968
rect 17184 9959 17186 9968
rect 17132 9930 17184 9936
rect 17420 9625 17448 12582
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17512 10810 17540 11698
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17512 10198 17540 10746
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17406 9616 17462 9625
rect 17224 9580 17276 9586
rect 17406 9551 17462 9560
rect 17224 9522 17276 9528
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17144 8945 17172 9318
rect 17236 9110 17264 9522
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17130 8936 17186 8945
rect 17130 8871 17186 8880
rect 17236 8634 17264 9046
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16960 3641 16988 6666
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 16946 3632 17002 3641
rect 16946 3567 17002 3576
rect 16960 2582 16988 3567
rect 17132 3528 17184 3534
rect 17130 3496 17132 3505
rect 17184 3496 17186 3505
rect 17130 3431 17186 3440
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16316 2106 16344 2246
rect 16304 2100 16356 2106
rect 16304 2042 16356 2048
rect 15212 1414 15792 1442
rect 15764 800 15792 1414
rect 16684 800 16712 2382
rect 17052 1465 17080 2790
rect 17236 2446 17264 6054
rect 17512 5778 17540 6598
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17420 3194 17448 4694
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17420 2990 17448 3130
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 1873 17356 2246
rect 17314 1864 17370 1873
rect 17314 1799 17370 1808
rect 17038 1456 17094 1465
rect 17038 1391 17094 1400
rect 17604 800 17632 13670
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17696 12306 17724 12786
rect 18050 12608 18106 12617
rect 18050 12543 18106 12552
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17696 12170 17724 12242
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17788 11898 17816 12174
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17788 11665 17816 11834
rect 17774 11656 17830 11665
rect 17774 11591 17830 11600
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17684 10736 17736 10742
rect 17684 10678 17736 10684
rect 17696 10266 17724 10678
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17696 8430 17724 10066
rect 17788 10062 17816 11086
rect 17880 10266 17908 11154
rect 17958 11112 18014 11121
rect 17958 11047 18014 11056
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17788 9466 17816 9998
rect 17788 9438 17908 9466
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9217 17816 9318
rect 17774 9208 17830 9217
rect 17880 9178 17908 9438
rect 17774 9143 17830 9152
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17880 8265 17908 8502
rect 17866 8256 17922 8265
rect 17866 8191 17922 8200
rect 17972 7342 18000 11047
rect 18064 9926 18092 12543
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18156 11898 18184 12242
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18156 10305 18184 11834
rect 18432 11354 18460 16759
rect 18786 16400 18842 17200
rect 18800 14550 18828 16400
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18142 10296 18198 10305
rect 18142 10231 18198 10240
rect 18432 10169 18460 11290
rect 18418 10160 18474 10169
rect 18418 10095 18474 10104
rect 18142 10024 18198 10033
rect 18142 9959 18198 9968
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18156 9518 18184 9959
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18050 7848 18106 7857
rect 18050 7783 18052 7792
rect 18104 7783 18106 7792
rect 18052 7754 18104 7760
rect 18236 7472 18288 7478
rect 18234 7440 18236 7449
rect 18288 7440 18290 7449
rect 18234 7375 18290 7384
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 18052 6656 18104 6662
rect 18050 6624 18052 6633
rect 18104 6624 18106 6633
rect 18050 6559 18106 6568
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 18234 6216 18290 6225
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17880 5273 17908 5510
rect 17866 5264 17922 5273
rect 17866 5199 17922 5208
rect 17972 4282 18000 6190
rect 18234 6151 18290 6160
rect 18248 6118 18276 6151
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18248 5370 18276 5714
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18340 4865 18368 8774
rect 18418 7032 18474 7041
rect 18418 6967 18474 6976
rect 18432 6730 18460 6967
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 18418 5672 18474 5681
rect 18418 5607 18420 5616
rect 18472 5607 18474 5616
rect 18420 5578 18472 5584
rect 18326 4856 18382 4865
rect 18326 4791 18382 4800
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18052 4480 18104 4486
rect 18050 4448 18052 4457
rect 18104 4448 18106 4457
rect 18050 4383 18106 4392
rect 18432 4282 18460 4558
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 18234 4040 18290 4049
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17696 3641 17724 3674
rect 17682 3632 17738 3641
rect 17682 3567 17738 3576
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17684 2304 17736 2310
rect 17788 2281 17816 2790
rect 17880 2689 17908 3334
rect 17972 2990 18000 4014
rect 18234 3975 18290 3984
rect 18248 3942 18276 3975
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18432 3602 18460 4218
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18432 3233 18460 3334
rect 18418 3224 18474 3233
rect 18418 3159 18474 3168
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 17866 2680 17922 2689
rect 17866 2615 17922 2624
rect 17868 2304 17920 2310
rect 17684 2246 17736 2252
rect 17774 2272 17830 2281
rect 17696 1057 17724 2246
rect 17868 2246 17920 2252
rect 17774 2207 17830 2216
rect 17682 1048 17738 1057
rect 17682 983 17738 992
rect 3422 640 3478 649
rect 3422 575 3478 584
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15750 0 15806 800
rect 16670 0 16726 800
rect 17590 0 17646 800
rect 17880 241 17908 2246
rect 18248 649 18276 2790
rect 18524 800 18552 13670
rect 18970 13424 19026 13433
rect 18970 13359 19026 13368
rect 18984 10742 19012 13359
rect 18972 10736 19024 10742
rect 18972 10678 19024 10684
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19444 800 19472 2858
rect 18234 640 18290 649
rect 18234 575 18290 584
rect 17866 232 17922 241
rect 17866 167 17922 176
rect 18510 0 18566 800
rect 19430 0 19486 800
<< via2 >>
rect 3238 16768 3294 16824
rect 1490 15952 1546 16008
rect 2134 14728 2190 14784
rect 2594 13504 2650 13560
rect 1582 6976 1638 7032
rect 1398 3848 1454 3904
rect 1582 3884 1584 3904
rect 1584 3884 1636 3904
rect 1636 3884 1638 3904
rect 1582 3848 1638 3884
rect 1582 2488 1638 2544
rect 2870 11328 2926 11384
rect 2778 11192 2834 11248
rect 2594 9560 2650 9616
rect 3422 16360 3478 16416
rect 4986 15136 5042 15192
rect 4066 14356 4068 14376
rect 4068 14356 4120 14376
rect 4120 14356 4122 14376
rect 4066 14320 4122 14356
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3790 13912 3846 13968
rect 3698 13096 3754 13152
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3974 12316 3976 12336
rect 3976 12316 4028 12336
rect 4028 12316 4030 12336
rect 3974 12280 4030 12316
rect 3606 12144 3662 12200
rect 3422 11872 3478 11928
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3514 11056 3570 11112
rect 1858 7656 1914 7712
rect 2502 7792 2558 7848
rect 1766 6840 1822 6896
rect 1950 6840 2006 6896
rect 2042 4936 2098 4992
rect 1766 4120 1822 4176
rect 2134 4020 2136 4040
rect 2136 4020 2188 4040
rect 2188 4020 2190 4040
rect 2134 3984 2190 4020
rect 1858 3440 1914 3496
rect 2318 3848 2374 3904
rect 2962 8880 3018 8936
rect 2778 6432 2834 6488
rect 2778 4664 2834 4720
rect 2226 2624 2282 2680
rect 3238 10376 3294 10432
rect 3698 10956 3700 10976
rect 3700 10956 3752 10976
rect 3752 10956 3754 10976
rect 3698 10920 3754 10956
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 3606 10104 3662 10160
rect 4158 10104 4214 10160
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 3514 9696 3570 9752
rect 3422 8880 3478 8936
rect 3422 8508 3424 8528
rect 3424 8508 3476 8528
rect 3476 8508 3478 8528
rect 3422 8472 3478 8508
rect 4158 9324 4160 9344
rect 4160 9324 4212 9344
rect 4212 9324 4214 9344
rect 4158 9288 4214 9324
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 3974 8372 3976 8392
rect 3976 8372 4028 8392
rect 4028 8372 4030 8392
rect 3974 8336 4030 8372
rect 4342 10240 4398 10296
rect 4894 10512 4950 10568
rect 4526 9560 4582 9616
rect 4526 9424 4582 9480
rect 4894 10376 4950 10432
rect 3790 8084 3846 8120
rect 3790 8064 3792 8084
rect 3792 8064 3844 8084
rect 3844 8064 3846 8084
rect 3698 7112 3754 7168
rect 3238 6024 3294 6080
rect 3698 5516 3700 5536
rect 3700 5516 3752 5536
rect 3752 5516 3754 5536
rect 3698 5480 3754 5516
rect 3146 5072 3202 5128
rect 2962 4256 3018 4312
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 4066 7248 4122 7304
rect 4434 6976 4490 7032
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 4434 4972 4436 4992
rect 4436 4972 4488 4992
rect 4488 4972 4490 4992
rect 4434 4936 4490 4972
rect 4526 4664 4582 4720
rect 1858 2216 1914 2272
rect 2870 3032 2926 3088
rect 2778 1808 2834 1864
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3882 4020 3884 4040
rect 3884 4020 3936 4040
rect 3936 4020 3938 4040
rect 3882 3984 3938 4020
rect 4342 4392 4398 4448
rect 3882 3460 3938 3496
rect 3882 3440 3884 3460
rect 3884 3440 3936 3460
rect 3936 3440 3938 3460
rect 4342 3440 4398 3496
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 3146 1400 3202 1456
rect 1398 176 1454 232
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 5446 10648 5502 10704
rect 6366 10260 6422 10296
rect 6366 10240 6368 10260
rect 6368 10240 6420 10260
rect 6420 10240 6422 10260
rect 6366 9968 6422 10024
rect 5998 7928 6054 7984
rect 5170 5208 5226 5264
rect 5446 4392 5502 4448
rect 6182 8744 6238 8800
rect 6274 8472 6330 8528
rect 6550 10412 6552 10432
rect 6552 10412 6604 10432
rect 6604 10412 6606 10432
rect 6550 10376 6606 10412
rect 6734 15544 6790 15600
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 7378 11056 7434 11112
rect 7562 11056 7618 11112
rect 5814 4120 5870 4176
rect 6826 9560 6882 9616
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 7470 9152 7526 9208
rect 7010 9016 7066 9072
rect 7286 9016 7342 9072
rect 7378 8608 7434 8664
rect 7010 8336 7066 8392
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6366 7112 6422 7168
rect 6366 6704 6422 6760
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 5998 3576 6054 3632
rect 6826 6316 6882 6352
rect 6826 6296 6828 6316
rect 6828 6296 6880 6316
rect 6880 6296 6882 6316
rect 6642 4936 6698 4992
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6918 5108 6920 5128
rect 6920 5108 6972 5128
rect 6972 5108 6974 5128
rect 7654 9152 7710 9208
rect 7470 7792 7526 7848
rect 6918 5072 6974 5108
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6918 4684 6974 4720
rect 6918 4664 6920 4684
rect 6920 4664 6972 4684
rect 6972 4664 6974 4684
rect 6642 3984 6698 4040
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 7654 6296 7710 6352
rect 7654 5072 7710 5128
rect 7562 4700 7564 4720
rect 7564 4700 7616 4720
rect 7616 4700 7618 4720
rect 7562 4664 7618 4700
rect 7746 4120 7802 4176
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 3790 992 3846 1048
rect 6918 2508 6974 2544
rect 6918 2488 6920 2508
rect 6920 2488 6972 2508
rect 6972 2488 6974 2508
rect 8298 11212 8354 11248
rect 8298 11192 8300 11212
rect 8300 11192 8352 11212
rect 8352 11192 8354 11212
rect 8206 10512 8262 10568
rect 8022 9968 8078 10024
rect 8022 9580 8078 9616
rect 8022 9560 8024 9580
rect 8024 9560 8076 9580
rect 8076 9560 8078 9580
rect 8574 9424 8630 9480
rect 8482 8744 8538 8800
rect 8482 4528 8538 4584
rect 8482 3984 8538 4040
rect 8758 12688 8814 12744
rect 13450 14728 13506 14784
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 10414 13776 10470 13832
rect 8758 8492 8814 8528
rect 8758 8472 8760 8492
rect 8760 8472 8812 8492
rect 8812 8472 8814 8492
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9494 12144 9550 12200
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 10138 11600 10194 11656
rect 9402 10124 9458 10160
rect 9402 10104 9404 10124
rect 9404 10104 9456 10124
rect 9456 10104 9458 10124
rect 8758 7928 8814 7984
rect 8666 5208 8722 5264
rect 8850 4392 8906 4448
rect 9310 7928 9366 7984
rect 9126 7248 9182 7304
rect 9126 6860 9182 6896
rect 9126 6840 9128 6860
rect 9128 6840 9180 6860
rect 9180 6840 9182 6860
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10138 8492 10194 8528
rect 10138 8472 10140 8492
rect 10140 8472 10192 8492
rect 10192 8472 10194 8492
rect 10046 7812 10102 7848
rect 10046 7792 10048 7812
rect 10048 7792 10100 7812
rect 10100 7792 10102 7812
rect 10690 11772 10692 11792
rect 10692 11772 10744 11792
rect 10744 11772 10746 11792
rect 10690 11736 10746 11772
rect 10322 9696 10378 9752
rect 10414 9016 10470 9072
rect 10690 9988 10746 10024
rect 10690 9968 10692 9988
rect 10692 9968 10744 9988
rect 10744 9968 10746 9988
rect 10598 8880 10654 8936
rect 10414 7928 10470 7984
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 10230 7520 10286 7576
rect 10506 7520 10562 7576
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9402 4564 9404 4584
rect 9404 4564 9456 4584
rect 9456 4564 9458 4584
rect 9402 4528 9458 4564
rect 9586 4120 9642 4176
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10322 5616 10378 5672
rect 10414 4800 10470 4856
rect 10230 4256 10286 4312
rect 9770 3712 9826 3768
rect 10414 3712 10470 3768
rect 9770 3440 9826 3496
rect 10598 6296 10654 6352
rect 10598 6180 10654 6216
rect 10598 6160 10600 6180
rect 10600 6160 10652 6180
rect 10652 6160 10654 6180
rect 10598 5208 10654 5264
rect 11150 12008 11206 12064
rect 11058 11756 11114 11792
rect 11058 11736 11060 11756
rect 11060 11736 11112 11756
rect 11112 11736 11114 11756
rect 11058 11600 11114 11656
rect 10874 10140 10876 10160
rect 10876 10140 10928 10160
rect 10928 10140 10930 10160
rect 10874 10104 10930 10140
rect 11610 10376 11666 10432
rect 10874 8336 10930 8392
rect 11058 8336 11114 8392
rect 10966 7692 10968 7712
rect 10968 7692 11020 7712
rect 11020 7692 11022 7712
rect 10966 7656 11022 7692
rect 11610 9560 11666 9616
rect 11334 7384 11390 7440
rect 11242 6840 11298 6896
rect 11242 6296 11298 6352
rect 11242 5752 11298 5808
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 13082 12824 13138 12880
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12346 12316 12348 12336
rect 12348 12316 12400 12336
rect 12400 12316 12402 12336
rect 12346 12280 12402 12316
rect 12530 12280 12586 12336
rect 11794 10240 11850 10296
rect 12070 10376 12126 10432
rect 12162 10104 12218 10160
rect 12622 11756 12678 11792
rect 12622 11736 12624 11756
rect 12624 11736 12676 11756
rect 12676 11736 12678 11756
rect 12438 10240 12494 10296
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12898 11056 12954 11112
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 10874 4120 10930 4176
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 10506 3304 10562 3360
rect 9126 2488 9182 2544
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 11610 4156 11612 4176
rect 11612 4156 11664 4176
rect 11664 4156 11666 4176
rect 11610 4120 11666 4156
rect 11242 2760 11298 2816
rect 11426 2644 11482 2680
rect 12438 9152 12494 9208
rect 12346 8880 12402 8936
rect 12530 8916 12532 8936
rect 12532 8916 12584 8936
rect 12584 8916 12586 8936
rect 12530 8880 12586 8916
rect 12438 8744 12494 8800
rect 12070 7384 12126 7440
rect 13266 9832 13322 9888
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 13174 9036 13230 9072
rect 13174 9016 13176 9036
rect 13176 9016 13228 9036
rect 13228 9016 13230 9036
rect 11978 5344 12034 5400
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 12530 6160 12586 6216
rect 12254 4548 12310 4584
rect 12254 4528 12256 4548
rect 12256 4528 12308 4548
rect 12308 4528 12310 4548
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12622 4800 12678 4856
rect 12622 4700 12624 4720
rect 12624 4700 12676 4720
rect 12676 4700 12678 4720
rect 12622 4664 12678 4700
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 12806 4528 12862 4584
rect 12622 4392 12678 4448
rect 13082 4156 13084 4176
rect 13084 4156 13136 4176
rect 13136 4156 13138 4176
rect 13082 4120 13138 4156
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12898 3596 12954 3632
rect 12898 3576 12900 3596
rect 12900 3576 12952 3596
rect 12952 3576 12954 3596
rect 11886 2760 11942 2816
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 11426 2624 11428 2644
rect 11428 2624 11480 2644
rect 11480 2624 11482 2644
rect 13266 7792 13322 7848
rect 16486 16360 16542 16416
rect 18418 16768 18474 16824
rect 14646 15952 14702 16008
rect 13542 10240 13598 10296
rect 13542 9696 13598 9752
rect 13818 11056 13874 11112
rect 13910 9832 13966 9888
rect 13634 8472 13690 8528
rect 13726 5752 13782 5808
rect 13542 5344 13598 5400
rect 14186 9596 14188 9616
rect 14188 9596 14240 9616
rect 14240 9596 14242 9616
rect 14186 9560 14242 9596
rect 14738 15544 14794 15600
rect 16394 15136 16450 15192
rect 14922 11600 14978 11656
rect 14646 10240 14702 10296
rect 13910 4256 13966 4312
rect 13910 4020 13912 4040
rect 13912 4020 13964 4040
rect 13964 4020 13966 4040
rect 13910 3984 13966 4020
rect 14554 6840 14610 6896
rect 15014 9560 15070 9616
rect 14738 8744 14794 8800
rect 14922 7692 14924 7712
rect 14924 7692 14976 7712
rect 14976 7692 14978 7712
rect 14922 7656 14978 7692
rect 16210 14220 16212 14240
rect 16212 14220 16264 14240
rect 16264 14220 16266 14240
rect 16210 14184 16266 14220
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15382 12824 15438 12880
rect 15934 12280 15990 12336
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 16118 11464 16174 11520
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 14554 5652 14556 5672
rect 14556 5652 14608 5672
rect 14608 5652 14610 5672
rect 14554 5616 14610 5652
rect 14462 4120 14518 4176
rect 14646 3984 14702 4040
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15474 7520 15530 7576
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15934 5208 15990 5264
rect 16394 11328 16450 11384
rect 16302 7384 16358 7440
rect 16578 11464 16634 11520
rect 16578 8780 16580 8800
rect 16580 8780 16632 8800
rect 16632 8780 16634 8800
rect 16578 8744 16634 8780
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15382 3304 15438 3360
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 16946 10376 17002 10432
rect 17130 9988 17186 10024
rect 17130 9968 17132 9988
rect 17132 9968 17184 9988
rect 17184 9968 17186 9988
rect 17406 9560 17462 9616
rect 17130 8880 17186 8936
rect 16946 3576 17002 3632
rect 17130 3476 17132 3496
rect 17132 3476 17184 3496
rect 17184 3476 17186 3496
rect 17130 3440 17186 3476
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 17314 1808 17370 1864
rect 17038 1400 17094 1456
rect 18050 12552 18106 12608
rect 17774 11600 17830 11656
rect 17958 11056 18014 11112
rect 17774 9152 17830 9208
rect 17866 8200 17922 8256
rect 18142 10240 18198 10296
rect 18418 10104 18474 10160
rect 18142 9968 18198 10024
rect 18050 7812 18106 7848
rect 18050 7792 18052 7812
rect 18052 7792 18104 7812
rect 18104 7792 18106 7812
rect 18234 7420 18236 7440
rect 18236 7420 18288 7440
rect 18288 7420 18290 7440
rect 18234 7384 18290 7420
rect 18050 6604 18052 6624
rect 18052 6604 18104 6624
rect 18104 6604 18106 6624
rect 18050 6568 18106 6604
rect 17866 5208 17922 5264
rect 18234 6160 18290 6216
rect 18418 6976 18474 7032
rect 18418 5636 18474 5672
rect 18418 5616 18420 5636
rect 18420 5616 18472 5636
rect 18472 5616 18474 5636
rect 18326 4800 18382 4856
rect 18050 4428 18052 4448
rect 18052 4428 18104 4448
rect 18104 4428 18106 4448
rect 18050 4392 18106 4428
rect 17682 3576 17738 3632
rect 18234 3984 18290 4040
rect 18418 3168 18474 3224
rect 17866 2624 17922 2680
rect 17774 2216 17830 2272
rect 17682 992 17738 1048
rect 3422 584 3478 640
rect 18970 13368 19026 13424
rect 18234 584 18290 640
rect 17866 176 17922 232
<< metal3 >>
rect 0 16826 800 16856
rect 3233 16826 3299 16829
rect 0 16824 3299 16826
rect 0 16768 3238 16824
rect 3294 16768 3299 16824
rect 0 16766 3299 16768
rect 0 16736 800 16766
rect 3233 16763 3299 16766
rect 18413 16826 18479 16829
rect 19200 16826 20000 16856
rect 18413 16824 20000 16826
rect 18413 16768 18418 16824
rect 18474 16768 20000 16824
rect 18413 16766 20000 16768
rect 18413 16763 18479 16766
rect 19200 16736 20000 16766
rect 0 16418 800 16448
rect 3417 16418 3483 16421
rect 0 16416 3483 16418
rect 0 16360 3422 16416
rect 3478 16360 3483 16416
rect 0 16358 3483 16360
rect 0 16328 800 16358
rect 3417 16355 3483 16358
rect 16481 16418 16547 16421
rect 19200 16418 20000 16448
rect 16481 16416 20000 16418
rect 16481 16360 16486 16416
rect 16542 16360 20000 16416
rect 16481 16358 20000 16360
rect 16481 16355 16547 16358
rect 19200 16328 20000 16358
rect 0 16010 800 16040
rect 1485 16010 1551 16013
rect 0 16008 1551 16010
rect 0 15952 1490 16008
rect 1546 15952 1551 16008
rect 0 15950 1551 15952
rect 0 15920 800 15950
rect 1485 15947 1551 15950
rect 14641 16010 14707 16013
rect 19200 16010 20000 16040
rect 14641 16008 20000 16010
rect 14641 15952 14646 16008
rect 14702 15952 20000 16008
rect 14641 15950 20000 15952
rect 14641 15947 14707 15950
rect 19200 15920 20000 15950
rect 0 15602 800 15632
rect 6729 15602 6795 15605
rect 0 15600 6795 15602
rect 0 15544 6734 15600
rect 6790 15544 6795 15600
rect 0 15542 6795 15544
rect 0 15512 800 15542
rect 6729 15539 6795 15542
rect 14733 15602 14799 15605
rect 19200 15602 20000 15632
rect 14733 15600 20000 15602
rect 14733 15544 14738 15600
rect 14794 15544 20000 15600
rect 14733 15542 20000 15544
rect 14733 15539 14799 15542
rect 19200 15512 20000 15542
rect 0 15194 800 15224
rect 4981 15194 5047 15197
rect 0 15192 5047 15194
rect 0 15136 4986 15192
rect 5042 15136 5047 15192
rect 0 15134 5047 15136
rect 0 15104 800 15134
rect 4981 15131 5047 15134
rect 16389 15194 16455 15197
rect 19200 15194 20000 15224
rect 16389 15192 20000 15194
rect 16389 15136 16394 15192
rect 16450 15136 20000 15192
rect 16389 15134 20000 15136
rect 16389 15131 16455 15134
rect 19200 15104 20000 15134
rect 0 14786 800 14816
rect 2129 14786 2195 14789
rect 0 14784 2195 14786
rect 0 14728 2134 14784
rect 2190 14728 2195 14784
rect 0 14726 2195 14728
rect 0 14696 800 14726
rect 2129 14723 2195 14726
rect 13445 14786 13511 14789
rect 19200 14786 20000 14816
rect 13445 14784 20000 14786
rect 13445 14728 13450 14784
rect 13506 14728 20000 14784
rect 13445 14726 20000 14728
rect 13445 14723 13511 14726
rect 6874 14720 7194 14721
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 19200 14696 20000 14726
rect 12805 14655 13125 14656
rect 0 14378 800 14408
rect 4061 14378 4127 14381
rect 0 14376 4127 14378
rect 0 14320 4066 14376
rect 4122 14320 4127 14376
rect 0 14318 4127 14320
rect 0 14288 800 14318
rect 4061 14315 4127 14318
rect 16205 14242 16271 14245
rect 19200 14242 20000 14272
rect 16205 14240 20000 14242
rect 16205 14184 16210 14240
rect 16266 14184 20000 14240
rect 16205 14182 20000 14184
rect 16205 14179 16271 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19200 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13970 800 14000
rect 3785 13970 3851 13973
rect 0 13968 3851 13970
rect 0 13912 3790 13968
rect 3846 13912 3851 13968
rect 0 13910 3851 13912
rect 0 13880 800 13910
rect 3785 13907 3851 13910
rect 10409 13834 10475 13837
rect 19200 13834 20000 13864
rect 10409 13832 20000 13834
rect 10409 13776 10414 13832
rect 10470 13776 20000 13832
rect 10409 13774 20000 13776
rect 10409 13771 10475 13774
rect 19200 13744 20000 13774
rect 6874 13632 7194 13633
rect 0 13562 800 13592
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 2589 13562 2655 13565
rect 0 13560 2655 13562
rect 0 13504 2594 13560
rect 2650 13504 2655 13560
rect 0 13502 2655 13504
rect 0 13472 800 13502
rect 2589 13499 2655 13502
rect 18965 13426 19031 13429
rect 19200 13426 20000 13456
rect 18965 13424 20000 13426
rect 18965 13368 18970 13424
rect 19026 13368 20000 13424
rect 18965 13366 20000 13368
rect 18965 13363 19031 13366
rect 19200 13336 20000 13366
rect 0 13154 800 13184
rect 3693 13154 3759 13157
rect 0 13152 3759 13154
rect 0 13096 3698 13152
rect 3754 13096 3759 13152
rect 0 13094 3759 13096
rect 0 13064 800 13094
rect 3693 13091 3759 13094
rect 3909 13088 4229 13089
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 19200 13018 20000 13048
rect 16208 12958 20000 13018
rect 13077 12882 13143 12885
rect 15377 12882 15443 12885
rect 16208 12882 16268 12958
rect 19200 12928 20000 12958
rect 13077 12880 16268 12882
rect 13077 12824 13082 12880
rect 13138 12824 15382 12880
rect 15438 12824 16268 12880
rect 13077 12822 16268 12824
rect 13077 12819 13143 12822
rect 15377 12819 15443 12822
rect 0 12746 800 12776
rect 8753 12746 8819 12749
rect 0 12744 8819 12746
rect 0 12688 8758 12744
rect 8814 12688 8819 12744
rect 0 12686 8819 12688
rect 0 12656 800 12686
rect 8753 12683 8819 12686
rect 18045 12610 18111 12613
rect 19200 12610 20000 12640
rect 18045 12608 20000 12610
rect 18045 12552 18050 12608
rect 18106 12552 20000 12608
rect 18045 12550 20000 12552
rect 18045 12547 18111 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 19200 12520 20000 12550
rect 12805 12479 13125 12480
rect 0 12338 800 12368
rect 3969 12338 4035 12341
rect 0 12336 4035 12338
rect 0 12280 3974 12336
rect 4030 12280 4035 12336
rect 0 12278 4035 12280
rect 0 12248 800 12278
rect 3969 12275 4035 12278
rect 12341 12338 12407 12341
rect 12525 12338 12591 12341
rect 12341 12336 12591 12338
rect 12341 12280 12346 12336
rect 12402 12280 12530 12336
rect 12586 12280 12591 12336
rect 12341 12278 12591 12280
rect 12341 12275 12407 12278
rect 12525 12275 12591 12278
rect 15510 12276 15516 12340
rect 15580 12338 15586 12340
rect 15929 12338 15995 12341
rect 15580 12336 15995 12338
rect 15580 12280 15934 12336
rect 15990 12280 15995 12336
rect 15580 12278 15995 12280
rect 15580 12276 15586 12278
rect 15929 12275 15995 12278
rect 3601 12202 3667 12205
rect 9489 12202 9555 12205
rect 19200 12202 20000 12232
rect 3601 12200 9555 12202
rect 3601 12144 3606 12200
rect 3662 12144 9494 12200
rect 9550 12144 9555 12200
rect 3601 12142 9555 12144
rect 3601 12139 3667 12142
rect 9489 12139 9555 12142
rect 14920 12142 20000 12202
rect 11145 12066 11211 12069
rect 14920 12066 14980 12142
rect 19200 12112 20000 12142
rect 11145 12064 14980 12066
rect 11145 12008 11150 12064
rect 11206 12008 14980 12064
rect 11145 12006 14980 12008
rect 11145 12003 11211 12006
rect 3909 12000 4229 12001
rect 0 11930 800 11960
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 3417 11930 3483 11933
rect 0 11928 3483 11930
rect 0 11872 3422 11928
rect 3478 11872 3483 11928
rect 0 11870 3483 11872
rect 0 11840 800 11870
rect 3417 11867 3483 11870
rect 10685 11794 10751 11797
rect 11053 11794 11119 11797
rect 10685 11792 11119 11794
rect 10685 11736 10690 11792
rect 10746 11736 11058 11792
rect 11114 11736 11119 11792
rect 10685 11734 11119 11736
rect 10685 11731 10751 11734
rect 11053 11731 11119 11734
rect 12617 11794 12683 11797
rect 19200 11794 20000 11824
rect 12617 11792 20000 11794
rect 12617 11736 12622 11792
rect 12678 11736 20000 11792
rect 12617 11734 20000 11736
rect 12617 11731 12683 11734
rect 19200 11704 20000 11734
rect 10133 11658 10199 11661
rect 11053 11658 11119 11661
rect 14917 11658 14983 11661
rect 17769 11658 17835 11661
rect 10133 11656 17835 11658
rect 10133 11600 10138 11656
rect 10194 11600 11058 11656
rect 11114 11600 14922 11656
rect 14978 11600 17774 11656
rect 17830 11600 17835 11656
rect 10133 11598 17835 11600
rect 10133 11595 10199 11598
rect 11053 11595 11119 11598
rect 14917 11595 14983 11598
rect 17769 11595 17835 11598
rect 16113 11522 16179 11525
rect 16573 11522 16639 11525
rect 16113 11520 16639 11522
rect 16113 11464 16118 11520
rect 16174 11464 16578 11520
rect 16634 11464 16639 11520
rect 16113 11462 16639 11464
rect 16113 11459 16179 11462
rect 16573 11459 16639 11462
rect 6874 11456 7194 11457
rect 0 11386 800 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 2865 11386 2931 11389
rect 0 11384 2931 11386
rect 0 11328 2870 11384
rect 2926 11328 2931 11384
rect 0 11326 2931 11328
rect 0 11296 800 11326
rect 2865 11323 2931 11326
rect 16389 11386 16455 11389
rect 16389 11384 16498 11386
rect 16389 11328 16394 11384
rect 16450 11328 16498 11384
rect 16389 11323 16498 11328
rect 2773 11250 2839 11253
rect 8293 11250 8359 11253
rect 2773 11248 8359 11250
rect 2773 11192 2778 11248
rect 2834 11192 8298 11248
rect 8354 11192 8359 11248
rect 2773 11190 8359 11192
rect 16438 11250 16498 11323
rect 19200 11250 20000 11280
rect 16438 11190 20000 11250
rect 2773 11187 2839 11190
rect 8293 11187 8359 11190
rect 19200 11160 20000 11190
rect 3509 11114 3575 11117
rect 7373 11114 7439 11117
rect 3509 11112 7439 11114
rect 3509 11056 3514 11112
rect 3570 11056 7378 11112
rect 7434 11056 7439 11112
rect 3509 11054 7439 11056
rect 3509 11051 3575 11054
rect 7373 11051 7439 11054
rect 7557 11116 7623 11117
rect 7557 11112 7604 11116
rect 7668 11114 7674 11116
rect 12893 11114 12959 11117
rect 7668 11112 12959 11114
rect 7557 11056 7562 11112
rect 7668 11056 12898 11112
rect 12954 11056 12959 11112
rect 7557 11052 7604 11056
rect 7668 11054 12959 11056
rect 7668 11052 7674 11054
rect 7557 11051 7623 11052
rect 12893 11051 12959 11054
rect 13813 11114 13879 11117
rect 17953 11114 18019 11117
rect 13813 11112 18019 11114
rect 13813 11056 13818 11112
rect 13874 11056 17958 11112
rect 18014 11056 18019 11112
rect 13813 11054 18019 11056
rect 13813 11051 13879 11054
rect 17953 11051 18019 11054
rect 0 10978 800 11008
rect 3693 10978 3759 10981
rect 0 10976 3759 10978
rect 0 10920 3698 10976
rect 3754 10920 3759 10976
rect 0 10918 3759 10920
rect 0 10888 800 10918
rect 3693 10915 3759 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 19200 10842 20000 10872
rect 16254 10782 20000 10842
rect 5441 10706 5507 10709
rect 4662 10704 5507 10706
rect 4662 10648 5446 10704
rect 5502 10648 5507 10704
rect 4662 10646 5507 10648
rect 0 10570 800 10600
rect 4662 10570 4722 10646
rect 5441 10643 5507 10646
rect 0 10510 4722 10570
rect 4889 10570 4955 10573
rect 8201 10570 8267 10573
rect 16254 10570 16314 10782
rect 19200 10752 20000 10782
rect 4889 10568 16314 10570
rect 4889 10512 4894 10568
rect 4950 10512 8206 10568
rect 8262 10512 16314 10568
rect 4889 10510 16314 10512
rect 0 10480 800 10510
rect 4889 10507 4955 10510
rect 8201 10507 8267 10510
rect 3233 10434 3299 10437
rect 4889 10434 4955 10437
rect 6545 10434 6611 10437
rect 3233 10432 6611 10434
rect 3233 10376 3238 10432
rect 3294 10376 4894 10432
rect 4950 10376 6550 10432
rect 6606 10376 6611 10432
rect 3233 10374 6611 10376
rect 3233 10371 3299 10374
rect 4889 10371 4955 10374
rect 6545 10371 6611 10374
rect 11605 10434 11671 10437
rect 12065 10434 12131 10437
rect 11605 10432 12131 10434
rect 11605 10376 11610 10432
rect 11666 10376 12070 10432
rect 12126 10376 12131 10432
rect 11605 10374 12131 10376
rect 11605 10371 11671 10374
rect 12065 10371 12131 10374
rect 16941 10434 17007 10437
rect 19200 10434 20000 10464
rect 16941 10432 20000 10434
rect 16941 10376 16946 10432
rect 17002 10376 20000 10432
rect 16941 10374 20000 10376
rect 16941 10371 17007 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19200 10344 20000 10374
rect 12805 10303 13125 10304
rect 4337 10298 4403 10301
rect 6361 10298 6427 10301
rect 4337 10296 6427 10298
rect 4337 10240 4342 10296
rect 4398 10240 6366 10296
rect 6422 10240 6427 10296
rect 4337 10238 6427 10240
rect 4337 10235 4403 10238
rect 6361 10235 6427 10238
rect 11789 10298 11855 10301
rect 12433 10298 12499 10301
rect 11789 10296 12499 10298
rect 11789 10240 11794 10296
rect 11850 10240 12438 10296
rect 12494 10240 12499 10296
rect 11789 10238 12499 10240
rect 11789 10235 11855 10238
rect 12433 10235 12499 10238
rect 13537 10298 13603 10301
rect 14641 10298 14707 10301
rect 18137 10298 18203 10301
rect 13537 10296 18203 10298
rect 13537 10240 13542 10296
rect 13598 10240 14646 10296
rect 14702 10240 18142 10296
rect 18198 10240 18203 10296
rect 13537 10238 18203 10240
rect 13537 10235 13603 10238
rect 14641 10235 14707 10238
rect 18137 10235 18203 10238
rect 0 10162 800 10192
rect 3601 10162 3667 10165
rect 4153 10162 4219 10165
rect 0 10160 4219 10162
rect 0 10104 3606 10160
rect 3662 10104 4158 10160
rect 4214 10104 4219 10160
rect 0 10102 4219 10104
rect 6364 10162 6424 10235
rect 9397 10162 9463 10165
rect 6364 10160 9463 10162
rect 6364 10104 9402 10160
rect 9458 10104 9463 10160
rect 6364 10102 9463 10104
rect 0 10072 800 10102
rect 3601 10099 3667 10102
rect 4153 10099 4219 10102
rect 9397 10099 9463 10102
rect 10869 10162 10935 10165
rect 12157 10162 12223 10165
rect 18413 10162 18479 10165
rect 10869 10160 18479 10162
rect 10869 10104 10874 10160
rect 10930 10104 12162 10160
rect 12218 10104 18418 10160
rect 18474 10104 18479 10160
rect 10869 10102 18479 10104
rect 10869 10099 10935 10102
rect 12157 10099 12223 10102
rect 18413 10099 18479 10102
rect 6361 10026 6427 10029
rect 8017 10026 8083 10029
rect 6361 10024 8083 10026
rect 6361 9968 6366 10024
rect 6422 9968 8022 10024
rect 8078 9968 8083 10024
rect 6361 9966 8083 9968
rect 6361 9963 6427 9966
rect 8017 9963 8083 9966
rect 10685 10026 10751 10029
rect 17125 10026 17191 10029
rect 10685 10024 17191 10026
rect 10685 9968 10690 10024
rect 10746 9968 17130 10024
rect 17186 9968 17191 10024
rect 10685 9966 17191 9968
rect 10685 9963 10751 9966
rect 17125 9963 17191 9966
rect 18137 10026 18203 10029
rect 19200 10026 20000 10056
rect 18137 10024 20000 10026
rect 18137 9968 18142 10024
rect 18198 9968 20000 10024
rect 18137 9966 20000 9968
rect 18137 9963 18203 9966
rect 19200 9936 20000 9966
rect 13261 9890 13327 9893
rect 13905 9890 13971 9893
rect 13261 9888 13971 9890
rect 13261 9832 13266 9888
rect 13322 9832 13910 9888
rect 13966 9832 13971 9888
rect 13261 9830 13971 9832
rect 13261 9827 13327 9830
rect 13905 9827 13971 9830
rect 3909 9824 4229 9825
rect 0 9754 800 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 9759 16090 9760
rect 3509 9754 3575 9757
rect 0 9752 3575 9754
rect 0 9696 3514 9752
rect 3570 9696 3575 9752
rect 0 9694 3575 9696
rect 0 9664 800 9694
rect 3509 9691 3575 9694
rect 10317 9754 10383 9757
rect 13537 9754 13603 9757
rect 10317 9752 13603 9754
rect 10317 9696 10322 9752
rect 10378 9696 13542 9752
rect 13598 9696 13603 9752
rect 10317 9694 13603 9696
rect 10317 9691 10383 9694
rect 13537 9691 13603 9694
rect 2589 9618 2655 9621
rect 4521 9618 4587 9621
rect 2589 9616 4587 9618
rect 2589 9560 2594 9616
rect 2650 9560 4526 9616
rect 4582 9560 4587 9616
rect 2589 9558 4587 9560
rect 2589 9555 2655 9558
rect 4521 9555 4587 9558
rect 6821 9618 6887 9621
rect 8017 9618 8083 9621
rect 6821 9616 8083 9618
rect 6821 9560 6826 9616
rect 6882 9560 8022 9616
rect 8078 9560 8083 9616
rect 6821 9558 8083 9560
rect 6821 9555 6887 9558
rect 8017 9555 8083 9558
rect 11605 9618 11671 9621
rect 14181 9618 14247 9621
rect 11605 9616 14247 9618
rect 11605 9560 11610 9616
rect 11666 9560 14186 9616
rect 14242 9560 14247 9616
rect 11605 9558 14247 9560
rect 11605 9555 11671 9558
rect 14181 9555 14247 9558
rect 15009 9618 15075 9621
rect 17401 9618 17467 9621
rect 19200 9618 20000 9648
rect 15009 9616 20000 9618
rect 15009 9560 15014 9616
rect 15070 9560 17406 9616
rect 17462 9560 20000 9616
rect 15009 9558 20000 9560
rect 15009 9555 15075 9558
rect 17401 9555 17467 9558
rect 19200 9528 20000 9558
rect 4521 9482 4587 9485
rect 8569 9482 8635 9485
rect 4521 9480 8635 9482
rect 4521 9424 4526 9480
rect 4582 9424 8574 9480
rect 8630 9424 8635 9480
rect 4521 9422 8635 9424
rect 4521 9419 4587 9422
rect 8569 9419 8635 9422
rect 0 9346 800 9376
rect 4153 9346 4219 9349
rect 0 9344 4219 9346
rect 0 9288 4158 9344
rect 4214 9288 4219 9344
rect 0 9286 4219 9288
rect 0 9256 800 9286
rect 4153 9283 4219 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 7465 9210 7531 9213
rect 7649 9210 7715 9213
rect 12433 9212 12499 9213
rect 7465 9208 7715 9210
rect 7465 9152 7470 9208
rect 7526 9152 7654 9208
rect 7710 9152 7715 9208
rect 7465 9150 7715 9152
rect 7465 9147 7531 9150
rect 7649 9147 7715 9150
rect 12382 9148 12388 9212
rect 12452 9210 12499 9212
rect 17769 9210 17835 9213
rect 19200 9210 20000 9240
rect 12452 9208 12544 9210
rect 12494 9152 12544 9208
rect 12452 9150 12544 9152
rect 17769 9208 20000 9210
rect 17769 9152 17774 9208
rect 17830 9152 20000 9208
rect 17769 9150 20000 9152
rect 12452 9148 12499 9150
rect 12433 9147 12499 9148
rect 17769 9147 17835 9150
rect 19200 9120 20000 9150
rect 7005 9074 7071 9077
rect 7281 9074 7347 9077
rect 10409 9076 10475 9077
rect 7005 9072 7347 9074
rect 7005 9016 7010 9072
rect 7066 9016 7286 9072
rect 7342 9016 7347 9072
rect 7005 9014 7347 9016
rect 7005 9011 7071 9014
rect 7281 9011 7347 9014
rect 10358 9012 10364 9076
rect 10428 9074 10475 9076
rect 13169 9074 13235 9077
rect 10428 9072 13235 9074
rect 10470 9016 13174 9072
rect 13230 9016 13235 9072
rect 10428 9014 13235 9016
rect 10428 9012 10475 9014
rect 10409 9011 10475 9012
rect 13169 9011 13235 9014
rect 0 8938 800 8968
rect 2957 8938 3023 8941
rect 0 8936 3023 8938
rect 0 8880 2962 8936
rect 3018 8880 3023 8936
rect 0 8878 3023 8880
rect 0 8848 800 8878
rect 2957 8875 3023 8878
rect 3417 8938 3483 8941
rect 10593 8938 10659 8941
rect 12341 8938 12407 8941
rect 12525 8940 12591 8941
rect 12525 8938 12572 8940
rect 3417 8936 10472 8938
rect 3417 8880 3422 8936
rect 3478 8880 10472 8936
rect 3417 8878 10472 8880
rect 3417 8875 3483 8878
rect 6177 8802 6243 8805
rect 8477 8802 8543 8805
rect 6177 8800 8543 8802
rect 6177 8744 6182 8800
rect 6238 8744 8482 8800
rect 8538 8744 8543 8800
rect 6177 8742 8543 8744
rect 10412 8802 10472 8878
rect 10593 8936 12407 8938
rect 10593 8880 10598 8936
rect 10654 8880 12346 8936
rect 12402 8880 12407 8936
rect 10593 8878 12407 8880
rect 12480 8936 12572 8938
rect 12636 8938 12642 8940
rect 17125 8938 17191 8941
rect 12636 8936 17191 8938
rect 12480 8880 12530 8936
rect 12636 8880 17130 8936
rect 17186 8880 17191 8936
rect 12480 8878 12572 8880
rect 10593 8875 10659 8878
rect 12341 8875 12407 8878
rect 12525 8876 12572 8878
rect 12636 8878 17191 8880
rect 12636 8876 12642 8878
rect 12525 8875 12591 8876
rect 17125 8875 17191 8878
rect 12433 8802 12499 8805
rect 10412 8800 12499 8802
rect 10412 8744 12438 8800
rect 12494 8744 12499 8800
rect 10412 8742 12499 8744
rect 6177 8739 6243 8742
rect 8477 8739 8543 8742
rect 12433 8739 12499 8742
rect 14733 8802 14799 8805
rect 15510 8802 15516 8804
rect 14733 8800 15516 8802
rect 14733 8744 14738 8800
rect 14794 8744 15516 8800
rect 14733 8742 15516 8744
rect 14733 8739 14799 8742
rect 15510 8740 15516 8742
rect 15580 8740 15586 8804
rect 16573 8802 16639 8805
rect 19200 8802 20000 8832
rect 16573 8800 20000 8802
rect 16573 8744 16578 8800
rect 16634 8744 20000 8800
rect 16573 8742 20000 8744
rect 16573 8739 16639 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 19200 8712 20000 8742
rect 15770 8671 16090 8672
rect 7373 8666 7439 8669
rect 7598 8666 7604 8668
rect 7373 8664 7604 8666
rect 7373 8608 7378 8664
rect 7434 8608 7604 8664
rect 7373 8606 7604 8608
rect 7373 8603 7439 8606
rect 7598 8604 7604 8606
rect 7668 8604 7674 8668
rect 0 8530 800 8560
rect 3417 8530 3483 8533
rect 0 8528 3483 8530
rect 0 8472 3422 8528
rect 3478 8472 3483 8528
rect 0 8470 3483 8472
rect 0 8440 800 8470
rect 3417 8467 3483 8470
rect 6269 8530 6335 8533
rect 8753 8530 8819 8533
rect 6269 8528 8819 8530
rect 6269 8472 6274 8528
rect 6330 8472 8758 8528
rect 8814 8472 8819 8528
rect 6269 8470 8819 8472
rect 6269 8467 6335 8470
rect 8753 8467 8819 8470
rect 10133 8530 10199 8533
rect 13629 8530 13695 8533
rect 10133 8528 13695 8530
rect 10133 8472 10138 8528
rect 10194 8472 13634 8528
rect 13690 8472 13695 8528
rect 10133 8470 13695 8472
rect 10133 8467 10199 8470
rect 13629 8467 13695 8470
rect 3969 8394 4035 8397
rect 7005 8394 7071 8397
rect 3969 8392 7071 8394
rect 3969 8336 3974 8392
rect 4030 8336 7010 8392
rect 7066 8336 7071 8392
rect 3969 8334 7071 8336
rect 3969 8331 4035 8334
rect 7005 8331 7071 8334
rect 10869 8394 10935 8397
rect 11053 8394 11119 8397
rect 10869 8392 11119 8394
rect 10869 8336 10874 8392
rect 10930 8336 11058 8392
rect 11114 8336 11119 8392
rect 10869 8334 11119 8336
rect 10869 8331 10935 8334
rect 11053 8331 11119 8334
rect 17861 8258 17927 8261
rect 19200 8258 20000 8288
rect 17861 8256 20000 8258
rect 17861 8200 17866 8256
rect 17922 8200 20000 8256
rect 17861 8198 20000 8200
rect 17861 8195 17927 8198
rect 6874 8192 7194 8193
rect 0 8122 800 8152
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 19200 8168 20000 8198
rect 12805 8127 13125 8128
rect 3785 8122 3851 8125
rect 0 8120 3851 8122
rect 0 8064 3790 8120
rect 3846 8064 3851 8120
rect 0 8062 3851 8064
rect 0 8032 800 8062
rect 3785 8059 3851 8062
rect 5993 7986 6059 7989
rect 8753 7986 8819 7989
rect 5993 7984 8819 7986
rect 5993 7928 5998 7984
rect 6054 7928 8758 7984
rect 8814 7928 8819 7984
rect 5993 7926 8819 7928
rect 5993 7923 6059 7926
rect 8753 7923 8819 7926
rect 9305 7986 9371 7989
rect 10409 7986 10475 7989
rect 9305 7984 10475 7986
rect 9305 7928 9310 7984
rect 9366 7928 10414 7984
rect 10470 7928 10475 7984
rect 9305 7926 10475 7928
rect 9305 7923 9371 7926
rect 10409 7923 10475 7926
rect 2497 7850 2563 7853
rect 7465 7850 7531 7853
rect 2497 7848 7531 7850
rect 2497 7792 2502 7848
rect 2558 7792 7470 7848
rect 7526 7792 7531 7848
rect 2497 7790 7531 7792
rect 2497 7787 2563 7790
rect 7465 7787 7531 7790
rect 10041 7850 10107 7853
rect 11462 7850 11468 7852
rect 10041 7848 11468 7850
rect 10041 7792 10046 7848
rect 10102 7792 11468 7848
rect 10041 7790 11468 7792
rect 10041 7787 10107 7790
rect 11462 7788 11468 7790
rect 11532 7850 11538 7852
rect 13261 7850 13327 7853
rect 11532 7848 13327 7850
rect 11532 7792 13266 7848
rect 13322 7792 13327 7848
rect 11532 7790 13327 7792
rect 11532 7788 11538 7790
rect 13261 7787 13327 7790
rect 18045 7850 18111 7853
rect 19200 7850 20000 7880
rect 18045 7848 20000 7850
rect 18045 7792 18050 7848
rect 18106 7792 20000 7848
rect 18045 7790 20000 7792
rect 18045 7787 18111 7790
rect 19200 7760 20000 7790
rect 0 7714 800 7744
rect 1853 7714 1919 7717
rect 0 7712 1919 7714
rect 0 7656 1858 7712
rect 1914 7656 1919 7712
rect 0 7654 1919 7656
rect 0 7624 800 7654
rect 1853 7651 1919 7654
rect 10961 7714 11027 7717
rect 14917 7714 14983 7717
rect 10961 7712 14983 7714
rect 10961 7656 10966 7712
rect 11022 7656 14922 7712
rect 14978 7656 14983 7712
rect 10961 7654 14983 7656
rect 10961 7651 11027 7654
rect 14917 7651 14983 7654
rect 3909 7648 4229 7649
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 10225 7578 10291 7581
rect 10358 7578 10364 7580
rect 10225 7576 10364 7578
rect 10225 7520 10230 7576
rect 10286 7520 10364 7576
rect 10225 7518 10364 7520
rect 10225 7515 10291 7518
rect 10358 7516 10364 7518
rect 10428 7516 10434 7580
rect 10501 7578 10567 7581
rect 15469 7578 15535 7581
rect 10501 7576 15535 7578
rect 10501 7520 10506 7576
rect 10562 7520 15474 7576
rect 15530 7520 15535 7576
rect 10501 7518 15535 7520
rect 10501 7515 10567 7518
rect 15469 7515 15535 7518
rect 11329 7442 11395 7445
rect 12065 7442 12131 7445
rect 16297 7442 16363 7445
rect 11329 7440 12131 7442
rect 11329 7384 11334 7440
rect 11390 7384 12070 7440
rect 12126 7384 12131 7440
rect 12390 7440 16363 7442
rect 12390 7408 16302 7440
rect 11329 7382 12131 7384
rect 11329 7379 11395 7382
rect 12065 7379 12131 7382
rect 12344 7384 16302 7408
rect 16358 7384 16363 7440
rect 12344 7382 16363 7384
rect 12344 7348 12450 7382
rect 16297 7379 16363 7382
rect 18229 7442 18295 7445
rect 19200 7442 20000 7472
rect 18229 7440 20000 7442
rect 18229 7384 18234 7440
rect 18290 7384 20000 7440
rect 18229 7382 20000 7384
rect 18229 7379 18295 7382
rect 19200 7352 20000 7382
rect 0 7306 800 7336
rect 4061 7306 4127 7309
rect 0 7304 4127 7306
rect 0 7248 4066 7304
rect 4122 7248 4127 7304
rect 0 7246 4127 7248
rect 0 7216 800 7246
rect 4061 7243 4127 7246
rect 9121 7306 9187 7309
rect 12344 7306 12404 7348
rect 9121 7304 12404 7306
rect 9121 7248 9126 7304
rect 9182 7248 12404 7304
rect 9121 7246 12404 7248
rect 9121 7243 9187 7246
rect 3693 7170 3759 7173
rect 6361 7170 6427 7173
rect 3693 7168 6427 7170
rect 3693 7112 3698 7168
rect 3754 7112 6366 7168
rect 6422 7112 6427 7168
rect 3693 7110 6427 7112
rect 3693 7107 3759 7110
rect 6361 7107 6427 7110
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 1577 7034 1643 7037
rect 4429 7034 4495 7037
rect 1577 7032 4495 7034
rect 1577 6976 1582 7032
rect 1638 6976 4434 7032
rect 4490 6976 4495 7032
rect 1577 6974 4495 6976
rect 1577 6971 1643 6974
rect 4429 6971 4495 6974
rect 18413 7034 18479 7037
rect 19200 7034 20000 7064
rect 18413 7032 20000 7034
rect 18413 6976 18418 7032
rect 18474 6976 20000 7032
rect 18413 6974 20000 6976
rect 18413 6971 18479 6974
rect 19200 6944 20000 6974
rect 0 6898 800 6928
rect 1761 6898 1827 6901
rect 0 6896 1827 6898
rect 0 6840 1766 6896
rect 1822 6840 1827 6896
rect 0 6838 1827 6840
rect 0 6808 800 6838
rect 1761 6835 1827 6838
rect 1945 6898 2011 6901
rect 9121 6898 9187 6901
rect 1945 6896 9187 6898
rect 1945 6840 1950 6896
rect 2006 6840 9126 6896
rect 9182 6840 9187 6896
rect 1945 6838 9187 6840
rect 1945 6835 2011 6838
rect 9121 6835 9187 6838
rect 11237 6898 11303 6901
rect 14549 6898 14615 6901
rect 11237 6896 14615 6898
rect 11237 6840 11242 6896
rect 11298 6840 14554 6896
rect 14610 6840 14615 6896
rect 11237 6838 14615 6840
rect 11237 6835 11303 6838
rect 14549 6835 14615 6838
rect 6361 6764 6427 6765
rect 6310 6700 6316 6764
rect 6380 6762 6427 6764
rect 6380 6760 6472 6762
rect 6422 6704 6472 6760
rect 6380 6702 6472 6704
rect 6380 6700 6427 6702
rect 6361 6699 6427 6700
rect 18045 6626 18111 6629
rect 19200 6626 20000 6656
rect 18045 6624 20000 6626
rect 18045 6568 18050 6624
rect 18106 6568 20000 6624
rect 18045 6566 20000 6568
rect 18045 6563 18111 6566
rect 3909 6560 4229 6561
rect 0 6490 800 6520
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 19200 6536 20000 6566
rect 15770 6495 16090 6496
rect 2773 6490 2839 6493
rect 0 6488 2839 6490
rect 0 6432 2778 6488
rect 2834 6432 2839 6488
rect 0 6430 2839 6432
rect 0 6400 800 6430
rect 2773 6427 2839 6430
rect 6821 6354 6887 6357
rect 7649 6354 7715 6357
rect 6821 6352 7715 6354
rect 6821 6296 6826 6352
rect 6882 6296 7654 6352
rect 7710 6296 7715 6352
rect 6821 6294 7715 6296
rect 6821 6291 6887 6294
rect 7649 6291 7715 6294
rect 10593 6354 10659 6357
rect 11237 6354 11303 6357
rect 10593 6352 11303 6354
rect 10593 6296 10598 6352
rect 10654 6296 11242 6352
rect 11298 6296 11303 6352
rect 10593 6294 11303 6296
rect 10593 6291 10659 6294
rect 11237 6291 11303 6294
rect 10593 6218 10659 6221
rect 12525 6218 12591 6221
rect 10593 6216 12591 6218
rect 10593 6160 10598 6216
rect 10654 6160 12530 6216
rect 12586 6160 12591 6216
rect 10593 6158 12591 6160
rect 10593 6155 10659 6158
rect 12525 6155 12591 6158
rect 18229 6218 18295 6221
rect 19200 6218 20000 6248
rect 18229 6216 20000 6218
rect 18229 6160 18234 6216
rect 18290 6160 20000 6216
rect 18229 6158 20000 6160
rect 18229 6155 18295 6158
rect 19200 6128 20000 6158
rect 0 6082 800 6112
rect 3233 6082 3299 6085
rect 0 6080 3299 6082
rect 0 6024 3238 6080
rect 3294 6024 3299 6080
rect 0 6022 3299 6024
rect 0 5992 800 6022
rect 3233 6019 3299 6022
rect 6874 6016 7194 6017
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 5951 13125 5952
rect 11237 5810 11303 5813
rect 13721 5810 13787 5813
rect 11237 5808 13787 5810
rect 11237 5752 11242 5808
rect 11298 5752 13726 5808
rect 13782 5752 13787 5808
rect 11237 5750 13787 5752
rect 11237 5747 11303 5750
rect 13721 5747 13787 5750
rect 10317 5674 10383 5677
rect 12382 5674 12388 5676
rect 10317 5672 12388 5674
rect 10317 5616 10322 5672
rect 10378 5616 12388 5672
rect 10317 5614 12388 5616
rect 10317 5611 10383 5614
rect 12382 5612 12388 5614
rect 12452 5674 12458 5676
rect 14549 5674 14615 5677
rect 12452 5672 14615 5674
rect 12452 5616 14554 5672
rect 14610 5616 14615 5672
rect 12452 5614 14615 5616
rect 12452 5612 12458 5614
rect 14549 5611 14615 5614
rect 18413 5674 18479 5677
rect 19200 5674 20000 5704
rect 18413 5672 20000 5674
rect 18413 5616 18418 5672
rect 18474 5616 20000 5672
rect 18413 5614 20000 5616
rect 18413 5611 18479 5614
rect 19200 5584 20000 5614
rect 0 5538 800 5568
rect 3693 5538 3759 5541
rect 0 5536 3759 5538
rect 0 5480 3698 5536
rect 3754 5480 3759 5536
rect 0 5478 3759 5480
rect 0 5448 800 5478
rect 3693 5475 3759 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 11973 5402 12039 5405
rect 13537 5402 13603 5405
rect 11973 5400 13603 5402
rect 11973 5344 11978 5400
rect 12034 5344 13542 5400
rect 13598 5344 13603 5400
rect 11973 5342 13603 5344
rect 11973 5339 12039 5342
rect 13537 5339 13603 5342
rect 5165 5266 5231 5269
rect 8661 5266 8727 5269
rect 5165 5264 8727 5266
rect 5165 5208 5170 5264
rect 5226 5208 8666 5264
rect 8722 5208 8727 5264
rect 5165 5206 8727 5208
rect 5165 5203 5231 5206
rect 8661 5203 8727 5206
rect 10593 5266 10659 5269
rect 15929 5266 15995 5269
rect 10593 5264 15995 5266
rect 10593 5208 10598 5264
rect 10654 5208 15934 5264
rect 15990 5208 15995 5264
rect 10593 5206 15995 5208
rect 10593 5203 10659 5206
rect 15929 5203 15995 5206
rect 17861 5266 17927 5269
rect 19200 5266 20000 5296
rect 17861 5264 20000 5266
rect 17861 5208 17866 5264
rect 17922 5208 20000 5264
rect 17861 5206 20000 5208
rect 17861 5203 17927 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 3141 5130 3207 5133
rect 0 5128 3207 5130
rect 0 5072 3146 5128
rect 3202 5072 3207 5128
rect 0 5070 3207 5072
rect 0 5040 800 5070
rect 3141 5067 3207 5070
rect 6913 5130 6979 5133
rect 7649 5130 7715 5133
rect 6913 5128 7715 5130
rect 6913 5072 6918 5128
rect 6974 5072 7654 5128
rect 7710 5072 7715 5128
rect 6913 5070 7715 5072
rect 6913 5067 6979 5070
rect 7649 5067 7715 5070
rect 2037 4994 2103 4997
rect 4429 4994 4495 4997
rect 6637 4994 6703 4997
rect 2037 4992 6703 4994
rect 2037 4936 2042 4992
rect 2098 4936 4434 4992
rect 4490 4936 6642 4992
rect 6698 4936 6703 4992
rect 2037 4934 6703 4936
rect 2037 4931 2103 4934
rect 4429 4931 4495 4934
rect 6637 4931 6703 4934
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 10409 4858 10475 4861
rect 12617 4858 12683 4861
rect 10409 4856 12683 4858
rect 10409 4800 10414 4856
rect 10470 4800 12622 4856
rect 12678 4800 12683 4856
rect 10409 4798 12683 4800
rect 10409 4795 10475 4798
rect 12617 4795 12683 4798
rect 18321 4858 18387 4861
rect 19200 4858 20000 4888
rect 18321 4856 20000 4858
rect 18321 4800 18326 4856
rect 18382 4800 20000 4856
rect 18321 4798 20000 4800
rect 18321 4795 18387 4798
rect 19200 4768 20000 4798
rect 0 4722 800 4752
rect 2773 4722 2839 4725
rect 0 4720 2839 4722
rect 0 4664 2778 4720
rect 2834 4664 2839 4720
rect 0 4662 2839 4664
rect 0 4632 800 4662
rect 2773 4659 2839 4662
rect 4521 4722 4587 4725
rect 6913 4722 6979 4725
rect 4521 4720 6979 4722
rect 4521 4664 4526 4720
rect 4582 4664 6918 4720
rect 6974 4664 6979 4720
rect 4521 4662 6979 4664
rect 4521 4659 4587 4662
rect 6913 4659 6979 4662
rect 7557 4722 7623 4725
rect 12617 4722 12683 4725
rect 7557 4720 12683 4722
rect 7557 4664 7562 4720
rect 7618 4664 12622 4720
rect 12678 4664 12683 4720
rect 7557 4662 12683 4664
rect 7557 4659 7623 4662
rect 12617 4659 12683 4662
rect 8477 4586 8543 4589
rect 9397 4586 9463 4589
rect 8477 4584 9463 4586
rect 8477 4528 8482 4584
rect 8538 4528 9402 4584
rect 9458 4528 9463 4584
rect 8477 4526 9463 4528
rect 8477 4523 8543 4526
rect 9397 4523 9463 4526
rect 12249 4586 12315 4589
rect 12801 4586 12867 4589
rect 12249 4584 12867 4586
rect 12249 4528 12254 4584
rect 12310 4528 12806 4584
rect 12862 4528 12867 4584
rect 12249 4526 12867 4528
rect 12249 4523 12315 4526
rect 12801 4523 12867 4526
rect 4337 4450 4403 4453
rect 5441 4450 5507 4453
rect 8845 4450 8911 4453
rect 12617 4452 12683 4453
rect 12566 4450 12572 4452
rect 4337 4448 8911 4450
rect 4337 4392 4342 4448
rect 4398 4392 5446 4448
rect 5502 4392 8850 4448
rect 8906 4392 8911 4448
rect 4337 4390 8911 4392
rect 12526 4390 12572 4450
rect 12636 4448 12683 4452
rect 12678 4392 12683 4448
rect 4337 4387 4403 4390
rect 5441 4387 5507 4390
rect 8845 4387 8911 4390
rect 12566 4388 12572 4390
rect 12636 4388 12683 4392
rect 12617 4387 12683 4388
rect 18045 4450 18111 4453
rect 19200 4450 20000 4480
rect 18045 4448 20000 4450
rect 18045 4392 18050 4448
rect 18106 4392 20000 4448
rect 18045 4390 20000 4392
rect 18045 4387 18111 4390
rect 3909 4384 4229 4385
rect 0 4314 800 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19200 4360 20000 4390
rect 15770 4319 16090 4320
rect 2957 4314 3023 4317
rect 0 4312 3023 4314
rect 0 4256 2962 4312
rect 3018 4256 3023 4312
rect 0 4254 3023 4256
rect 0 4224 800 4254
rect 2957 4251 3023 4254
rect 10225 4314 10291 4317
rect 13905 4314 13971 4317
rect 10225 4312 13971 4314
rect 10225 4256 10230 4312
rect 10286 4256 13910 4312
rect 13966 4256 13971 4312
rect 10225 4254 13971 4256
rect 10225 4251 10291 4254
rect 13905 4251 13971 4254
rect 1761 4178 1827 4181
rect 5809 4178 5875 4181
rect 7741 4178 7807 4181
rect 9581 4178 9647 4181
rect 1761 4176 5875 4178
rect 1761 4120 1766 4176
rect 1822 4120 5814 4176
rect 5870 4120 5875 4176
rect 1761 4118 5875 4120
rect 1761 4115 1827 4118
rect 5809 4115 5875 4118
rect 5950 4176 9647 4178
rect 5950 4120 7746 4176
rect 7802 4120 9586 4176
rect 9642 4120 9647 4176
rect 5950 4118 9647 4120
rect 2129 4042 2195 4045
rect 3877 4042 3943 4045
rect 2129 4040 3943 4042
rect 2129 3984 2134 4040
rect 2190 3984 3882 4040
rect 3938 3984 3943 4040
rect 2129 3982 3943 3984
rect 2129 3979 2195 3982
rect 3877 3979 3943 3982
rect 0 3906 800 3936
rect 1393 3906 1459 3909
rect 0 3904 1459 3906
rect 0 3848 1398 3904
rect 1454 3848 1459 3904
rect 0 3846 1459 3848
rect 0 3816 800 3846
rect 1393 3843 1459 3846
rect 1577 3906 1643 3909
rect 2313 3906 2379 3909
rect 5950 3906 6010 4118
rect 7741 4115 7807 4118
rect 9581 4115 9647 4118
rect 10869 4178 10935 4181
rect 11605 4178 11671 4181
rect 10869 4176 11671 4178
rect 10869 4120 10874 4176
rect 10930 4120 11610 4176
rect 11666 4120 11671 4176
rect 10869 4118 11671 4120
rect 10869 4115 10935 4118
rect 11605 4115 11671 4118
rect 13077 4178 13143 4181
rect 14457 4178 14523 4181
rect 13077 4176 14523 4178
rect 13077 4120 13082 4176
rect 13138 4120 14462 4176
rect 14518 4120 14523 4176
rect 13077 4118 14523 4120
rect 13077 4115 13143 4118
rect 14457 4115 14523 4118
rect 6637 4042 6703 4045
rect 8477 4042 8543 4045
rect 6637 4040 8543 4042
rect 6637 3984 6642 4040
rect 6698 3984 8482 4040
rect 8538 3984 8543 4040
rect 6637 3982 8543 3984
rect 6637 3979 6703 3982
rect 8477 3979 8543 3982
rect 13905 4042 13971 4045
rect 14641 4042 14707 4045
rect 13905 4040 14707 4042
rect 13905 3984 13910 4040
rect 13966 3984 14646 4040
rect 14702 3984 14707 4040
rect 13905 3982 14707 3984
rect 13905 3979 13971 3982
rect 14641 3979 14707 3982
rect 18229 4042 18295 4045
rect 19200 4042 20000 4072
rect 18229 4040 20000 4042
rect 18229 3984 18234 4040
rect 18290 3984 20000 4040
rect 18229 3982 20000 3984
rect 18229 3979 18295 3982
rect 19200 3952 20000 3982
rect 1577 3904 6010 3906
rect 1577 3848 1582 3904
rect 1638 3848 2318 3904
rect 2374 3848 6010 3904
rect 1577 3846 6010 3848
rect 1577 3843 1643 3846
rect 2313 3843 2379 3846
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 9765 3770 9831 3773
rect 10409 3770 10475 3773
rect 9765 3768 10475 3770
rect 9765 3712 9770 3768
rect 9826 3712 10414 3768
rect 10470 3712 10475 3768
rect 9765 3710 10475 3712
rect 9765 3707 9831 3710
rect 10409 3707 10475 3710
rect 5993 3634 6059 3637
rect 12893 3634 12959 3637
rect 16941 3634 17007 3637
rect 5993 3632 12818 3634
rect 5993 3576 5998 3632
rect 6054 3576 12818 3632
rect 5993 3574 12818 3576
rect 5993 3571 6059 3574
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 3877 3498 3943 3501
rect 4337 3498 4403 3501
rect 6310 3498 6316 3500
rect 3877 3496 6316 3498
rect 3877 3440 3882 3496
rect 3938 3440 4342 3496
rect 4398 3440 6316 3496
rect 3877 3438 6316 3440
rect 3877 3435 3943 3438
rect 4337 3435 4403 3438
rect 6310 3436 6316 3438
rect 6380 3498 6386 3500
rect 9765 3498 9831 3501
rect 6380 3496 9831 3498
rect 6380 3440 9770 3496
rect 9826 3440 9831 3496
rect 6380 3438 9831 3440
rect 12758 3498 12818 3574
rect 12893 3632 17007 3634
rect 12893 3576 12898 3632
rect 12954 3576 16946 3632
rect 17002 3576 17007 3632
rect 12893 3574 17007 3576
rect 12893 3571 12959 3574
rect 16941 3571 17007 3574
rect 17677 3634 17743 3637
rect 19200 3634 20000 3664
rect 17677 3632 20000 3634
rect 17677 3576 17682 3632
rect 17738 3576 20000 3632
rect 17677 3574 20000 3576
rect 17677 3571 17743 3574
rect 19200 3544 20000 3574
rect 17125 3498 17191 3501
rect 12758 3496 17191 3498
rect 12758 3440 17130 3496
rect 17186 3440 17191 3496
rect 12758 3438 17191 3440
rect 6380 3436 6386 3438
rect 9765 3435 9831 3438
rect 17125 3435 17191 3438
rect 10501 3362 10567 3365
rect 15377 3362 15443 3365
rect 10501 3360 15443 3362
rect 10501 3304 10506 3360
rect 10562 3304 15382 3360
rect 15438 3304 15443 3360
rect 10501 3302 15443 3304
rect 10501 3299 10567 3302
rect 15377 3299 15443 3302
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 18413 3226 18479 3229
rect 19200 3226 20000 3256
rect 18413 3224 20000 3226
rect 18413 3168 18418 3224
rect 18474 3168 20000 3224
rect 18413 3166 20000 3168
rect 18413 3163 18479 3166
rect 19200 3136 20000 3166
rect 0 3090 800 3120
rect 2865 3090 2931 3093
rect 0 3088 2931 3090
rect 0 3032 2870 3088
rect 2926 3032 2931 3088
rect 0 3030 2931 3032
rect 0 3000 800 3030
rect 2865 3027 2931 3030
rect 11237 2818 11303 2821
rect 11881 2818 11947 2821
rect 11237 2816 11947 2818
rect 11237 2760 11242 2816
rect 11298 2760 11886 2816
rect 11942 2760 11947 2816
rect 11237 2758 11947 2760
rect 11237 2755 11303 2758
rect 11881 2755 11947 2758
rect 6874 2752 7194 2753
rect 0 2682 800 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 2221 2682 2287 2685
rect 11421 2684 11487 2685
rect 11421 2682 11468 2684
rect 0 2680 2287 2682
rect 0 2624 2226 2680
rect 2282 2624 2287 2680
rect 0 2622 2287 2624
rect 11376 2680 11468 2682
rect 11376 2624 11426 2680
rect 11376 2622 11468 2624
rect 0 2592 800 2622
rect 2221 2619 2287 2622
rect 11421 2620 11468 2622
rect 11532 2620 11538 2684
rect 17861 2682 17927 2685
rect 19200 2682 20000 2712
rect 17861 2680 20000 2682
rect 17861 2624 17866 2680
rect 17922 2624 20000 2680
rect 17861 2622 20000 2624
rect 11421 2619 11487 2620
rect 17861 2619 17927 2622
rect 19200 2592 20000 2622
rect 1577 2546 1643 2549
rect 6913 2546 6979 2549
rect 9121 2546 9187 2549
rect 1577 2544 9187 2546
rect 1577 2488 1582 2544
rect 1638 2488 6918 2544
rect 6974 2488 9126 2544
rect 9182 2488 9187 2544
rect 1577 2486 9187 2488
rect 1577 2483 1643 2486
rect 6913 2483 6979 2486
rect 9121 2483 9187 2486
rect 0 2274 800 2304
rect 1853 2274 1919 2277
rect 0 2272 1919 2274
rect 0 2216 1858 2272
rect 1914 2216 1919 2272
rect 0 2214 1919 2216
rect 0 2184 800 2214
rect 1853 2211 1919 2214
rect 17769 2274 17835 2277
rect 19200 2274 20000 2304
rect 17769 2272 20000 2274
rect 17769 2216 17774 2272
rect 17830 2216 20000 2272
rect 17769 2214 20000 2216
rect 17769 2211 17835 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19200 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 800 1896
rect 2773 1866 2839 1869
rect 0 1864 2839 1866
rect 0 1808 2778 1864
rect 2834 1808 2839 1864
rect 0 1806 2839 1808
rect 0 1776 800 1806
rect 2773 1803 2839 1806
rect 17309 1866 17375 1869
rect 19200 1866 20000 1896
rect 17309 1864 20000 1866
rect 17309 1808 17314 1864
rect 17370 1808 20000 1864
rect 17309 1806 20000 1808
rect 17309 1803 17375 1806
rect 19200 1776 20000 1806
rect 0 1458 800 1488
rect 3141 1458 3207 1461
rect 0 1456 3207 1458
rect 0 1400 3146 1456
rect 3202 1400 3207 1456
rect 0 1398 3207 1400
rect 0 1368 800 1398
rect 3141 1395 3207 1398
rect 17033 1458 17099 1461
rect 19200 1458 20000 1488
rect 17033 1456 20000 1458
rect 17033 1400 17038 1456
rect 17094 1400 20000 1456
rect 17033 1398 20000 1400
rect 17033 1395 17099 1398
rect 19200 1368 20000 1398
rect 0 1050 800 1080
rect 3785 1050 3851 1053
rect 0 1048 3851 1050
rect 0 992 3790 1048
rect 3846 992 3851 1048
rect 0 990 3851 992
rect 0 960 800 990
rect 3785 987 3851 990
rect 17677 1050 17743 1053
rect 19200 1050 20000 1080
rect 17677 1048 20000 1050
rect 17677 992 17682 1048
rect 17738 992 20000 1048
rect 17677 990 20000 992
rect 17677 987 17743 990
rect 19200 960 20000 990
rect 0 642 800 672
rect 3417 642 3483 645
rect 0 640 3483 642
rect 0 584 3422 640
rect 3478 584 3483 640
rect 0 582 3483 584
rect 0 552 800 582
rect 3417 579 3483 582
rect 18229 642 18295 645
rect 19200 642 20000 672
rect 18229 640 20000 642
rect 18229 584 18234 640
rect 18290 584 20000 640
rect 18229 582 20000 584
rect 18229 579 18295 582
rect 19200 552 20000 582
rect 0 234 800 264
rect 1393 234 1459 237
rect 0 232 1459 234
rect 0 176 1398 232
rect 1454 176 1459 232
rect 0 174 1459 176
rect 0 144 800 174
rect 1393 171 1459 174
rect 17861 234 17927 237
rect 19200 234 20000 264
rect 17861 232 20000 234
rect 17861 176 17866 232
rect 17922 176 20000 232
rect 17861 174 20000 176
rect 17861 171 17927 174
rect 19200 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 15516 12276 15580 12340
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 7604 11112 7668 11116
rect 7604 11056 7618 11112
rect 7618 11056 7668 11112
rect 7604 11052 7668 11056
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 12388 9208 12452 9212
rect 12388 9152 12438 9208
rect 12438 9152 12452 9208
rect 12388 9148 12452 9152
rect 10364 9072 10428 9076
rect 10364 9016 10414 9072
rect 10414 9016 10428 9072
rect 10364 9012 10428 9016
rect 12572 8936 12636 8940
rect 12572 8880 12586 8936
rect 12586 8880 12636 8936
rect 12572 8876 12636 8880
rect 15516 8740 15580 8804
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 7604 8604 7668 8668
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 11468 7788 11532 7852
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 10364 7516 10428 7580
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 6316 6760 6380 6764
rect 6316 6704 6366 6760
rect 6366 6704 6380 6760
rect 6316 6700 6380 6704
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 12388 5612 12452 5676
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 12572 4448 12636 4452
rect 12572 4392 12622 4448
rect 12622 4392 12636 4448
rect 12572 4388 12636 4392
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 6316 3436 6380 3500
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 11468 2680 11532 2684
rect 11468 2624 11482 2680
rect 11482 2624 11532 2680
rect 11468 2620 11532 2624
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 7603 11116 7669 11117
rect 7603 11052 7604 11116
rect 7668 11052 7669 11116
rect 7603 11051 7669 11052
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 7606 8669 7666 11051
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 15770 14176 16091 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16091 14176
rect 15770 13088 16091 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16091 13088
rect 15515 12340 15581 12341
rect 15515 12276 15516 12340
rect 15580 12276 15581 12340
rect 15515 12275 15581 12276
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12387 9212 12453 9213
rect 12387 9148 12388 9212
rect 12452 9148 12453 9212
rect 12387 9147 12453 9148
rect 10363 9076 10429 9077
rect 10363 9012 10364 9076
rect 10428 9012 10429 9076
rect 10363 9011 10429 9012
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 7603 8668 7669 8669
rect 7603 8604 7604 8668
rect 7668 8604 7669 8668
rect 7603 8603 7669 8604
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6315 6764 6381 6765
rect 6315 6700 6316 6764
rect 6380 6700 6381 6764
rect 6315 6699 6381 6700
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 6318 3501 6378 6699
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6315 3500 6381 3501
rect 6315 3436 6316 3500
rect 6380 3436 6381 3500
rect 6315 3435 6381 3436
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 10366 7581 10426 9011
rect 11467 7852 11533 7853
rect 11467 7788 11468 7852
rect 11532 7788 11533 7852
rect 11467 7787 11533 7788
rect 10363 7580 10429 7581
rect 10363 7516 10364 7580
rect 10428 7516 10429 7580
rect 10363 7515 10429 7516
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 11470 2685 11530 7787
rect 12390 5677 12450 9147
rect 12571 8940 12637 8941
rect 12571 8876 12572 8940
rect 12636 8876 12637 8940
rect 12571 8875 12637 8876
rect 12387 5676 12453 5677
rect 12387 5612 12388 5676
rect 12452 5612 12453 5676
rect 12387 5611 12453 5612
rect 12574 4453 12634 8875
rect 12805 8192 13125 9216
rect 15518 8805 15578 12275
rect 15770 12000 16091 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16091 12000
rect 15770 10912 16091 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16091 10912
rect 15770 9824 16091 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16091 9824
rect 15515 8804 15581 8805
rect 15515 8740 15516 8804
rect 15580 8740 15581 8804
rect 15515 8739 15581 8740
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12571 4452 12637 4453
rect 12571 4388 12572 4452
rect 12636 4388 12637 4452
rect 12571 4387 12637 4388
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 11467 2684 11533 2685
rect 11467 2620 11468 2684
rect 11532 2620 11533 2684
rect 11467 2619 11533 2620
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 2128 13125 2688
rect 15770 8736 16091 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16091 8736
rect 15770 7648 16091 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16091 7648
rect 15770 6560 16091 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16091 6560
rect 15770 5472 16091 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16091 5472
rect 15770 4384 16091 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16091 4384
rect 15770 3296 16091 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16091 3296
rect 15770 2208 16091 3232
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16091 2208
rect 15770 2128 16091 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1564 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1564 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2116 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _40_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608910539
transform 1 0 2668 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3864 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3036 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608910539
transform 1 0 3220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4600 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4692 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1608910539
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_43
timestamp 1608910539
transform 1 0 5060 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1608910539
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 6072 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 5520 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5152 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8464 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8556 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_104
timestamp 1608910539
transform 1 0 10672 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1608910539
transform 1 0 9016 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9936 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_114
timestamp 1608910539
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1608910539
transform 1 0 11592 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1608910539
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1608910539
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1608910539
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11684 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13156 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_135 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 13524 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_141
timestamp 1608910539
transform 1 0 14076 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1608910539
transform 1 0 14076 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14168 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14352 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15824 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_148 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14720 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_162
timestamp 1608910539
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1608910539
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608910539
transform 1 0 16100 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_168
timestamp 1608910539
transform 1 0 16560 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_167
timestamp 1608910539
transform 1 0 16468 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1608910539
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1608910539
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608910539
transform 1 0 16836 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1608910539
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608910539
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1608910539
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608910539
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608910539
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608910539
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1608910539
transform 1 0 18492 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1608910539
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1608910539
transform 1 0 1472 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1608910539
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608910539
transform 1 0 2392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608910539
transform 1 0 2024 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608910539
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1608910539
transform 1 0 4876 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 6716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5704 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_65
timestamp 1608910539
transform 1 0 7084 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8188 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 9752 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9936 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10948 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11776 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13248 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_166
timestamp 1608910539
transform 1 0 16376 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1608910539
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1608910539
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1608910539
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608910539
transform 1 0 17480 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608910539
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608910539
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1608910539
transform 1 0 1472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1608910539
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2208 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608910539
transform 1 0 1656 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 3864 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608910539
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 5336 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _32_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6164 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7636 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1608910539
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9108 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 10488 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608910539
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12512 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12696 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14352 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_155
timestamp 1608910539
transform 1 0 15364 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1608910539
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_167
timestamp 1608910539
transform 1 0 16468 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1608910539
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1608910539
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1608910539
transform 1 0 1472 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1656 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2484 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5888 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5060 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 1608910539
transform 1 0 7084 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8188 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_118
timestamp 1608910539
transform 1 0 11960 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11132 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1608910539
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1608910539
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13708 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1608910539
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608910539
transform 1 0 14536 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1608910539
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_178
timestamp 1608910539
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1608910539
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608910539
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1472 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 3128 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4784 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3956 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608910539
transform 1 0 5612 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6900 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10028 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9200 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_118
timestamp 1608910539
transform 1 0 11960 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 10856 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1608910539
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_139
timestamp 1608910539
transform 1 0 13892 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13984 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1608910539
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_186
timestamp 1608910539
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1608910539
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_167
timestamp 1608910539
transform 1 0 16468 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1608910539
transform 1 0 1472 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608910539
transform 1 0 2024 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608910539
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1608910539
transform 1 0 2760 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608910539
transform 1 0 2392 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1472 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3772 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608910539
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_45
timestamp 1608910539
transform 1 0 5244 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 5612 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 6808 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5336 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608910539
transform 1 0 5244 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_82
timestamp 1608910539
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_76
timestamp 1608910539
transform 1 0 8096 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1608910539
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1608910539
transform 1 0 7912 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 7636 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 8188 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8740 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_101
timestamp 1608910539
transform 1 0 10396 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9844 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608910539
transform 1 0 9016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_113
timestamp 1608910539
transform 1 0 11500 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11776 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10856 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12604 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_126
timestamp 1608910539
transform 1 0 12696 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13156 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1608910539
transform 1 0 14076 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13984 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_158
timestamp 1608910539
transform 1 0 15640 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1608910539
transform 1 0 15456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1608910539
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1608910539
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_170
timestamp 1608910539
transform 1 0 16744 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1608910539
transform 1 0 16560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1608910539
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608910539
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608910539
transform 1 0 17848 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1608910539
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1608910539
transform 1 0 1472 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1656 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2484 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_41
timestamp 1608910539
transform 1 0 4876 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 4968 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5244 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6072 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8740 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6900 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 1608910539
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 10120 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_114
timestamp 1608910539
transform 1 0 11592 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1608910539
transform 1 0 12236 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1608910539
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13892 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_161
timestamp 1608910539
transform 1 0 15916 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1608910539
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14904 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14720 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608910539
transform 1 0 15456 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_177
timestamp 1608910539
transform 1 0 17388 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_173
timestamp 1608910539
transform 1 0 17020 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1608910539
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1608910539
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608910539
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608910539
transform 1 0 17848 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1564 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_25
timestamp 1608910539
transform 1 0 3404 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1608910539
transform 1 0 3496 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608910539
transform 1 0 4324 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608910539
transform 1 0 3036 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 8096 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608910539
transform 1 0 7636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_92
timestamp 1608910539
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9844 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1608910539
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1608910539
transform 1 0 11500 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_132
timestamp 1608910539
transform 1 0 13248 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1608910539
transform 1 0 14168 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13340 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1608910539
transform 1 0 15824 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14996 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1608910539
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1608910539
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2760 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608910539
transform 1 0 1564 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608910539
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_45
timestamp 1608910539
transform 1 0 5244 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1608910539
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5520 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 8188 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 7360 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_86
timestamp 1608910539
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10488 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1608910539
transform 1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11316 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13248 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608910539
transform 1 0 12788 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1608910539
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14904 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1608910539
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp 1608910539
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_170
timestamp 1608910539
transform 1 0 16744 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1608910539
transform 1 0 17664 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608910539
transform 1 0 17848 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_19
timestamp 1608910539
transform 1 0 2852 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3128 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4600 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608910539
transform 1 0 3956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608910539
transform 1 0 4324 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1608910539
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1608910539
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7544 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 9016 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608910539
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_106
timestamp 1608910539
transform 1 0 10856 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 11960 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11132 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13248 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14076 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_159
timestamp 1608910539
transform 1 0 15732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1608910539
transform 1 0 14904 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15824 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1608910539
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_176
timestamp 1608910539
transform 1 0 17296 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1608910539
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_10
timestamp 1608910539
transform 1 0 2024 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 1472 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 2116 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608910539
transform 1 0 1656 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4140 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5336 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1608910539
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11132 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1608910539
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_138
timestamp 1608910539
transform 1 0 13800 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14352 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12788 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1608910539
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16560 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608910539
transform 1 0 18032 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1608910539
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1608910539
transform 1 0 2852 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1932 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608910539
transform 1 0 1564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4140 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4876 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3404 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_42
timestamp 1608910539
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_74
timestamp 1608910539
transform 1 0 7912 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8188 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1608910539
transform 1 0 6900 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1608910539
transform 1 0 7636 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1608910539
transform 1 0 9016 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1608910539
transform 1 0 10304 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9844 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1608910539
transform 1 0 10028 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11960 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_127
timestamp 1608910539
transform 1 0 12788 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_141
timestamp 1608910539
transform 1 0 14076 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 12880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14168 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13340 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1608910539
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_149
timestamp 1608910539
transform 1 0 14812 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15364 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15824 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16192 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_173
timestamp 1608910539
transform 1 0 17020 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1608910539
transform 1 0 17296 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16652 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_186
timestamp 1608910539
transform 1 0 18216 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1608910539
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608910539
transform 1 0 18124 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_21
timestamp 1608910539
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3128 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 3956 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4784 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_82
timestamp 1608910539
transform 1 0 8648 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1608910539
transform 1 0 7636 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8924 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9752 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 11224 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_144
timestamp 1608910539
transform 1 0 14352 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 14444 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608910539
transform 1 0 13892 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 16100 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_15_184
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1608910539
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1608910539
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1608910539
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2116 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_38
timestamp 1608910539
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1608910539
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 3588 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_46
timestamp 1608910539
transform 1 0 5336 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5428 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1608910539
transform 1 0 6900 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7728 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1608910539
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10120 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_111
timestamp 1608910539
transform 1 0 11316 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11592 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14076 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1608910539
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15456 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_174
timestamp 1608910539
transform 1 0 17112 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1608910539
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1608910539
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 2208 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_28
timestamp 1608910539
transform 1 0 3680 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3772 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1608910539
transform 1 0 3036 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_45
timestamp 1608910539
transform 1 0 5244 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_79
timestamp 1608910539
transform 1 0 8372 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6900 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 7084 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7360 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10396 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8924 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608910539
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12512 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11224 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_138
timestamp 1608910539
transform 1 0 13800 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1608910539
transform 1 0 13524 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14260 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12696 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_152
timestamp 1608910539
transform 1 0 15088 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15180 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1608910539
transform 1 0 16008 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1608910539
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1608910539
transform 1 0 16836 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_12
timestamp 1608910539
transform 1 0 2208 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1608910539
transform 1 0 1932 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1608910539
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_24
timestamp 1608910539
transform 1 0 3312 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5704 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 6532 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_82
timestamp 1608910539
transform 1 0 8648 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 7360 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1608910539
transform 1 0 8188 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10212 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_122
timestamp 1608910539
transform 1 0 12328 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_110
timestamp 1608910539
transform 1 0 11224 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1608910539
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1608910539
transform 1 0 14260 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12696 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1608910539
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15456 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16284 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1608910539
transform 1 0 17756 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1608910539
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608910539
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608910539
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1608910539
transform 1 0 3588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4600 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4324 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_19_51
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 6072 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 7728 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6900 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7820 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_101
timestamp 1608910539
transform 1 0 10396 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_89
timestamp 1608910539
transform 1 0 9292 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1608910539
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1608910539
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1608910539
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1608910539
transform 1 0 11500 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_129
timestamp 1608910539
transform 1 0 12972 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1608910539
transform 1 0 12788 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1608910539
transform 1 0 13616 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 14444 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13064 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1608910539
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1608910539
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16100 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608910539
transform 1 0 14536 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1608910539
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_186
timestamp 1608910539
transform 1 0 18216 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1608910539
transform 1 0 17112 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1608910539
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1608910539
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1608910539
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_51
timestamp 1608910539
transform 1 0 5796 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_64
timestamp 1608910539
transform 1 0 6992 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7084 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_97
timestamp 1608910539
transform 1 0 10028 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_85
timestamp 1608910539
transform 1 0 8924 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1608910539
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_109
timestamp 1608910539
transform 1 0 11132 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_141
timestamp 1608910539
transform 1 0 14076 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1608910539
transform 1 0 12972 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 13248 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 1608910539
transform 1 0 15548 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1608910539
transform 1 0 15180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15916 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15640 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1608910539
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 17664 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1608910539
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608910539
transform 1 0 17112 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1608910539
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1608910539
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608910539
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1608910539
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608910539
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_81
timestamp 1608910539
transform 1 0 8556 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_69
timestamp 1608910539
transform 1 0 7452 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 6900 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1608910539
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1608910539
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1608910539
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1608910539
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1608910539
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_156
timestamp 1608910539
transform 1 0 15456 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1608910539
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 15732 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1608910539
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_174
timestamp 1608910539
transform 1 0 17112 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 16928 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 1122 16400 1178 17200 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 SC_IN_BOT
port 1 nsew signal input
rlabel metal2 s 3330 16400 3386 17200 6 SC_IN_TOP
port 2 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 SC_OUT_BOT
port 3 nsew signal tristate
rlabel metal2 s 5538 16400 5594 17200 6 SC_OUT_TOP
port 4 nsew signal tristate
rlabel metal2 s 1214 0 1270 800 6 bottom_grid_pin_0_
port 5 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 bottom_grid_pin_10_
port 6 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 bottom_grid_pin_11_
port 7 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 bottom_grid_pin_12_
port 8 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 bottom_grid_pin_13_
port 9 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 bottom_grid_pin_14_
port 10 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 bottom_grid_pin_15_
port 11 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_1_
port 12 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 bottom_grid_pin_2_
port 13 nsew signal tristate
rlabel metal2 s 3974 0 4030 800 6 bottom_grid_pin_3_
port 14 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 bottom_grid_pin_4_
port 15 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 bottom_grid_pin_5_
port 16 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 bottom_grid_pin_6_
port 17 nsew signal tristate
rlabel metal2 s 7562 0 7618 800 6 bottom_grid_pin_7_
port 18 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 bottom_grid_pin_8_
port 19 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 bottom_grid_pin_9_
port 20 nsew signal tristate
rlabel metal2 s 15750 0 15806 800 6 bottom_width_0_height_0__pin_0_
port 21 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 bottom_width_0_height_0__pin_1_lower
port 22 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 bottom_width_0_height_0__pin_1_upper
port 23 nsew signal tristate
rlabel metal2 s 7746 16400 7802 17200 6 ccff_head
port 24 nsew signal input
rlabel metal2 s 9954 16400 10010 17200 6 ccff_tail
port 25 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[0]
port 26 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[10]
port 27 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_in[11]
port 28 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 chanx_left_in[12]
port 29 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 chanx_left_in[13]
port 30 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 chanx_left_in[14]
port 31 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 chanx_left_in[15]
port 32 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 chanx_left_in[16]
port 33 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 chanx_left_in[17]
port 34 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 chanx_left_in[18]
port 35 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 chanx_left_in[19]
port 36 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[1]
port 37 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[2]
port 38 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[3]
port 39 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[4]
port 40 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[5]
port 41 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[6]
port 42 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[7]
port 43 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[8]
port 44 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[9]
port 45 nsew signal input
rlabel metal3 s 0 552 800 672 6 chanx_left_out[0]
port 46 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[10]
port 47 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[11]
port 48 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 chanx_left_out[12]
port 49 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[13]
port 50 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[14]
port 51 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 chanx_left_out[15]
port 52 nsew signal tristate
rlabel metal3 s 0 7216 800 7336 6 chanx_left_out[16]
port 53 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 chanx_left_out[17]
port 54 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 chanx_left_out[18]
port 55 nsew signal tristate
rlabel metal3 s 0 8440 800 8560 6 chanx_left_out[19]
port 56 nsew signal tristate
rlabel metal3 s 0 960 800 1080 6 chanx_left_out[1]
port 57 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[2]
port 58 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[3]
port 59 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 chanx_left_out[4]
port 60 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 chanx_left_out[5]
port 61 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[6]
port 62 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[7]
port 63 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_out[8]
port 64 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 chanx_left_out[9]
port 65 nsew signal tristate
rlabel metal3 s 19200 8712 20000 8832 6 chanx_right_in[0]
port 66 nsew signal input
rlabel metal3 s 19200 12928 20000 13048 6 chanx_right_in[10]
port 67 nsew signal input
rlabel metal3 s 19200 13336 20000 13456 6 chanx_right_in[11]
port 68 nsew signal input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[12]
port 69 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[13]
port 70 nsew signal input
rlabel metal3 s 19200 14696 20000 14816 6 chanx_right_in[14]
port 71 nsew signal input
rlabel metal3 s 19200 15104 20000 15224 6 chanx_right_in[15]
port 72 nsew signal input
rlabel metal3 s 19200 15512 20000 15632 6 chanx_right_in[16]
port 73 nsew signal input
rlabel metal3 s 19200 15920 20000 16040 6 chanx_right_in[17]
port 74 nsew signal input
rlabel metal3 s 19200 16328 20000 16448 6 chanx_right_in[18]
port 75 nsew signal input
rlabel metal3 s 19200 16736 20000 16856 6 chanx_right_in[19]
port 76 nsew signal input
rlabel metal3 s 19200 9120 20000 9240 6 chanx_right_in[1]
port 77 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 chanx_right_in[2]
port 78 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[3]
port 79 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[4]
port 80 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[5]
port 81 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[6]
port 82 nsew signal input
rlabel metal3 s 19200 11704 20000 11824 6 chanx_right_in[7]
port 83 nsew signal input
rlabel metal3 s 19200 12112 20000 12232 6 chanx_right_in[8]
port 84 nsew signal input
rlabel metal3 s 19200 12520 20000 12640 6 chanx_right_in[9]
port 85 nsew signal input
rlabel metal3 s 19200 144 20000 264 6 chanx_right_out[0]
port 86 nsew signal tristate
rlabel metal3 s 19200 4360 20000 4480 6 chanx_right_out[10]
port 87 nsew signal tristate
rlabel metal3 s 19200 4768 20000 4888 6 chanx_right_out[11]
port 88 nsew signal tristate
rlabel metal3 s 19200 5176 20000 5296 6 chanx_right_out[12]
port 89 nsew signal tristate
rlabel metal3 s 19200 5584 20000 5704 6 chanx_right_out[13]
port 90 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[14]
port 91 nsew signal tristate
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[15]
port 92 nsew signal tristate
rlabel metal3 s 19200 6944 20000 7064 6 chanx_right_out[16]
port 93 nsew signal tristate
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[17]
port 94 nsew signal tristate
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[18]
port 95 nsew signal tristate
rlabel metal3 s 19200 8168 20000 8288 6 chanx_right_out[19]
port 96 nsew signal tristate
rlabel metal3 s 19200 552 20000 672 6 chanx_right_out[1]
port 97 nsew signal tristate
rlabel metal3 s 19200 960 20000 1080 6 chanx_right_out[2]
port 98 nsew signal tristate
rlabel metal3 s 19200 1368 20000 1488 6 chanx_right_out[3]
port 99 nsew signal tristate
rlabel metal3 s 19200 1776 20000 1896 6 chanx_right_out[4]
port 100 nsew signal tristate
rlabel metal3 s 19200 2184 20000 2304 6 chanx_right_out[5]
port 101 nsew signal tristate
rlabel metal3 s 19200 2592 20000 2712 6 chanx_right_out[6]
port 102 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 chanx_right_out[7]
port 103 nsew signal tristate
rlabel metal3 s 19200 3544 20000 3664 6 chanx_right_out[8]
port 104 nsew signal tristate
rlabel metal3 s 19200 3952 20000 4072 6 chanx_right_out[9]
port 105 nsew signal tristate
rlabel metal2 s 14370 16400 14426 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 106 nsew signal tristate
rlabel metal2 s 16578 16400 16634 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 107 nsew signal input
rlabel metal2 s 18786 16400 18842 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 108 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 prog_clk_0_S_in
port 109 nsew signal input
rlabel metal3 s 0 144 800 264 6 prog_clk_0_W_out
port 110 nsew signal tristate
rlabel metal2 s 12162 16400 12218 17200 6 top_grid_pin_0_
port 111 nsew signal tristate
rlabel metal4 s 15771 2128 16091 14736 6 VPWR
port 112 nsew power bidirectional
rlabel metal4 s 9840 2128 10160 14736 6 VPWR
port 113 nsew power bidirectional
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 114 nsew power bidirectional
rlabel metal4 s 12805 2128 13125 14736 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
