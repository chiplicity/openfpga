* NGSPICE file created from sb_0__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt sb_0__0_ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10] chanx_right_in[11]
+ chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16]
+ chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11]
+ chanx_right_out[12] chanx_right_out[13] chanx_right_out[14] chanx_right_out[15]
+ chanx_right_out[16] chanx_right_out[17] chanx_right_out[18] chanx_right_out[19]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_top_in[0]
+ chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14]
+ chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19]
+ chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0]
+ chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14]
+ chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19]
+ chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9] prog_clk_0_E_in
+ right_bottom_grid_pin_11_ right_bottom_grid_pin_13_ right_bottom_grid_pin_15_ right_bottom_grid_pin_17_
+ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_
+ right_bottom_grid_pin_9_ top_left_grid_pin_1_ VPWR VGND
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_right_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_20.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_83_ _83_/A VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
XFILLER_3_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_66_ _66_/A VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
Xmux_right_track_36.sky130_fd_sc_hd__buf_4_0_ mux_right_track_36.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _49_/A sky130_fd_sc_hd__buf_4
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_8.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_49_ _49_/A VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_38.mux_l1_in_0_ right_bottom_grid_pin_15_ chany_top_in[18] mux_right_track_38.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_38.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_82_ chanx_right_in[6] VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_65_ _65_/A VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_right_track_26.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_right_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_48_ _48_/A VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
Xclkbuf_2_2_0_mem_right_track_0.prog_clk clkbuf_2_3_0_mem_right_track_0.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_2_0_mem_right_track_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_81_ chanx_right_in[7] VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
XFILLER_8_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_64_ _64_/A VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_right_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_47_ VGND VGND VPWR VPWR _47_/HI _47_/LO sky130_fd_sc_hd__conb_1
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_80_ chanx_right_in[8] VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_63_ _63_/A VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_0_FTB00 prog_clk_0_E_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_46_ VGND VGND VPWR VPWR _46_/HI _46_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_10.mux_l2_in_0_ _37_/HI mux_right_track_10.mux_l1_in_0_/X mux_right_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_29_ VGND VGND VPWR VPWR _29_/HI _29_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_62_ _62_/A VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_45_ VGND VGND VPWR VPWR _45_/HI _45_/LO sky130_fd_sc_hd__conb_1
X_28_ VGND VGND VPWR VPWR _28_/HI _28_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_12.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _87_/A sky130_fd_sc_hd__buf_4
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_10.mux_l1_in_0_ right_bottom_grid_pin_3_ chany_top_in[4] mux_right_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l2_in_0_ _32_/HI mux_top_track_0.mux_l1_in_0_/X mux_top_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_22.mux_l2_in_0_ _44_/HI mux_right_track_22.mux_l1_in_0_/X mux_right_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l1_in_1_ _31_/HI right_bottom_grid_pin_17_ mux_right_track_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_61_ _61_/A VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_44_ VGND VGND VPWR VPWR _44_/HI _44_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_27_ VGND VGND VPWR VPWR _27_/HI _27_/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_10.sky130_fd_sc_hd__buf_4_0_ mux_right_track_10.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _62_/A sky130_fd_sc_hd__buf_4
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_10.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l1_in_0_ right_bottom_grid_pin_1_ chany_top_in[3] mux_right_track_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_60_ _60_/A VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_18.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_22.mux_l1_in_0_ right_bottom_grid_pin_15_ chany_top_in[10] mux_right_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l1_in_0_ chanx_right_in[1] top_left_grid_pin_1_ mux_top_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_34.mux_l2_in_0_ _26_/HI mux_right_track_34.mux_l1_in_0_/X mux_right_track_34.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _63_/A sky130_fd_sc_hd__buf_4
X_43_ VGND VGND VPWR VPWR _43_/HI _43_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_26_ VGND VGND VPWR VPWR _26_/HI _26_/LO sky130_fd_sc_hd__conb_1
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _51_/A sky130_fd_sc_hd__buf_4
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_26.sky130_fd_sc_hd__buf_4_0_ mux_right_track_26.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _54_/A sky130_fd_sc_hd__buf_4
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_42_ VGND VGND VPWR VPWR _42_/HI _42_/LO sky130_fd_sc_hd__conb_1
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_30.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_34.mux_l1_in_0_ right_bottom_grid_pin_11_ chany_top_in[16] mux_right_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_25_ VGND VGND VPWR VPWR _25_/HI _25_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_41_ VGND VGND VPWR VPWR _41_/HI _41_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_28.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_24_ VGND VGND VPWR VPWR _24_/HI _24_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_36.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_mem_right_track_0.prog_clk clkbuf_2_3_0_mem_right_track_0.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_3_0_mem_right_track_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_40_ VGND VGND VPWR VPWR _40_/HI _40_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_34.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_right_track_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l2_in_1_ _29_/HI mux_right_track_4.mux_l1_in_2_/X mux_right_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_17_ right_bottom_grid_pin_13_
+ mux_right_track_4.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_right_track_4.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l2_in_0_ _40_/HI mux_right_track_16.mux_l1_in_0_/X mux_right_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_9_ right_bottom_grid_pin_5_
+ mux_right_track_4.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_22.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.mux_l1_in_0_ right_bottom_grid_pin_9_ chany_top_in[7] mux_right_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ right_bottom_grid_pin_1_ chany_top_in[1] mux_right_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_28.mux_l2_in_0_ _47_/HI mux_right_track_28.mux_l1_in_0_/X mux_right_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _65_/A sky130_fd_sc_hd__buf_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_30.mux_l2_in_0_ _24_/HI mux_right_track_30.mux_l1_in_0_/X mux_right_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_22.sky130_fd_sc_hd__buf_4_0_ mux_right_track_22.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _56_/A sky130_fd_sc_hd__buf_4
X_79_ chanx_right_in[9] VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_28.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _59_/A sky130_fd_sc_hd__buf_4
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_28.mux_l1_in_0_ right_bottom_grid_pin_5_ chany_top_in[13] mux_right_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_30.mux_l1_in_0_ right_bottom_grid_pin_7_ chany_top_in[14] mux_right_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_78_ chanx_right_in[10] VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_26.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_38.sky130_fd_sc_hd__buf_4_0_ mux_right_track_38.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _48_/A sky130_fd_sc_hd__buf_4
XFILLER_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_77_ chanx_right_in[11] VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_76_ chanx_right_in[12] VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_59_ _59_/A VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_0.mux_l2_in_1_ _36_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_14.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_2_ right_bottom_grid_pin_17_ right_bottom_grid_pin_13_
+ mux_right_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_75_ _75_/A VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xmux_top_track_24.mux_l2_in_0_ _33_/HI mux_top_track_24.mux_l1_in_0_/X mux_top_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_58_ _58_/A VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_12.mux_l2_in_0_ _38_/HI mux_right_track_12.mux_l1_in_0_/X mux_right_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_12.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_9_ right_bottom_grid_pin_5_
+ mux_right_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_74_ chanx_right_in[14] VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _75_/A sky130_fd_sc_hd__buf_4
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_57_ _57_/A VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[13] top_left_grid_pin_1_ mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _67_/A sky130_fd_sc_hd__buf_4
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_1_ chany_top_in[19] mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_12.mux_l1_in_0_ right_bottom_grid_pin_5_ chany_top_in[5] mux_right_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_73_ chanx_right_in[15] VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_56_ _56_/A VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
Xmux_right_track_24.mux_l1_in_1_ _45_/HI right_bottom_grid_pin_17_ mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_39_ VGND VGND VPWR VPWR _39_/HI _39_/LO sky130_fd_sc_hd__conb_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_12.sky130_fd_sc_hd__buf_4_0_ mux_right_track_12.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _61_/A sky130_fd_sc_hd__buf_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_72_ chanx_right_in[16] VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0_mem_right_track_0.prog_clk clkbuf_0_mem_right_track_0.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_right_track_0.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_top_track_0.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_55_ _55_/A VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_1_ chany_top_in[11] mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_36.mux_l2_in_0_ _27_/HI mux_right_track_36.mux_l1_in_0_/X mux_right_track_36.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_30.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_38_ VGND VGND VPWR VPWR _38_/HI _38_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_38.mux_l1_in_0_/S VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_34.sky130_fd_sc_hd__buf_4_0_ mux_right_track_34.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _50_/A sky130_fd_sc_hd__buf_4
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_71_ chanx_right_in[17] VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ ccff_head VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_54_ _54_/A VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xmux_right_track_28.sky130_fd_sc_hd__buf_4_0_ mux_right_track_28.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _53_/A sky130_fd_sc_hd__buf_4
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ VGND VGND VPWR VPWR _37_/HI _37_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_36.mux_l1_in_0_ right_bottom_grid_pin_13_ chany_top_in[17] mux_right_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_0_0_mem_right_track_0.prog_clk clkbuf_2_1_0_mem_right_track_0.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_0_0_mem_right_track_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_36.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_38.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_right_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_70_ chanx_right_in[18] VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_53_ _53_/A VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_36_ VGND VGND VPWR VPWR _36_/HI _36_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_52_ _52_/A VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_right_track_6.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35_ VGND VGND VPWR VPWR _35_/HI _35_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_51_ _51_/A VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34_ VGND VGND VPWR VPWR _34_/HI _34_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_1_ _30_/HI right_bottom_grid_pin_15_ mux_right_track_6.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_50_ _50_/A VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_33_ VGND VGND VPWR VPWR _33_/HI _33_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_18.mux_l2_in_0_ _41_/HI mux_right_track_18.mux_l1_in_0_/X mux_right_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_20.mux_l2_in_0_ _43_/HI mux_right_track_20.mux_l1_in_0_/X mux_right_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l1_in_1_ right_bottom_grid_pin_11_ right_bottom_grid_pin_7_
+ mux_right_track_6.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ VGND VGND VPWR VPWR _32_/HI _32_/LO sky130_fd_sc_hd__conb_1
XFILLER_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_18.mux_l1_in_0_ right_bottom_grid_pin_11_ chany_top_in[8] mux_right_track_18.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_20.mux_l1_in_0_ right_bottom_grid_pin_13_ chany_top_in[9] mux_right_track_20.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_6.mux_l1_in_0_ right_bottom_grid_pin_3_ chany_top_in[2] mux_right_track_6.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l2_in_0_ _35_/HI mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_32.mux_l2_in_0_ _25_/HI mux_right_track_32.mux_l1_in_0_/X mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_6.sky130_fd_sc_hd__buf_4_0_ mux_right_track_6.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _64_/A sky130_fd_sc_hd__buf_4
XFILLER_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _83_/A sky130_fd_sc_hd__buf_4
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31_ VGND VGND VPWR VPWR _31_/HI _31_/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_30.sky130_fd_sc_hd__buf_4_0_ mux_right_track_30.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _52_/A sky130_fd_sc_hd__buf_4
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_mem_right_track_0.prog_clk clkbuf_0_mem_right_track_0.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_right_track_0.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _55_/A sky130_fd_sc_hd__buf_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_18.sky130_fd_sc_hd__buf_4_0_ mux_right_track_18.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _58_/A sky130_fd_sc_hd__buf_4
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[5] top_left_grid_pin_1_ mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_32.mux_l1_in_0_ right_bottom_grid_pin_9_ chany_top_in[15] mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30_ VGND VGND VPWR VPWR _30_/HI _30_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_right_track_0.prog_clk/X
+ mux_right_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_16.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_mem_right_track_0.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_right_track_0.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_mem_right_track_0.prog_clk clkbuf_2_1_0_mem_right_track_0.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_1_0_mem_right_track_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_right_track_0.prog_clk/X
+ mux_right_track_14.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ _42_/HI right_bottom_grid_pin_15_ mux_right_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_87_ _87_/A VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
XFILLER_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_34.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_14.mux_l2_in_0_ _39_/HI mux_right_track_14.mux_l1_in_0_/X mux_right_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_86_ chanx_right_in[2] VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_11_ right_bottom_grid_pin_7_
+ mux_right_track_2.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_69_ chanx_right_in[19] VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_right_track_0.prog_clk/X
+ mux_right_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_right_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_85_ _85_/A VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_14.mux_l1_in_0_ right_bottom_grid_pin_7_ chany_top_in[6] mux_right_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _66_/A sky130_fd_sc_hd__buf_4
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l1_in_0_ right_bottom_grid_pin_3_ chany_top_in[0] mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_26.mux_l2_in_0_ _46_/HI mux_right_track_26.mux_l1_in_0_/X mux_right_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_0_ _34_/HI mux_top_track_4.mux_l1_in_0_/X mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_68_ chanx_right_in[0] VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _85_/A sky130_fd_sc_hd__buf_4
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_top_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_20.sky130_fd_sc_hd__buf_4_0_ mux_right_track_20.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _57_/A sky130_fd_sc_hd__buf_4
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_right_track_2.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_84_ chanx_right_in[4] VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_14.sky130_fd_sc_hd__buf_4_0_ mux_right_track_14.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _60_/A sky130_fd_sc_hd__buf_4
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_67_ _67_/A VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_0_ chanx_right_in[3] top_left_grid_pin_1_ mux_top_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_26.mux_l1_in_0_ right_bottom_grid_pin_3_ chany_top_in[12] mux_right_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_38.mux_l2_in_0_ _28_/HI mux_right_track_38.mux_l1_in_0_/X ccff_tail
+ VGND VGND VPWR VPWR mux_right_track_38.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_right_track_0.prog_clk/X
+ mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

