magic
tech EFS8A
magscale 1 2
timestamp 1603803831
<< locali >>
rect 11621 5219 11655 5321
rect 12173 4607 12207 4709
<< viali >>
rect 1593 11305 1627 11339
rect 35633 11305 35667 11339
rect 1409 11169 1443 11203
rect 35449 11169 35483 11203
rect 1593 10761 1627 10795
rect 35449 10421 35483 10455
rect 1593 10217 1627 10251
rect 35633 10217 35667 10251
rect 1409 10081 1443 10115
rect 35449 10081 35483 10115
rect 35449 9469 35483 9503
rect 1685 9333 1719 9367
rect 1593 9129 1627 9163
rect 35633 9129 35667 9163
rect 1409 8993 1443 9027
rect 2580 8993 2614 9027
rect 35449 8993 35483 9027
rect 2651 8789 2685 8823
rect 1593 8585 1627 8619
rect 2053 8585 2087 8619
rect 3433 8585 3467 8619
rect 35357 8585 35391 8619
rect 35633 8585 35667 8619
rect 2651 8517 2685 8551
rect 4675 8517 4709 8551
rect 3985 8449 4019 8483
rect 5089 8449 5123 8483
rect 1409 8381 1443 8415
rect 2329 8381 2363 8415
rect 2580 8381 2614 8415
rect 3065 8381 3099 8415
rect 3560 8381 3594 8415
rect 3663 8381 3697 8415
rect 4604 8381 4638 8415
rect 35449 8381 35483 8415
rect 36001 8381 36035 8415
rect 1593 8041 1627 8075
rect 2697 8041 2731 8075
rect 5089 8041 5123 8075
rect 5779 8041 5813 8075
rect 35633 8041 35667 8075
rect 4261 7973 4295 8007
rect 1409 7905 1443 7939
rect 2513 7905 2547 7939
rect 5708 7905 5742 7939
rect 9908 7905 9942 7939
rect 14232 7905 14266 7939
rect 19165 7905 19199 7939
rect 35449 7905 35483 7939
rect 4169 7837 4203 7871
rect 4813 7837 4847 7871
rect 3157 7701 3191 7735
rect 10011 7701 10045 7735
rect 14335 7701 14369 7735
rect 14657 7701 14691 7735
rect 19349 7701 19383 7735
rect 1593 7497 1627 7531
rect 2053 7497 2087 7531
rect 5641 7497 5675 7531
rect 13921 7497 13955 7531
rect 16635 7497 16669 7531
rect 19533 7497 19567 7531
rect 35357 7497 35391 7531
rect 35633 7497 35667 7531
rect 36737 7497 36771 7531
rect 2605 7429 2639 7463
rect 2973 7361 3007 7395
rect 4169 7361 4203 7395
rect 4721 7361 4755 7395
rect 5181 7361 5215 7395
rect 14473 7361 14507 7395
rect 1409 7293 1443 7327
rect 3801 7293 3835 7327
rect 10308 7293 10342 7327
rect 13420 7293 13454 7327
rect 16564 7293 16598 7327
rect 16957 7293 16991 7327
rect 19108 7293 19142 7327
rect 19901 7293 19935 7327
rect 20152 7293 20186 7327
rect 21465 7293 21499 7327
rect 21649 7293 21683 7327
rect 35449 7293 35483 7327
rect 36001 7293 36035 7327
rect 36553 7293 36587 7327
rect 37105 7293 37139 7327
rect 3157 7225 3191 7259
rect 3249 7225 3283 7259
rect 4813 7225 4847 7259
rect 13507 7225 13541 7259
rect 14565 7225 14599 7259
rect 15117 7225 15151 7259
rect 20637 7225 20671 7259
rect 4445 7157 4479 7191
rect 6009 7157 6043 7191
rect 9873 7157 9907 7191
rect 10379 7157 10413 7191
rect 10701 7157 10735 7191
rect 14289 7157 14323 7191
rect 15485 7157 15519 7191
rect 18981 7157 19015 7191
rect 19211 7157 19245 7191
rect 20223 7157 20257 7191
rect 20913 7157 20947 7191
rect 21833 7157 21867 7191
rect 1685 6953 1719 6987
rect 23443 6953 23477 6987
rect 2599 6885 2633 6919
rect 4261 6885 4295 6919
rect 5825 6885 5859 6919
rect 10333 6885 10367 6919
rect 10425 6885 10459 6919
rect 13829 6885 13863 6919
rect 15485 6885 15519 6919
rect 19441 6885 19475 6919
rect 21097 6885 21131 6919
rect 12684 6817 12718 6851
rect 16865 6817 16899 6851
rect 18280 6817 18314 6851
rect 23372 6817 23406 6851
rect 24501 6817 24535 6851
rect 35449 6817 35483 6851
rect 2237 6749 2271 6783
rect 4169 6749 4203 6783
rect 5089 6749 5123 6783
rect 5733 6749 5767 6783
rect 6009 6749 6043 6783
rect 6837 6749 6871 6783
rect 8585 6749 8619 6783
rect 12771 6749 12805 6783
rect 13185 6749 13219 6783
rect 13737 6749 13771 6783
rect 14013 6749 14047 6783
rect 15393 6749 15427 6783
rect 15669 6749 15703 6783
rect 19349 6749 19383 6783
rect 20637 6749 20671 6783
rect 21005 6749 21039 6783
rect 3433 6681 3467 6715
rect 4721 6681 4755 6715
rect 10885 6681 10919 6715
rect 18383 6681 18417 6715
rect 19901 6681 19935 6715
rect 21557 6681 21591 6715
rect 21925 6681 21959 6715
rect 35633 6681 35667 6715
rect 2145 6613 2179 6647
rect 3157 6613 3191 6647
rect 11345 6613 11379 6647
rect 13553 6613 13587 6647
rect 14749 6613 14783 6647
rect 15117 6613 15151 6647
rect 17049 6613 17083 6647
rect 18705 6613 18739 6647
rect 19073 6613 19107 6647
rect 20269 6613 20303 6647
rect 24593 6613 24627 6647
rect 25329 6613 25363 6647
rect 1593 6409 1627 6443
rect 3433 6409 3467 6443
rect 4077 6409 4111 6443
rect 6009 6409 6043 6443
rect 8769 6409 8803 6443
rect 10333 6409 10367 6443
rect 13001 6409 13035 6443
rect 15301 6409 15335 6443
rect 18245 6409 18279 6443
rect 18567 6409 18601 6443
rect 22385 6409 22419 6443
rect 23121 6409 23155 6443
rect 24501 6409 24535 6443
rect 2421 6341 2455 6375
rect 5273 6341 5307 6375
rect 5641 6341 5675 6375
rect 9597 6341 9631 6375
rect 11161 6341 11195 6375
rect 16037 6341 16071 6375
rect 20085 6341 20119 6375
rect 21649 6341 21683 6375
rect 24961 6341 24995 6375
rect 35449 6341 35483 6375
rect 2513 6273 2547 6307
rect 4353 6273 4387 6307
rect 4629 6273 4663 6307
rect 6929 6273 6963 6307
rect 7205 6273 7239 6307
rect 9045 6273 9079 6307
rect 10609 6273 10643 6307
rect 15485 6273 15519 6307
rect 17095 6273 17129 6307
rect 17509 6273 17543 6307
rect 19533 6273 19567 6307
rect 22017 6273 22051 6307
rect 25145 6273 25179 6307
rect 25421 6273 25455 6307
rect 1409 6205 1443 6239
rect 12265 6205 12299 6239
rect 12449 6205 12483 6239
rect 13645 6205 13679 6239
rect 17008 6205 17042 6239
rect 18464 6205 18498 6239
rect 18889 6205 18923 6239
rect 22636 6205 22670 6239
rect 2875 6137 2909 6171
rect 3801 6137 3835 6171
rect 4445 6137 4479 6171
rect 7021 6137 7055 6171
rect 9137 6137 9171 6171
rect 10701 6137 10735 6171
rect 11529 6137 11563 6171
rect 13553 6137 13587 6171
rect 14007 6137 14041 6171
rect 14933 6137 14967 6171
rect 15577 6137 15611 6171
rect 19625 6137 19659 6171
rect 20545 6137 20579 6171
rect 21097 6137 21131 6171
rect 21189 6137 21223 6171
rect 23489 6137 23523 6171
rect 25237 6137 25271 6171
rect 2053 6069 2087 6103
rect 6561 6069 6595 6103
rect 12633 6069 12667 6103
rect 14565 6069 14599 6103
rect 16405 6069 16439 6103
rect 16773 6069 16807 6103
rect 17877 6069 17911 6103
rect 19257 6069 19291 6103
rect 20821 6069 20855 6103
rect 22707 6069 22741 6103
rect 24041 6069 24075 6103
rect 6837 5865 6871 5899
rect 9045 5865 9079 5899
rect 10333 5865 10367 5899
rect 14013 5865 14047 5899
rect 14289 5865 14323 5899
rect 18429 5865 18463 5899
rect 19165 5865 19199 5899
rect 2558 5797 2592 5831
rect 3893 5797 3927 5831
rect 4398 5797 4432 5831
rect 6279 5797 6313 5831
rect 7849 5797 7883 5831
rect 10793 5797 10827 5831
rect 12817 5797 12851 5831
rect 13455 5797 13489 5831
rect 15485 5797 15519 5831
rect 16313 5797 16347 5831
rect 17830 5797 17864 5831
rect 19349 5797 19383 5831
rect 19441 5797 19475 5831
rect 21275 5797 21309 5831
rect 22569 5797 22603 5831
rect 22753 5797 22787 5831
rect 22845 5797 22879 5831
rect 24593 5797 24627 5831
rect 3157 5729 3191 5763
rect 11345 5729 11379 5763
rect 18705 5729 18739 5763
rect 26617 5729 26651 5763
rect 2237 5661 2271 5695
rect 4077 5661 4111 5695
rect 5917 5661 5951 5695
rect 7757 5661 7791 5695
rect 8033 5661 8067 5695
rect 10701 5661 10735 5695
rect 13093 5661 13127 5695
rect 14657 5661 14691 5695
rect 15393 5661 15427 5695
rect 15761 5661 15795 5695
rect 17509 5661 17543 5695
rect 20913 5661 20947 5695
rect 23029 5661 23063 5695
rect 24501 5661 24535 5695
rect 26525 5661 26559 5695
rect 27629 5661 27663 5695
rect 1777 5593 1811 5627
rect 12541 5593 12575 5627
rect 19901 5593 19935 5627
rect 25053 5593 25087 5627
rect 2145 5525 2179 5559
rect 3525 5525 3559 5559
rect 4997 5525 5031 5559
rect 7573 5525 7607 5559
rect 15025 5525 15059 5559
rect 16773 5525 16807 5559
rect 17417 5525 17451 5559
rect 20361 5525 20395 5559
rect 21833 5525 21867 5559
rect 22109 5525 22143 5559
rect 23673 5525 23707 5559
rect 25421 5525 25455 5559
rect 27905 5525 27939 5559
rect 1593 5321 1627 5355
rect 2421 5321 2455 5355
rect 5917 5321 5951 5355
rect 7389 5321 7423 5355
rect 8769 5321 8803 5355
rect 10517 5321 10551 5355
rect 10793 5321 10827 5355
rect 11161 5321 11195 5355
rect 11529 5321 11563 5355
rect 11621 5321 11655 5355
rect 12265 5321 12299 5355
rect 15669 5321 15703 5355
rect 16037 5321 16071 5355
rect 18981 5321 19015 5355
rect 20729 5321 20763 5355
rect 22937 5321 22971 5355
rect 24225 5321 24259 5355
rect 24593 5321 24627 5355
rect 27261 5321 27295 5355
rect 35633 5321 35667 5355
rect 9505 5253 9539 5287
rect 23811 5253 23845 5287
rect 2053 5185 2087 5219
rect 6837 5185 6871 5219
rect 7849 5185 7883 5219
rect 11621 5185 11655 5219
rect 21649 5185 21683 5219
rect 22293 5185 22327 5219
rect 25053 5185 25087 5219
rect 27537 5185 27571 5219
rect 1409 5117 1443 5151
rect 2513 5117 2547 5151
rect 3249 5117 3283 5151
rect 3525 5117 3559 5151
rect 3801 5117 3835 5151
rect 4997 5117 5031 5151
rect 9137 5117 9171 5151
rect 9597 5117 9631 5151
rect 11345 5117 11379 5151
rect 12541 5117 12575 5151
rect 13093 5117 13127 5151
rect 13277 5117 13311 5151
rect 13737 5117 13771 5151
rect 14749 5117 14783 5151
rect 16681 5117 16715 5151
rect 17325 5117 17359 5151
rect 18061 5117 18095 5151
rect 19809 5117 19843 5151
rect 23740 5117 23774 5151
rect 26468 5117 26502 5151
rect 26893 5117 26927 5151
rect 35449 5117 35483 5151
rect 36001 5117 36035 5151
rect 4353 5049 4387 5083
rect 4905 5049 4939 5083
rect 5359 5049 5393 5083
rect 6285 5049 6319 5083
rect 7757 5049 7791 5083
rect 8211 5049 8245 5083
rect 9959 5049 9993 5083
rect 14197 5049 14231 5083
rect 14657 5049 14691 5083
rect 15111 5049 15145 5083
rect 16405 5049 16439 5083
rect 16497 5049 16531 5083
rect 17049 5049 17083 5083
rect 17877 5049 17911 5083
rect 18423 5049 18457 5083
rect 19717 5049 19751 5083
rect 20171 5049 20205 5083
rect 21741 5049 21775 5083
rect 24777 5049 24811 5083
rect 24869 5049 24903 5083
rect 25697 5049 25731 5083
rect 27629 5049 27663 5083
rect 28181 5049 28215 5083
rect 2789 4981 2823 5015
rect 6653 4981 6687 5015
rect 11805 4981 11839 5015
rect 13645 4981 13679 5015
rect 19349 4981 19383 5015
rect 21005 4981 21039 5015
rect 21373 4981 21407 5015
rect 22661 4981 22695 5015
rect 23489 4981 23523 5015
rect 26571 4981 26605 5015
rect 1961 4777 1995 4811
rect 3801 4777 3835 4811
rect 4215 4777 4249 4811
rect 5089 4777 5123 4811
rect 5273 4777 5307 4811
rect 7665 4777 7699 4811
rect 8769 4777 8803 4811
rect 9781 4777 9815 4811
rect 15117 4777 15151 4811
rect 18061 4777 18095 4811
rect 20729 4777 20763 4811
rect 23489 4777 23523 4811
rect 24501 4777 24535 4811
rect 25513 4777 25547 4811
rect 26663 4777 26697 4811
rect 8211 4709 8245 4743
rect 12173 4709 12207 4743
rect 12265 4709 12299 4743
rect 13921 4709 13955 4743
rect 17693 4709 17727 4743
rect 19993 4709 20027 4743
rect 20269 4709 20303 4743
rect 21051 4709 21085 4743
rect 21373 4709 21407 4743
rect 24914 4709 24948 4743
rect 27629 4709 27663 4743
rect 27721 4709 27755 4743
rect 28273 4709 28307 4743
rect 1777 4641 1811 4675
rect 2421 4641 2455 4675
rect 2697 4641 2731 4675
rect 3065 4641 3099 4675
rect 4144 4641 4178 4675
rect 5181 4641 5215 4675
rect 5917 4641 5951 4675
rect 6193 4641 6227 4675
rect 6561 4641 6595 4675
rect 9965 4641 9999 4675
rect 10149 4641 10183 4675
rect 10517 4641 10551 4675
rect 10885 4641 10919 4675
rect 12449 4641 12483 4675
rect 13093 4641 13127 4675
rect 13277 4641 13311 4675
rect 13645 4641 13679 4675
rect 16221 4641 16255 4675
rect 16957 4641 16991 4675
rect 17049 4641 17083 4675
rect 17417 4641 17451 4675
rect 18521 4641 18555 4675
rect 18981 4641 19015 4675
rect 19349 4641 19383 4675
rect 19717 4641 19751 4675
rect 20964 4641 20998 4675
rect 22385 4641 22419 4675
rect 22753 4641 22787 4675
rect 23305 4641 23339 4675
rect 23581 4641 23615 4675
rect 26592 4641 26626 4675
rect 29193 4641 29227 4675
rect 30700 4641 30734 4675
rect 7849 4573 7883 4607
rect 12173 4573 12207 4607
rect 14289 4573 14323 4607
rect 15761 4573 15795 4607
rect 18429 4573 18463 4607
rect 24041 4573 24075 4607
rect 24593 4573 24627 4607
rect 27353 4505 27387 4539
rect 3525 4437 3559 4471
rect 4537 4437 4571 4471
rect 9137 4437 9171 4471
rect 11529 4437 11563 4471
rect 11897 4437 11931 4471
rect 14657 4437 14691 4471
rect 16037 4437 16071 4471
rect 21833 4437 21867 4471
rect 22201 4437 22235 4471
rect 26985 4437 27019 4471
rect 29561 4437 29595 4471
rect 30803 4437 30837 4471
rect 2237 4233 2271 4267
rect 7941 4233 7975 4267
rect 10609 4233 10643 4267
rect 15485 4233 15519 4267
rect 21281 4233 21315 4267
rect 22661 4233 22695 4267
rect 26433 4233 26467 4267
rect 28089 4233 28123 4267
rect 29101 4233 29135 4267
rect 31309 4233 31343 4267
rect 11529 4165 11563 4199
rect 4813 4097 4847 4131
rect 5457 4097 5491 4131
rect 7573 4097 7607 4131
rect 17141 4097 17175 4131
rect 19809 4097 19843 4131
rect 21925 4097 21959 4131
rect 23029 4097 23063 4131
rect 23673 4097 23707 4131
rect 30113 4097 30147 4131
rect 2421 4029 2455 4063
rect 3065 4029 3099 4063
rect 3433 4029 3467 4063
rect 3801 4029 3835 4063
rect 8401 4029 8435 4063
rect 9137 4029 9171 4063
rect 9413 4029 9447 4063
rect 9597 4029 9631 4063
rect 10885 4029 10919 4063
rect 11345 4029 11379 4063
rect 12449 4029 12483 4063
rect 13093 4029 13127 4063
rect 13277 4029 13311 4063
rect 13645 4029 13679 4063
rect 15669 4029 15703 4063
rect 16405 4029 16439 4063
rect 16681 4029 16715 4063
rect 17049 4029 17083 4063
rect 18153 4029 18187 4063
rect 18797 4029 18831 4063
rect 18889 4029 18923 4063
rect 19257 4029 19291 4063
rect 20361 4029 20395 4063
rect 22109 4029 22143 4063
rect 24593 4029 24627 4063
rect 25456 4029 25490 4063
rect 25881 4029 25915 4063
rect 26525 4029 26559 4063
rect 27445 4029 27479 4063
rect 29320 4029 29354 4063
rect 29745 4029 29779 4063
rect 4905 3961 4939 3995
rect 5733 3961 5767 3995
rect 6193 3961 6227 3995
rect 7205 3961 7239 3995
rect 14841 3961 14875 3995
rect 20269 3961 20303 3995
rect 20723 3961 20757 3995
rect 21649 3961 21683 3995
rect 23994 3961 24028 3995
rect 25237 3961 25271 3995
rect 26846 3961 26880 3995
rect 29423 3961 29457 3995
rect 30389 3961 30423 3995
rect 30481 3961 30515 3995
rect 31033 3961 31067 3995
rect 1869 3893 1903 3927
rect 2513 3893 2547 3927
rect 4261 3893 4295 3927
rect 4629 3893 4663 3927
rect 6469 3893 6503 3927
rect 8217 3893 8251 3927
rect 8493 3893 8527 3927
rect 10241 3893 10275 3927
rect 11805 3893 11839 3927
rect 12265 3893 12299 3927
rect 13645 3893 13679 3927
rect 14473 3893 14507 3927
rect 15209 3893 15243 3927
rect 17417 3893 17451 3927
rect 17785 3893 17819 3927
rect 18153 3893 18187 3927
rect 22293 3893 22327 3927
rect 23489 3893 23523 3927
rect 24869 3893 24903 3927
rect 25559 3893 25593 3927
rect 27813 3893 27847 3927
rect 1777 3689 1811 3723
rect 2651 3689 2685 3723
rect 3065 3689 3099 3723
rect 4813 3689 4847 3723
rect 5089 3689 5123 3723
rect 6653 3689 6687 3723
rect 9137 3689 9171 3723
rect 9873 3689 9907 3723
rect 12541 3689 12575 3723
rect 16313 3689 16347 3723
rect 16773 3689 16807 3723
rect 19257 3689 19291 3723
rect 20269 3689 20303 3723
rect 22017 3689 22051 3723
rect 25881 3689 25915 3723
rect 28181 3689 28215 3723
rect 30389 3689 30423 3723
rect 2145 3621 2179 3655
rect 8769 3621 8803 3655
rect 15117 3621 15151 3655
rect 15301 3621 15335 3655
rect 16037 3621 16071 3655
rect 18981 3621 19015 3655
rect 21005 3621 21039 3655
rect 21097 3621 21131 3655
rect 23949 3621 23983 3655
rect 24961 3621 24995 3655
rect 25053 3621 25087 3655
rect 26846 3621 26880 3655
rect 28365 3621 28399 3655
rect 28457 3621 28491 3655
rect 30021 3621 30055 3655
rect 30573 3621 30607 3655
rect 30665 3621 30699 3655
rect 32137 3621 32171 3655
rect 2580 3553 2614 3587
rect 3433 3553 3467 3587
rect 5273 3553 5307 3587
rect 6009 3553 6043 3587
rect 6285 3553 6319 3587
rect 6653 3553 6687 3587
rect 8677 3553 8711 3587
rect 9689 3553 9723 3587
rect 10149 3553 10183 3587
rect 11805 3553 11839 3587
rect 14289 3553 14323 3587
rect 17325 3553 17359 3587
rect 17509 3553 17543 3587
rect 17969 3553 18003 3587
rect 18337 3553 18371 3587
rect 18705 3553 18739 3587
rect 19625 3553 19659 3587
rect 22661 3553 22695 3587
rect 22937 3553 22971 3587
rect 23489 3553 23523 3587
rect 23765 3553 23799 3587
rect 32229 3553 32263 3587
rect 11897 3485 11931 3519
rect 14381 3485 14415 3519
rect 15669 3485 15703 3519
rect 19809 3485 19843 3519
rect 21281 3485 21315 3519
rect 25237 3485 25271 3519
rect 26525 3485 26559 3519
rect 29009 3485 29043 3519
rect 29285 3485 29319 3519
rect 31033 3485 31067 3519
rect 7941 3417 7975 3451
rect 11069 3417 11103 3451
rect 15439 3417 15473 3451
rect 15577 3417 15611 3451
rect 12909 3349 12943 3383
rect 13277 3349 13311 3383
rect 14749 3349 14783 3383
rect 20729 3349 20763 3383
rect 22385 3349 22419 3383
rect 24225 3349 24259 3383
rect 24593 3349 24627 3383
rect 26249 3349 26283 3383
rect 27445 3349 27479 3383
rect 33149 3349 33183 3383
rect 1777 3145 1811 3179
rect 2605 3145 2639 3179
rect 4537 3145 4571 3179
rect 7205 3145 7239 3179
rect 9781 3145 9815 3179
rect 13737 3145 13771 3179
rect 14546 3145 14580 3179
rect 14657 3145 14691 3179
rect 15485 3145 15519 3179
rect 17141 3145 17175 3179
rect 17509 3145 17543 3179
rect 19809 3145 19843 3179
rect 21097 3145 21131 3179
rect 23029 3145 23063 3179
rect 25421 3145 25455 3179
rect 27169 3145 27203 3179
rect 28549 3145 28583 3179
rect 30573 3145 30607 3179
rect 32229 3145 32263 3179
rect 2145 3077 2179 3111
rect 4077 3077 4111 3111
rect 5825 3077 5859 3111
rect 7481 3077 7515 3111
rect 22661 3077 22695 3111
rect 26065 3077 26099 3111
rect 4905 3009 4939 3043
rect 11529 3009 11563 3043
rect 12449 3009 12483 3043
rect 14749 3009 14783 3043
rect 15945 3009 15979 3043
rect 23489 3009 23523 3043
rect 26249 3009 26283 3043
rect 29285 3009 29319 3043
rect 30941 3009 30975 3043
rect 31585 3009 31619 3043
rect 32505 3009 32539 3043
rect 32781 3009 32815 3043
rect 2973 2941 3007 2975
rect 3341 2941 3375 2975
rect 3525 2941 3559 2975
rect 4077 2941 4111 2975
rect 4997 2941 5031 2975
rect 6653 2941 6687 2975
rect 7021 2941 7055 2975
rect 8033 2941 8067 2975
rect 8769 2941 8803 2975
rect 9045 2941 9079 2975
rect 9229 2941 9263 2975
rect 11161 2941 11195 2975
rect 12265 2941 12299 2975
rect 12541 2941 12575 2975
rect 14289 2941 14323 2975
rect 15853 2941 15887 2975
rect 16589 2941 16623 2975
rect 18061 2941 18095 2975
rect 18521 2941 18555 2975
rect 18889 2941 18923 2975
rect 19257 2941 19291 2975
rect 20177 2941 20211 2975
rect 20545 2941 20579 2975
rect 21557 2941 21591 2975
rect 21925 2941 21959 2975
rect 22293 2941 22327 2975
rect 22661 2941 22695 2975
rect 23673 2941 23707 2975
rect 24133 2941 24167 2975
rect 24593 2941 24627 2975
rect 24869 2941 24903 2975
rect 25145 2941 25179 2975
rect 27813 2941 27847 2975
rect 28089 2941 28123 2975
rect 29101 2941 29135 2975
rect 29377 2941 29411 2975
rect 10885 2873 10919 2907
rect 10977 2873 11011 2907
rect 11897 2873 11931 2907
rect 14381 2873 14415 2907
rect 15117 2873 15151 2907
rect 26570 2873 26604 2907
rect 31033 2873 31067 2907
rect 32597 2873 32631 2907
rect 33425 2873 33459 2907
rect 5181 2805 5215 2839
rect 5549 2805 5583 2839
rect 7941 2805 7975 2839
rect 8309 2805 8343 2839
rect 18337 2805 18371 2839
rect 27445 2805 27479 2839
rect 3065 2601 3099 2635
rect 3433 2601 3467 2635
rect 7849 2601 7883 2635
rect 8585 2601 8619 2635
rect 8861 2601 8895 2635
rect 12449 2601 12483 2635
rect 12817 2601 12851 2635
rect 13737 2601 13771 2635
rect 14933 2601 14967 2635
rect 16313 2601 16347 2635
rect 18153 2601 18187 2635
rect 19901 2601 19935 2635
rect 20223 2601 20257 2635
rect 20637 2601 20671 2635
rect 29101 2601 29135 2635
rect 29561 2601 29595 2635
rect 30941 2601 30975 2635
rect 31309 2601 31343 2635
rect 31631 2601 31665 2635
rect 32045 2601 32079 2635
rect 2789 2533 2823 2567
rect 5273 2533 5307 2567
rect 7573 2533 7607 2567
rect 11437 2533 11471 2567
rect 16865 2533 16899 2567
rect 18658 2533 18692 2567
rect 19533 2533 19567 2567
rect 21465 2533 21499 2567
rect 23121 2533 23155 2567
rect 23857 2533 23891 2567
rect 26249 2533 26283 2567
rect 26617 2533 26651 2567
rect 27214 2533 27248 2567
rect 28457 2533 28491 2567
rect 29837 2533 29871 2567
rect 29929 2533 29963 2567
rect 1777 2465 1811 2499
rect 7665 2465 7699 2499
rect 8677 2465 8711 2499
rect 9137 2465 9171 2499
rect 10793 2465 10827 2499
rect 12633 2465 12667 2499
rect 13829 2465 13863 2499
rect 13976 2465 14010 2499
rect 15485 2465 15519 2499
rect 17417 2465 17451 2499
rect 18337 2465 18371 2499
rect 20120 2465 20154 2499
rect 21005 2465 21039 2499
rect 21649 2465 21683 2499
rect 22109 2465 22143 2499
rect 22477 2465 22511 2499
rect 23029 2465 23063 2499
rect 23489 2465 23523 2499
rect 24041 2465 24075 2499
rect 24777 2465 24811 2499
rect 25053 2465 25087 2499
rect 25237 2465 25271 2499
rect 25513 2465 25547 2499
rect 26893 2465 26927 2499
rect 27813 2465 27847 2499
rect 28708 2465 28742 2499
rect 31560 2465 31594 2499
rect 32413 2465 32447 2499
rect 32689 2465 32723 2499
rect 12081 2397 12115 2431
rect 13369 2397 13403 2431
rect 14197 2397 14231 2431
rect 15301 2397 15335 2431
rect 15945 2397 15979 2431
rect 16773 2397 16807 2431
rect 25881 2397 25915 2431
rect 28089 2397 28123 2431
rect 30113 2397 30147 2431
rect 32597 2397 32631 2431
rect 34161 2397 34195 2431
rect 8217 2329 8251 2363
rect 10517 2329 10551 2363
rect 14105 2329 14139 2363
rect 15669 2329 15703 2363
rect 17693 2329 17727 2363
rect 19257 2329 19291 2363
rect 28779 2329 28813 2363
rect 14289 2261 14323 2295
<< metal1 >>
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 35618 11336 35624 11348
rect 35579 11308 35624 11336
rect 35618 11296 35624 11308
rect 35676 11296 35682 11348
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 35434 11200 35440 11212
rect 35395 11172 35440 11200
rect 35434 11160 35440 11172
rect 35492 11160 35498 11212
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1452 10764 1593 10792
rect 1452 10752 1458 10764
rect 1581 10761 1593 10764
rect 1627 10792 1639 10795
rect 2682 10792 2688 10804
rect 1627 10764 2688 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 35434 10452 35440 10464
rect 35395 10424 35440 10452
rect 35434 10412 35440 10424
rect 35492 10412 35498 10464
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 35618 10248 35624 10260
rect 35579 10220 35624 10248
rect 35618 10208 35624 10220
rect 35676 10208 35682 10260
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1670 10112 1676 10124
rect 1443 10084 1676 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 35434 10112 35440 10124
rect 35395 10084 35440 10112
rect 35434 10072 35440 10084
rect 35492 10072 35498 10124
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 35434 9500 35440 9512
rect 35395 9472 35440 9500
rect 35434 9460 35440 9472
rect 35492 9460 35498 9512
rect 1670 9364 1676 9376
rect 1631 9336 1676 9364
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1544 9132 1593 9160
rect 1544 9120 1550 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 35621 9163 35679 9169
rect 35621 9129 35633 9163
rect 35667 9160 35679 9163
rect 35710 9160 35716 9172
rect 35667 9132 35716 9160
rect 35667 9129 35679 9132
rect 35621 9123 35679 9129
rect 35710 9120 35716 9132
rect 35768 9120 35774 9172
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2038 9024 2044 9036
rect 1443 8996 2044 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 2568 9027 2626 9033
rect 2568 8993 2580 9027
rect 2614 9024 2626 9027
rect 2682 9024 2688 9036
rect 2614 8996 2688 9024
rect 2614 8993 2626 8996
rect 2568 8987 2626 8993
rect 2682 8984 2688 8996
rect 2740 9024 2746 9036
rect 3418 9024 3424 9036
rect 2740 8996 3424 9024
rect 2740 8984 2746 8996
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 35434 9024 35440 9036
rect 35395 8996 35440 9024
rect 35434 8984 35440 8996
rect 35492 8984 35498 9036
rect 2682 8829 2688 8832
rect 2639 8823 2688 8829
rect 2639 8789 2651 8823
rect 2685 8789 2688 8823
rect 2639 8783 2688 8789
rect 2682 8780 2688 8783
rect 2740 8780 2746 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1762 8616 1768 8628
rect 1627 8588 1768 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 3418 8616 3424 8628
rect 3379 8588 3424 8616
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 35345 8619 35403 8625
rect 35345 8585 35357 8619
rect 35391 8616 35403 8619
rect 35434 8616 35440 8628
rect 35391 8588 35440 8616
rect 35391 8585 35403 8588
rect 35345 8579 35403 8585
rect 35434 8576 35440 8588
rect 35492 8576 35498 8628
rect 35618 8616 35624 8628
rect 35579 8588 35624 8616
rect 35618 8576 35624 8588
rect 35676 8576 35682 8628
rect 2590 8508 2596 8560
rect 2648 8557 2654 8560
rect 2648 8551 2697 8557
rect 2648 8517 2651 8551
rect 2685 8517 2697 8551
rect 2648 8511 2697 8517
rect 4663 8551 4721 8557
rect 4663 8517 4675 8551
rect 4709 8548 4721 8551
rect 5442 8548 5448 8560
rect 4709 8520 5448 8548
rect 4709 8517 4721 8520
rect 4663 8511 4721 8517
rect 2648 8508 2654 8511
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 3970 8480 3976 8492
rect 3528 8452 3976 8480
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2317 8415 2375 8421
rect 2317 8412 2329 8415
rect 1443 8384 2329 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2317 8381 2329 8384
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 2568 8415 2626 8421
rect 2568 8381 2580 8415
rect 2614 8412 2626 8415
rect 2866 8412 2872 8424
rect 2614 8384 2872 8412
rect 2614 8381 2626 8384
rect 2568 8375 2626 8381
rect 2332 8344 2360 8375
rect 2866 8372 2872 8384
rect 2924 8412 2930 8424
rect 3050 8412 3056 8424
rect 2924 8384 3056 8412
rect 2924 8372 2930 8384
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 3528 8421 3556 8452
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 5074 8480 5080 8492
rect 5035 8452 5080 8480
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 3528 8415 3606 8421
rect 3528 8384 3560 8415
rect 3548 8381 3560 8384
rect 3594 8381 3606 8415
rect 3548 8375 3606 8381
rect 3651 8415 3709 8421
rect 3651 8381 3663 8415
rect 3697 8412 3709 8415
rect 4062 8412 4068 8424
rect 3697 8384 4068 8412
rect 3697 8381 3709 8384
rect 3651 8375 3709 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4592 8415 4650 8421
rect 4592 8412 4604 8415
rect 4356 8384 4604 8412
rect 4356 8344 4384 8384
rect 4592 8381 4604 8384
rect 4638 8412 4650 8415
rect 5092 8412 5120 8440
rect 35434 8412 35440 8424
rect 4638 8384 5120 8412
rect 35395 8384 35440 8412
rect 4638 8381 4650 8384
rect 4592 8375 4650 8381
rect 35434 8372 35440 8384
rect 35492 8412 35498 8424
rect 35989 8415 36047 8421
rect 35989 8412 36001 8415
rect 35492 8384 36001 8412
rect 35492 8372 35498 8384
rect 35989 8381 36001 8384
rect 36035 8381 36047 8415
rect 35989 8375 36047 8381
rect 2332 8316 4384 8344
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 2498 8032 2504 8084
rect 2556 8072 2562 8084
rect 2685 8075 2743 8081
rect 2685 8072 2697 8075
rect 2556 8044 2697 8072
rect 2556 8032 2562 8044
rect 2685 8041 2697 8044
rect 2731 8041 2743 8075
rect 5074 8072 5080 8084
rect 5035 8044 5080 8072
rect 2685 8035 2743 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5767 8075 5825 8081
rect 5767 8041 5779 8075
rect 5813 8072 5825 8075
rect 6638 8072 6644 8084
rect 5813 8044 6644 8072
rect 5813 8041 5825 8044
rect 5767 8035 5825 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 35526 8032 35532 8084
rect 35584 8072 35590 8084
rect 35621 8075 35679 8081
rect 35621 8072 35633 8075
rect 35584 8044 35633 8072
rect 35584 8032 35590 8044
rect 35621 8041 35633 8044
rect 35667 8041 35679 8075
rect 35621 8035 35679 8041
rect 4246 8004 4252 8016
rect 4207 7976 4252 8004
rect 4246 7964 4252 7976
rect 4304 7964 4310 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 2038 7936 2044 7948
rect 1443 7908 2044 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 2498 7936 2504 7948
rect 2459 7908 2504 7936
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 5696 7939 5754 7945
rect 5696 7905 5708 7939
rect 5742 7936 5754 7939
rect 5902 7936 5908 7948
rect 5742 7908 5908 7936
rect 5742 7905 5754 7908
rect 5696 7899 5754 7905
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 9858 7896 9864 7948
rect 9916 7945 9922 7948
rect 9916 7939 9954 7945
rect 9942 7905 9954 7939
rect 9916 7899 9954 7905
rect 9916 7896 9922 7899
rect 14182 7896 14188 7948
rect 14240 7945 14246 7948
rect 14240 7939 14278 7945
rect 14266 7905 14278 7939
rect 19150 7936 19156 7948
rect 19111 7908 19156 7936
rect 14240 7899 14278 7905
rect 14240 7896 14246 7899
rect 19150 7896 19156 7908
rect 19208 7896 19214 7948
rect 35434 7936 35440 7948
rect 35395 7908 35440 7936
rect 35434 7896 35440 7908
rect 35492 7896 35498 7948
rect 4154 7868 4160 7880
rect 4115 7840 4160 7868
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 5166 7868 5172 7880
rect 4847 7840 5172 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 3142 7732 3148 7744
rect 3103 7704 3148 7732
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 9999 7735 10057 7741
rect 9999 7701 10011 7735
rect 10045 7732 10057 7735
rect 10318 7732 10324 7744
rect 10045 7704 10324 7732
rect 10045 7701 10057 7704
rect 9999 7695 10057 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 14323 7735 14381 7741
rect 14323 7701 14335 7735
rect 14369 7732 14381 7735
rect 14458 7732 14464 7744
rect 14369 7704 14464 7732
rect 14369 7701 14381 7704
rect 14323 7695 14381 7701
rect 14458 7692 14464 7704
rect 14516 7732 14522 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14516 7704 14657 7732
rect 14516 7692 14522 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 14645 7695 14703 7701
rect 19337 7735 19395 7741
rect 19337 7701 19349 7735
rect 19383 7732 19395 7735
rect 20438 7732 20444 7744
rect 19383 7704 20444 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 1854 7528 1860 7540
rect 1627 7500 1860 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 1854 7488 1860 7500
rect 1912 7488 1918 7540
rect 2038 7528 2044 7540
rect 1999 7500 2044 7528
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 5629 7531 5687 7537
rect 5629 7528 5641 7531
rect 4212 7500 5641 7528
rect 4212 7488 4218 7500
rect 5629 7497 5641 7500
rect 5675 7497 5687 7531
rect 5629 7491 5687 7497
rect 13909 7531 13967 7537
rect 13909 7497 13921 7531
rect 13955 7528 13967 7531
rect 14366 7528 14372 7540
rect 13955 7500 14372 7528
rect 13955 7497 13967 7500
rect 13909 7491 13967 7497
rect 2498 7420 2504 7472
rect 2556 7460 2562 7472
rect 2593 7463 2651 7469
rect 2593 7460 2605 7463
rect 2556 7432 2605 7460
rect 2556 7420 2562 7432
rect 2593 7429 2605 7432
rect 2639 7460 2651 7463
rect 3694 7460 3700 7472
rect 2639 7432 3700 7460
rect 2639 7429 2651 7432
rect 2593 7423 2651 7429
rect 3694 7420 3700 7432
rect 3752 7420 3758 7472
rect 5074 7460 5080 7472
rect 4724 7432 5080 7460
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3234 7392 3240 7404
rect 3007 7364 3240 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3234 7352 3240 7364
rect 3292 7392 3298 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3292 7364 4169 7392
rect 3292 7352 3298 7364
rect 4157 7361 4169 7364
rect 4203 7392 4215 7395
rect 4246 7392 4252 7404
rect 4203 7364 4252 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 4724 7401 4752 7432
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 5166 7392 5172 7404
rect 5127 7364 5172 7392
rect 4709 7355 4767 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 1670 7324 1676 7336
rect 1443 7296 1676 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7324 3847 7327
rect 4430 7324 4436 7336
rect 3835 7296 4436 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 10296 7327 10354 7333
rect 10296 7293 10308 7327
rect 10342 7324 10354 7327
rect 10342 7296 10732 7324
rect 10342 7293 10354 7296
rect 10296 7287 10354 7293
rect 3142 7256 3148 7268
rect 3055 7228 3148 7256
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 4801 7259 4859 7265
rect 3292 7228 3337 7256
rect 3292 7216 3298 7228
rect 4801 7225 4813 7259
rect 4847 7225 4859 7259
rect 4801 7219 4859 7225
rect 3160 7188 3188 7216
rect 3970 7188 3976 7200
rect 3160 7160 3976 7188
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 4212 7160 4445 7188
rect 4212 7148 4218 7160
rect 4433 7157 4445 7160
rect 4479 7188 4491 7191
rect 4816 7188 4844 7219
rect 10704 7200 10732 7296
rect 13078 7284 13084 7336
rect 13136 7324 13142 7336
rect 13408 7327 13466 7333
rect 13408 7324 13420 7327
rect 13136 7296 13420 7324
rect 13136 7284 13142 7296
rect 13408 7293 13420 7296
rect 13454 7324 13466 7327
rect 13924 7324 13952 7491
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 16666 7537 16672 7540
rect 16623 7531 16672 7537
rect 16623 7497 16635 7531
rect 16669 7497 16672 7531
rect 16623 7491 16672 7497
rect 16666 7488 16672 7491
rect 16724 7488 16730 7540
rect 19150 7488 19156 7540
rect 19208 7528 19214 7540
rect 19521 7531 19579 7537
rect 19521 7528 19533 7531
rect 19208 7500 19533 7528
rect 19208 7488 19214 7500
rect 19521 7497 19533 7500
rect 19567 7528 19579 7531
rect 19794 7528 19800 7540
rect 19567 7500 19800 7528
rect 19567 7497 19579 7500
rect 19521 7491 19579 7497
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 35345 7531 35403 7537
rect 35345 7497 35357 7531
rect 35391 7528 35403 7531
rect 35434 7528 35440 7540
rect 35391 7500 35440 7528
rect 35391 7497 35403 7500
rect 35345 7491 35403 7497
rect 35434 7488 35440 7500
rect 35492 7488 35498 7540
rect 35621 7531 35679 7537
rect 35621 7497 35633 7531
rect 35667 7528 35679 7531
rect 35802 7528 35808 7540
rect 35667 7500 35808 7528
rect 35667 7497 35679 7500
rect 35621 7491 35679 7497
rect 35802 7488 35808 7500
rect 35860 7488 35866 7540
rect 36722 7528 36728 7540
rect 36683 7500 36728 7528
rect 36722 7488 36728 7500
rect 36780 7488 36786 7540
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 13454 7296 13952 7324
rect 16552 7327 16610 7333
rect 13454 7293 13466 7296
rect 13408 7287 13466 7293
rect 16552 7293 16564 7327
rect 16598 7324 16610 7327
rect 16666 7324 16672 7336
rect 16598 7296 16672 7324
rect 16598 7293 16610 7296
rect 16552 7287 16610 7293
rect 16666 7284 16672 7296
rect 16724 7324 16730 7336
rect 16945 7327 17003 7333
rect 16945 7324 16957 7327
rect 16724 7296 16957 7324
rect 16724 7284 16730 7296
rect 16945 7293 16957 7296
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 19058 7284 19064 7336
rect 19116 7333 19122 7336
rect 19116 7327 19154 7333
rect 19142 7324 19154 7327
rect 19886 7324 19892 7336
rect 19142 7296 19892 7324
rect 19142 7293 19154 7296
rect 19116 7287 19154 7293
rect 19116 7284 19122 7287
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 19978 7284 19984 7336
rect 20036 7324 20042 7336
rect 20140 7327 20198 7333
rect 20140 7324 20152 7327
rect 20036 7296 20152 7324
rect 20036 7284 20042 7296
rect 20140 7293 20152 7296
rect 20186 7293 20198 7327
rect 20140 7287 20198 7293
rect 21453 7327 21511 7333
rect 21453 7293 21465 7327
rect 21499 7324 21511 7327
rect 21634 7324 21640 7336
rect 21499 7296 21640 7324
rect 21499 7293 21511 7296
rect 21453 7287 21511 7293
rect 13495 7259 13553 7265
rect 13495 7225 13507 7259
rect 13541 7256 13553 7259
rect 13722 7256 13728 7268
rect 13541 7228 13728 7256
rect 13541 7225 13553 7228
rect 13495 7219 13553 7225
rect 13722 7216 13728 7228
rect 13780 7216 13786 7268
rect 14553 7259 14611 7265
rect 14553 7225 14565 7259
rect 14599 7256 14611 7259
rect 14826 7256 14832 7268
rect 14599 7228 14832 7256
rect 14599 7225 14611 7228
rect 14553 7219 14611 7225
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 15105 7259 15163 7265
rect 15105 7225 15117 7259
rect 15151 7225 15163 7259
rect 20155 7256 20183 7287
rect 21634 7284 21640 7296
rect 21692 7284 21698 7336
rect 34974 7284 34980 7336
rect 35032 7324 35038 7336
rect 35437 7327 35495 7333
rect 35437 7324 35449 7327
rect 35032 7296 35449 7324
rect 35032 7284 35038 7296
rect 35437 7293 35449 7296
rect 35483 7324 35495 7327
rect 35989 7327 36047 7333
rect 35989 7324 36001 7327
rect 35483 7296 36001 7324
rect 35483 7293 35495 7296
rect 35437 7287 35495 7293
rect 35989 7293 36001 7296
rect 36035 7293 36047 7327
rect 36538 7324 36544 7336
rect 36499 7296 36544 7324
rect 35989 7287 36047 7293
rect 36538 7284 36544 7296
rect 36596 7324 36602 7336
rect 37093 7327 37151 7333
rect 37093 7324 37105 7327
rect 36596 7296 37105 7324
rect 36596 7284 36602 7296
rect 37093 7293 37105 7296
rect 37139 7293 37151 7327
rect 37093 7287 37151 7293
rect 20625 7259 20683 7265
rect 20625 7256 20637 7259
rect 20155 7228 20637 7256
rect 15105 7219 15163 7225
rect 20625 7225 20637 7228
rect 20671 7256 20683 7259
rect 23014 7256 23020 7268
rect 20671 7228 23020 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 4479 7160 4844 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 5902 7148 5908 7200
rect 5960 7188 5966 7200
rect 5997 7191 6055 7197
rect 5997 7188 6009 7191
rect 5960 7160 6009 7188
rect 5960 7148 5966 7160
rect 5997 7157 6009 7160
rect 6043 7157 6055 7191
rect 9858 7188 9864 7200
rect 9819 7160 9864 7188
rect 5997 7151 6055 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10367 7191 10425 7197
rect 10367 7157 10379 7191
rect 10413 7188 10425 7191
rect 10502 7188 10508 7200
rect 10413 7160 10508 7188
rect 10413 7157 10425 7160
rect 10367 7151 10425 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10686 7188 10692 7200
rect 10647 7160 10692 7188
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 14277 7191 14335 7197
rect 14277 7188 14289 7191
rect 14240 7160 14289 7188
rect 14240 7148 14246 7160
rect 14277 7157 14289 7160
rect 14323 7188 14335 7191
rect 15010 7188 15016 7200
rect 14323 7160 15016 7188
rect 14323 7157 14335 7160
rect 14277 7151 14335 7157
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15120 7188 15148 7219
rect 23014 7216 23020 7228
rect 23072 7216 23078 7268
rect 15473 7191 15531 7197
rect 15473 7188 15485 7191
rect 15120 7160 15485 7188
rect 15473 7157 15485 7160
rect 15519 7188 15531 7191
rect 15562 7188 15568 7200
rect 15519 7160 15568 7188
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 18966 7188 18972 7200
rect 18927 7160 18972 7188
rect 18966 7148 18972 7160
rect 19024 7148 19030 7200
rect 19242 7197 19248 7200
rect 19199 7191 19248 7197
rect 19199 7157 19211 7191
rect 19245 7157 19248 7191
rect 19199 7151 19248 7157
rect 19242 7148 19248 7151
rect 19300 7148 19306 7200
rect 20162 7148 20168 7200
rect 20220 7197 20226 7200
rect 20220 7191 20269 7197
rect 20220 7157 20223 7191
rect 20257 7157 20269 7191
rect 20898 7188 20904 7200
rect 20859 7160 20904 7188
rect 20220 7151 20269 7157
rect 20220 7148 20226 7151
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 21821 7191 21879 7197
rect 21821 7157 21833 7191
rect 21867 7188 21879 7191
rect 21910 7188 21916 7200
rect 21867 7160 21916 7188
rect 21867 7157 21879 7160
rect 21821 7151 21879 7157
rect 21910 7148 21916 7160
rect 21968 7148 21974 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 1670 6984 1676 6996
rect 1583 6956 1676 6984
rect 1670 6944 1676 6956
rect 1728 6984 1734 6996
rect 9490 6984 9496 6996
rect 1728 6956 9496 6984
rect 1728 6944 1734 6956
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 9732 6956 16988 6984
rect 9732 6944 9738 6956
rect 2587 6919 2645 6925
rect 2587 6885 2599 6919
rect 2633 6885 2645 6919
rect 4246 6916 4252 6928
rect 4207 6888 4252 6916
rect 2587 6879 2645 6885
rect 2406 6808 2412 6860
rect 2464 6848 2470 6860
rect 2608 6848 2636 6879
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 5166 6876 5172 6928
rect 5224 6916 5230 6928
rect 5810 6916 5816 6928
rect 5224 6888 5488 6916
rect 5771 6888 5816 6916
rect 5224 6876 5230 6888
rect 2464 6820 2636 6848
rect 5460 6848 5488 6888
rect 5810 6876 5816 6888
rect 5868 6876 5874 6928
rect 10318 6916 10324 6928
rect 10279 6888 10324 6916
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 10410 6876 10416 6928
rect 10468 6916 10474 6928
rect 13817 6919 13875 6925
rect 10468 6888 10513 6916
rect 10468 6876 10474 6888
rect 13817 6885 13829 6919
rect 13863 6916 13875 6919
rect 15470 6916 15476 6928
rect 13863 6888 14412 6916
rect 13863 6885 13875 6888
rect 13817 6879 13875 6885
rect 12672 6851 12730 6857
rect 5460 6820 5580 6848
rect 2464 6808 2470 6820
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 2240 6644 2268 6743
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3936 6752 4169 6780
rect 3936 6740 3942 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4396 6752 5089 6780
rect 4396 6740 4402 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 2774 6672 2780 6724
rect 2832 6712 2838 6724
rect 3421 6715 3479 6721
rect 3421 6712 3433 6715
rect 2832 6684 3433 6712
rect 2832 6672 2838 6684
rect 3421 6681 3433 6684
rect 3467 6681 3479 6715
rect 3421 6675 3479 6681
rect 4430 6672 4436 6724
rect 4488 6712 4494 6724
rect 4709 6715 4767 6721
rect 4709 6712 4721 6715
rect 4488 6684 4721 6712
rect 4488 6672 4494 6684
rect 4709 6681 4721 6684
rect 4755 6681 4767 6715
rect 5552 6712 5580 6820
rect 12672 6817 12684 6851
rect 12718 6848 12730 6851
rect 12986 6848 12992 6860
rect 12718 6820 12992 6848
rect 12718 6817 12730 6820
rect 12672 6811 12730 6817
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 14384 6848 14412 6888
rect 15212 6888 15476 6916
rect 15212 6848 15240 6888
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 14384 6820 15240 6848
rect 5718 6780 5724 6792
rect 5679 6752 5724 6780
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6043 6752 6837 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6825 6749 6837 6752
rect 6871 6780 6883 6783
rect 6914 6780 6920 6792
rect 6871 6752 6920 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 6012 6712 6040 6743
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 8754 6780 8760 6792
rect 8619 6752 8760 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 12759 6783 12817 6789
rect 12759 6749 12771 6783
rect 12805 6780 12817 6783
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 12805 6752 13185 6780
rect 12805 6749 12817 6752
rect 12759 6743 12817 6749
rect 13173 6749 13185 6752
rect 13219 6780 13231 6783
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 13219 6752 13737 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 13998 6780 14004 6792
rect 13959 6752 14004 6780
rect 13725 6743 13783 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 14384 6780 14412 6820
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 16853 6851 16911 6857
rect 16853 6848 16865 6851
rect 16632 6820 16865 6848
rect 16632 6808 16638 6820
rect 16853 6817 16865 6820
rect 16899 6817 16911 6851
rect 16960 6848 16988 6956
rect 23382 6944 23388 6996
rect 23440 6993 23446 6996
rect 23440 6987 23489 6993
rect 23440 6953 23443 6987
rect 23477 6953 23489 6987
rect 23440 6947 23489 6953
rect 23440 6944 23446 6947
rect 19429 6919 19487 6925
rect 19429 6916 19441 6919
rect 19168 6888 19441 6916
rect 18230 6848 18236 6860
rect 18288 6857 18294 6860
rect 18288 6851 18326 6857
rect 16960 6820 18236 6848
rect 16853 6811 16911 6817
rect 18230 6808 18236 6820
rect 18314 6817 18326 6851
rect 18288 6811 18326 6817
rect 18288 6808 18294 6811
rect 19058 6808 19064 6860
rect 19116 6848 19122 6860
rect 19168 6848 19196 6888
rect 19429 6885 19441 6888
rect 19475 6885 19487 6919
rect 21085 6919 21143 6925
rect 21085 6916 21097 6919
rect 19429 6879 19487 6885
rect 20824 6888 21097 6916
rect 19116 6820 19196 6848
rect 19116 6808 19122 6820
rect 20714 6808 20720 6860
rect 20772 6848 20778 6860
rect 20824 6848 20852 6888
rect 21085 6885 21097 6888
rect 21131 6885 21143 6919
rect 21085 6879 21143 6885
rect 20772 6820 20852 6848
rect 23360 6851 23418 6857
rect 20772 6808 20778 6820
rect 23360 6817 23372 6851
rect 23406 6848 23418 6851
rect 23474 6848 23480 6860
rect 23406 6820 23480 6848
rect 23406 6817 23418 6820
rect 23360 6811 23418 6817
rect 23474 6808 23480 6820
rect 23532 6808 23538 6860
rect 24486 6848 24492 6860
rect 24447 6820 24492 6848
rect 24486 6808 24492 6820
rect 24544 6808 24550 6860
rect 35434 6848 35440 6860
rect 35395 6820 35440 6848
rect 35434 6808 35440 6820
rect 35492 6808 35498 6860
rect 15378 6780 15384 6792
rect 14148 6752 14412 6780
rect 15339 6752 15384 6780
rect 14148 6740 14154 6752
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 15657 6783 15715 6789
rect 15657 6780 15669 6783
rect 15620 6752 15669 6780
rect 15620 6740 15626 6752
rect 15657 6749 15669 6752
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 19337 6783 19395 6789
rect 19337 6780 19349 6783
rect 18656 6752 19349 6780
rect 18656 6740 18662 6752
rect 19337 6749 19349 6752
rect 19383 6780 19395 6783
rect 20625 6783 20683 6789
rect 20625 6780 20637 6783
rect 19383 6752 20637 6780
rect 19383 6749 19395 6752
rect 19337 6743 19395 6749
rect 20625 6749 20637 6752
rect 20671 6749 20683 6783
rect 20625 6743 20683 6749
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20864 6752 21005 6780
rect 20864 6740 20870 6752
rect 20993 6749 21005 6752
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 5552 6684 6040 6712
rect 10873 6715 10931 6721
rect 4709 6675 4767 6681
rect 10873 6681 10885 6715
rect 10919 6681 10931 6715
rect 10873 6675 10931 6681
rect 18371 6715 18429 6721
rect 18371 6681 18383 6715
rect 18417 6712 18429 6715
rect 18966 6712 18972 6724
rect 18417 6684 18972 6712
rect 18417 6681 18429 6684
rect 18371 6675 18429 6681
rect 2498 6644 2504 6656
rect 2179 6616 2504 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 4062 6644 4068 6656
rect 3191 6616 4068 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 10888 6644 10916 6675
rect 18966 6672 18972 6684
rect 19024 6672 19030 6724
rect 19886 6712 19892 6724
rect 19847 6684 19892 6712
rect 19886 6672 19892 6684
rect 19944 6712 19950 6724
rect 20898 6712 20904 6724
rect 19944 6684 20904 6712
rect 19944 6672 19950 6684
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 21542 6712 21548 6724
rect 21503 6684 21548 6712
rect 21542 6672 21548 6684
rect 21600 6712 21606 6724
rect 21913 6715 21971 6721
rect 21913 6712 21925 6715
rect 21600 6684 21925 6712
rect 21600 6672 21606 6684
rect 21913 6681 21925 6684
rect 21959 6681 21971 6715
rect 21913 6675 21971 6681
rect 35250 6672 35256 6724
rect 35308 6712 35314 6724
rect 35621 6715 35679 6721
rect 35621 6712 35633 6715
rect 35308 6684 35633 6712
rect 35308 6672 35314 6684
rect 35621 6681 35633 6684
rect 35667 6681 35679 6715
rect 35621 6675 35679 6681
rect 11330 6644 11336 6656
rect 10652 6616 11336 6644
rect 10652 6604 10658 6616
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13630 6644 13636 6656
rect 13587 6616 13636 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6644 14795 6647
rect 14826 6644 14832 6656
rect 14783 6616 14832 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15102 6644 15108 6656
rect 15063 6616 15108 6644
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 17034 6644 17040 6656
rect 16995 6616 17040 6644
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19058 6644 19064 6656
rect 19019 6616 19064 6644
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 20162 6644 20168 6656
rect 19392 6616 20168 6644
rect 19392 6604 19398 6616
rect 20162 6604 20168 6616
rect 20220 6644 20226 6656
rect 20257 6647 20315 6653
rect 20257 6644 20269 6647
rect 20220 6616 20269 6644
rect 20220 6604 20226 6616
rect 20257 6613 20269 6616
rect 20303 6613 20315 6647
rect 24578 6644 24584 6656
rect 24539 6616 24584 6644
rect 20257 6607 20315 6613
rect 24578 6604 24584 6616
rect 24636 6604 24642 6656
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25317 6647 25375 6653
rect 25317 6644 25329 6647
rect 24912 6616 25329 6644
rect 24912 6604 24918 6616
rect 25317 6613 25329 6616
rect 25363 6613 25375 6647
rect 25317 6607 25375 6613
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1946 6440 1952 6452
rect 1627 6412 1952 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 3292 6412 3433 6440
rect 3292 6400 3298 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 4062 6440 4068 6452
rect 4023 6412 4068 6440
rect 3421 6403 3479 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5776 6412 6009 6440
rect 5776 6400 5782 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 8754 6440 8760 6452
rect 8715 6412 8760 6440
rect 5997 6403 6055 6409
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 10321 6443 10379 6449
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 10410 6440 10416 6452
rect 10367 6412 10416 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 12986 6440 12992 6452
rect 12947 6412 12992 6440
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 15289 6443 15347 6449
rect 15289 6409 15301 6443
rect 15335 6440 15347 6443
rect 15470 6440 15476 6452
rect 15335 6412 15476 6440
rect 15335 6409 15347 6412
rect 15289 6403 15347 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 18230 6440 18236 6452
rect 18191 6412 18236 6440
rect 18230 6400 18236 6412
rect 18288 6400 18294 6452
rect 18598 6449 18604 6452
rect 18555 6443 18604 6449
rect 18555 6409 18567 6443
rect 18601 6409 18604 6443
rect 18555 6403 18604 6409
rect 18598 6400 18604 6403
rect 18656 6400 18662 6452
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 22373 6443 22431 6449
rect 22373 6440 22385 6443
rect 21324 6412 22385 6440
rect 21324 6400 21330 6412
rect 22373 6409 22385 6412
rect 22419 6409 22431 6443
rect 22373 6403 22431 6409
rect 23109 6443 23167 6449
rect 23109 6409 23121 6443
rect 23155 6440 23167 6443
rect 23290 6440 23296 6452
rect 23155 6412 23296 6440
rect 23155 6409 23167 6412
rect 23109 6403 23167 6409
rect 2406 6372 2412 6384
rect 2367 6344 2412 6372
rect 2406 6332 2412 6344
rect 2464 6332 2470 6384
rect 4246 6332 4252 6384
rect 4304 6372 4310 6384
rect 5261 6375 5319 6381
rect 5261 6372 5273 6375
rect 4304 6344 5273 6372
rect 4304 6332 4310 6344
rect 5261 6341 5273 6344
rect 5307 6372 5319 6375
rect 5629 6375 5687 6381
rect 5629 6372 5641 6375
rect 5307 6344 5641 6372
rect 5307 6341 5319 6344
rect 5261 6335 5319 6341
rect 5629 6341 5641 6344
rect 5675 6372 5687 6375
rect 5810 6372 5816 6384
rect 5675 6344 5816 6372
rect 5675 6341 5687 6344
rect 5629 6335 5687 6341
rect 5810 6332 5816 6344
rect 5868 6332 5874 6384
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6304 2559 6307
rect 2774 6304 2780 6316
rect 2547 6276 2780 6304
rect 2547 6273 2559 6276
rect 2501 6267 2559 6273
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 4338 6304 4344 6316
rect 4299 6276 4344 6304
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4430 6264 4436 6316
rect 4488 6304 4494 6316
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4488 6276 4629 6304
rect 4488 6264 4494 6276
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 6914 6304 6920 6316
rect 6875 6276 6920 6304
rect 4617 6267 4675 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7190 6304 7196 6316
rect 7151 6276 7196 6304
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 8772 6304 8800 6400
rect 9585 6375 9643 6381
rect 9585 6341 9597 6375
rect 9631 6372 9643 6375
rect 11146 6372 11152 6384
rect 9631 6344 11152 6372
rect 9631 6341 9643 6344
rect 9585 6335 9643 6341
rect 11146 6332 11152 6344
rect 11204 6332 11210 6384
rect 13998 6332 14004 6384
rect 14056 6372 14062 6384
rect 16025 6375 16083 6381
rect 16025 6372 16037 6375
rect 14056 6344 16037 6372
rect 14056 6332 14062 6344
rect 16025 6341 16037 6344
rect 16071 6341 16083 6375
rect 16025 6335 16083 6341
rect 20073 6375 20131 6381
rect 20073 6341 20085 6375
rect 20119 6372 20131 6375
rect 21542 6372 21548 6384
rect 20119 6344 21548 6372
rect 20119 6341 20131 6344
rect 20073 6335 20131 6341
rect 21542 6332 21548 6344
rect 21600 6372 21606 6384
rect 21637 6375 21695 6381
rect 21637 6372 21649 6375
rect 21600 6344 21649 6372
rect 21600 6332 21606 6344
rect 21637 6341 21649 6344
rect 21683 6341 21695 6375
rect 21637 6335 21695 6341
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 8772 6276 9045 6304
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 10594 6304 10600 6316
rect 10555 6276 10600 6304
rect 9033 6267 9091 6273
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 15473 6307 15531 6313
rect 15473 6304 15485 6307
rect 15160 6276 15485 6304
rect 15160 6264 15166 6276
rect 15473 6273 15485 6276
rect 15519 6304 15531 6307
rect 17083 6307 17141 6313
rect 17083 6304 17095 6307
rect 15519 6276 17095 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 17083 6273 17095 6276
rect 17129 6273 17141 6307
rect 17494 6304 17500 6316
rect 17455 6276 17500 6304
rect 17083 6267 17141 6273
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19521 6307 19579 6313
rect 19521 6304 19533 6307
rect 19024 6276 19533 6304
rect 19024 6264 19030 6276
rect 19521 6273 19533 6276
rect 19567 6273 19579 6307
rect 19521 6267 19579 6273
rect 20806 6264 20812 6316
rect 20864 6304 20870 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 20864 6276 22017 6304
rect 20864 6264 20870 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 12253 6239 12311 6245
rect 1443 6208 2084 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2056 6112 2084 6208
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 12434 6236 12440 6248
rect 12299 6208 12440 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 12434 6196 12440 6208
rect 12492 6236 12498 6248
rect 13630 6236 13636 6248
rect 12492 6208 12537 6236
rect 13591 6208 13636 6236
rect 12492 6196 12498 6208
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 16996 6239 17054 6245
rect 16996 6205 17008 6239
rect 17042 6236 17054 6239
rect 17512 6236 17540 6264
rect 17042 6208 17540 6236
rect 17042 6205 17054 6208
rect 16996 6199 17054 6205
rect 18414 6196 18420 6248
rect 18472 6245 18478 6248
rect 18472 6239 18510 6245
rect 18498 6236 18510 6239
rect 18874 6236 18880 6248
rect 18498 6208 18880 6236
rect 18498 6205 18510 6208
rect 18472 6199 18510 6205
rect 18472 6196 18478 6199
rect 18874 6196 18880 6208
rect 18932 6196 18938 6248
rect 22624 6239 22682 6245
rect 22624 6205 22636 6239
rect 22670 6236 22682 6239
rect 23124 6236 23152 6403
rect 23290 6400 23296 6412
rect 23348 6400 23354 6452
rect 24486 6440 24492 6452
rect 24447 6412 24492 6440
rect 24486 6400 24492 6412
rect 24544 6440 24550 6452
rect 24670 6440 24676 6452
rect 24544 6412 24676 6440
rect 24544 6400 24550 6412
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 24949 6375 25007 6381
rect 24949 6341 24961 6375
rect 24995 6372 25007 6375
rect 25222 6372 25228 6384
rect 24995 6344 25228 6372
rect 24995 6341 25007 6344
rect 24949 6335 25007 6341
rect 25222 6332 25228 6344
rect 25280 6332 25286 6384
rect 35434 6372 35440 6384
rect 35395 6344 35440 6372
rect 35434 6332 35440 6344
rect 35492 6332 35498 6384
rect 24854 6264 24860 6316
rect 24912 6304 24918 6316
rect 25133 6307 25191 6313
rect 25133 6304 25145 6307
rect 24912 6276 25145 6304
rect 24912 6264 24918 6276
rect 25133 6273 25145 6276
rect 25179 6273 25191 6307
rect 25406 6304 25412 6316
rect 25367 6276 25412 6304
rect 25133 6267 25191 6273
rect 25406 6264 25412 6276
rect 25464 6264 25470 6316
rect 22670 6208 23152 6236
rect 22670 6205 22682 6208
rect 22624 6199 22682 6205
rect 2314 6128 2320 6180
rect 2372 6168 2378 6180
rect 2863 6171 2921 6177
rect 2863 6168 2875 6171
rect 2372 6140 2875 6168
rect 2372 6128 2378 6140
rect 2863 6137 2875 6140
rect 2909 6168 2921 6171
rect 3789 6171 3847 6177
rect 3789 6168 3801 6171
rect 2909 6140 3801 6168
rect 2909 6137 2921 6140
rect 2863 6131 2921 6137
rect 3789 6137 3801 6140
rect 3835 6168 3847 6171
rect 4338 6168 4344 6180
rect 3835 6140 4344 6168
rect 3835 6137 3847 6140
rect 3789 6131 3847 6137
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 4433 6171 4491 6177
rect 4433 6137 4445 6171
rect 4479 6137 4491 6171
rect 4433 6131 4491 6137
rect 7009 6171 7067 6177
rect 7009 6137 7021 6171
rect 7055 6137 7067 6171
rect 9122 6168 9128 6180
rect 9083 6140 9128 6168
rect 7009 6131 7067 6137
rect 2038 6100 2044 6112
rect 1999 6072 2044 6100
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4448 6100 4476 6131
rect 6546 6100 6552 6112
rect 4120 6072 4476 6100
rect 6507 6072 6552 6100
rect 4120 6060 4126 6072
rect 6546 6060 6552 6072
rect 6604 6100 6610 6112
rect 7024 6100 7052 6131
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 9674 6128 9680 6180
rect 9732 6168 9738 6180
rect 10689 6171 10747 6177
rect 10689 6168 10701 6171
rect 9732 6140 10701 6168
rect 9732 6128 9738 6140
rect 10689 6137 10701 6140
rect 10735 6168 10747 6171
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 10735 6140 11529 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 11517 6137 11529 6140
rect 11563 6137 11575 6171
rect 13538 6168 13544 6180
rect 13451 6140 13544 6168
rect 11517 6131 11575 6137
rect 13538 6128 13544 6140
rect 13596 6168 13602 6180
rect 13995 6171 14053 6177
rect 13995 6168 14007 6171
rect 13596 6140 14007 6168
rect 13596 6128 13602 6140
rect 13995 6137 14007 6140
rect 14041 6168 14053 6171
rect 14642 6168 14648 6180
rect 14041 6140 14648 6168
rect 14041 6137 14053 6140
rect 13995 6131 14053 6137
rect 14642 6128 14648 6140
rect 14700 6128 14706 6180
rect 14826 6128 14832 6180
rect 14884 6168 14890 6180
rect 14921 6171 14979 6177
rect 14921 6168 14933 6171
rect 14884 6140 14933 6168
rect 14884 6128 14890 6140
rect 14921 6137 14933 6140
rect 14967 6168 14979 6171
rect 15565 6171 15623 6177
rect 15565 6168 15577 6171
rect 14967 6140 15577 6168
rect 14967 6137 14979 6140
rect 14921 6131 14979 6137
rect 15565 6137 15577 6140
rect 15611 6168 15623 6171
rect 15654 6168 15660 6180
rect 15611 6140 15660 6168
rect 15611 6137 15623 6140
rect 15565 6131 15623 6137
rect 15654 6128 15660 6140
rect 15712 6128 15718 6180
rect 19613 6171 19671 6177
rect 19613 6137 19625 6171
rect 19659 6137 19671 6171
rect 19613 6131 19671 6137
rect 12618 6100 12624 6112
rect 6604 6072 7052 6100
rect 12579 6072 12624 6100
rect 6604 6060 6610 6072
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 14553 6103 14611 6109
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 14734 6100 14740 6112
rect 14599 6072 14740 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 14734 6060 14740 6072
rect 14792 6060 14798 6112
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 16393 6103 16451 6109
rect 16393 6100 16405 6103
rect 15436 6072 16405 6100
rect 15436 6060 15442 6072
rect 16393 6069 16405 6072
rect 16439 6069 16451 6103
rect 16393 6063 16451 6069
rect 16574 6060 16580 6112
rect 16632 6100 16638 6112
rect 16761 6103 16819 6109
rect 16761 6100 16773 6103
rect 16632 6072 16773 6100
rect 16632 6060 16638 6072
rect 16761 6069 16773 6072
rect 16807 6069 16819 6103
rect 17862 6100 17868 6112
rect 17823 6072 17868 6100
rect 16761 6063 16819 6069
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 18966 6060 18972 6112
rect 19024 6100 19030 6112
rect 19245 6103 19303 6109
rect 19245 6100 19257 6103
rect 19024 6072 19257 6100
rect 19024 6060 19030 6072
rect 19245 6069 19257 6072
rect 19291 6100 19303 6103
rect 19628 6100 19656 6131
rect 19702 6128 19708 6180
rect 19760 6168 19766 6180
rect 20533 6171 20591 6177
rect 20533 6168 20545 6171
rect 19760 6140 20545 6168
rect 19760 6128 19766 6140
rect 20533 6137 20545 6140
rect 20579 6168 20591 6171
rect 21082 6168 21088 6180
rect 20579 6140 20944 6168
rect 21043 6140 21088 6168
rect 20579 6137 20591 6140
rect 20533 6131 20591 6137
rect 19291 6072 19656 6100
rect 19291 6069 19303 6072
rect 19245 6063 19303 6069
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 20809 6103 20867 6109
rect 20809 6100 20821 6103
rect 20772 6072 20821 6100
rect 20772 6060 20778 6072
rect 20809 6069 20821 6072
rect 20855 6069 20867 6103
rect 20916 6100 20944 6140
rect 21082 6128 21088 6140
rect 21140 6128 21146 6180
rect 21177 6171 21235 6177
rect 21177 6137 21189 6171
rect 21223 6137 21235 6171
rect 23474 6168 23480 6180
rect 23387 6140 23480 6168
rect 21177 6131 21235 6137
rect 21192 6100 21220 6131
rect 23474 6128 23480 6140
rect 23532 6168 23538 6180
rect 25222 6168 25228 6180
rect 23532 6140 25084 6168
rect 25183 6140 25228 6168
rect 23532 6128 23538 6140
rect 25056 6112 25084 6140
rect 25222 6128 25228 6140
rect 25280 6128 25286 6180
rect 22738 6109 22744 6112
rect 20916 6072 21220 6100
rect 22695 6103 22744 6109
rect 20809 6063 20867 6069
rect 22695 6069 22707 6103
rect 22741 6069 22744 6103
rect 22695 6063 22744 6069
rect 22738 6060 22744 6063
rect 22796 6060 22802 6112
rect 24026 6100 24032 6112
rect 23987 6072 24032 6100
rect 24026 6060 24032 6072
rect 24084 6060 24090 6112
rect 25038 6060 25044 6112
rect 25096 6060 25102 6112
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5865 6883 5899
rect 6825 5859 6883 5865
rect 9033 5899 9091 5905
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 9122 5896 9128 5908
rect 9079 5868 9128 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 2406 5788 2412 5840
rect 2464 5828 2470 5840
rect 2546 5831 2604 5837
rect 2546 5828 2558 5831
rect 2464 5800 2558 5828
rect 2464 5788 2470 5800
rect 2546 5797 2558 5800
rect 2592 5797 2604 5831
rect 3878 5828 3884 5840
rect 3839 5800 3884 5828
rect 2546 5791 2604 5797
rect 3878 5788 3884 5800
rect 3936 5788 3942 5840
rect 4338 5788 4344 5840
rect 4396 5837 4402 5840
rect 6270 5837 6276 5840
rect 4396 5831 4444 5837
rect 4396 5797 4398 5831
rect 4432 5797 4444 5831
rect 6267 5828 6276 5837
rect 6231 5800 6276 5828
rect 4396 5791 4444 5797
rect 6267 5791 6276 5800
rect 4396 5788 4402 5791
rect 6270 5788 6276 5791
rect 6328 5788 6334 5840
rect 6840 5828 6868 5859
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 10318 5896 10324 5908
rect 10279 5868 10324 5896
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 14001 5899 14059 5905
rect 14001 5865 14013 5899
rect 14047 5896 14059 5899
rect 14090 5896 14096 5908
rect 14047 5868 14096 5896
rect 14047 5865 14059 5868
rect 14001 5859 14059 5865
rect 14090 5856 14096 5868
rect 14148 5896 14154 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 14148 5868 14289 5896
rect 14148 5856 14154 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 18417 5899 18475 5905
rect 18417 5865 18429 5899
rect 18463 5896 18475 5899
rect 19153 5899 19211 5905
rect 19153 5896 19165 5899
rect 18463 5868 19165 5896
rect 18463 5865 18475 5868
rect 18417 5859 18475 5865
rect 19153 5865 19165 5868
rect 19199 5896 19211 5899
rect 19199 5868 19472 5896
rect 19199 5865 19211 5868
rect 19153 5859 19211 5865
rect 7466 5828 7472 5840
rect 6840 5800 7472 5828
rect 7466 5788 7472 5800
rect 7524 5828 7530 5840
rect 7837 5831 7895 5837
rect 7837 5828 7849 5831
rect 7524 5800 7849 5828
rect 7524 5788 7530 5800
rect 7837 5797 7849 5800
rect 7883 5797 7895 5831
rect 7837 5791 7895 5797
rect 10410 5788 10416 5840
rect 10468 5828 10474 5840
rect 10781 5831 10839 5837
rect 10781 5828 10793 5831
rect 10468 5800 10793 5828
rect 10468 5788 10474 5800
rect 10781 5797 10793 5800
rect 10827 5797 10839 5831
rect 10781 5791 10839 5797
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 12805 5831 12863 5837
rect 12805 5828 12817 5831
rect 12584 5800 12817 5828
rect 12584 5788 12590 5800
rect 12805 5797 12817 5800
rect 12851 5797 12863 5831
rect 12805 5791 12863 5797
rect 12894 5788 12900 5840
rect 12952 5828 12958 5840
rect 13443 5831 13501 5837
rect 13443 5828 13455 5831
rect 12952 5800 13455 5828
rect 12952 5788 12958 5800
rect 13443 5797 13455 5800
rect 13489 5828 13501 5831
rect 13538 5828 13544 5840
rect 13489 5800 13544 5828
rect 13489 5797 13501 5800
rect 13443 5791 13501 5797
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 14734 5788 14740 5840
rect 14792 5828 14798 5840
rect 15473 5831 15531 5837
rect 15473 5828 15485 5831
rect 14792 5800 15485 5828
rect 14792 5788 14798 5800
rect 15473 5797 15485 5800
rect 15519 5828 15531 5831
rect 16301 5831 16359 5837
rect 16301 5828 16313 5831
rect 15519 5800 16313 5828
rect 15519 5797 15531 5800
rect 15473 5791 15531 5797
rect 16301 5797 16313 5800
rect 16347 5797 16359 5831
rect 16301 5791 16359 5797
rect 17770 5788 17776 5840
rect 17828 5837 17834 5840
rect 17828 5831 17876 5837
rect 17828 5797 17830 5831
rect 17864 5797 17876 5831
rect 19334 5828 19340 5840
rect 19295 5800 19340 5828
rect 17828 5791 17876 5797
rect 17828 5788 17834 5791
rect 19334 5788 19340 5800
rect 19392 5788 19398 5840
rect 19444 5837 19472 5868
rect 19429 5831 19487 5837
rect 19429 5797 19441 5831
rect 19475 5828 19487 5831
rect 19702 5828 19708 5840
rect 19475 5800 19708 5828
rect 19475 5797 19487 5800
rect 19429 5791 19487 5797
rect 19702 5788 19708 5800
rect 19760 5788 19766 5840
rect 21266 5837 21272 5840
rect 21263 5828 21272 5837
rect 21227 5800 21272 5828
rect 21263 5791 21272 5800
rect 21266 5788 21272 5791
rect 21324 5788 21330 5840
rect 22557 5831 22615 5837
rect 22557 5797 22569 5831
rect 22603 5828 22615 5831
rect 22738 5828 22744 5840
rect 22603 5800 22744 5828
rect 22603 5797 22615 5800
rect 22557 5791 22615 5797
rect 22738 5788 22744 5800
rect 22796 5788 22802 5840
rect 22830 5788 22836 5840
rect 22888 5828 22894 5840
rect 24578 5828 24584 5840
rect 22888 5800 22933 5828
rect 24539 5800 24584 5828
rect 22888 5788 22894 5800
rect 24578 5788 24584 5800
rect 24636 5788 24642 5840
rect 3145 5763 3203 5769
rect 3145 5729 3157 5763
rect 3191 5760 3203 5763
rect 4246 5760 4252 5772
rect 3191 5732 4252 5760
rect 3191 5729 3203 5732
rect 3145 5723 3203 5729
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 11333 5763 11391 5769
rect 11333 5729 11345 5763
rect 11379 5760 11391 5763
rect 11379 5732 15240 5760
rect 11379 5729 11391 5732
rect 11333 5723 11391 5729
rect 2222 5692 2228 5704
rect 2183 5664 2228 5692
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 4062 5692 4068 5704
rect 4023 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 6638 5692 6644 5704
rect 5951 5664 6644 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7745 5695 7803 5701
rect 7745 5692 7757 5695
rect 7432 5664 7757 5692
rect 7432 5652 7438 5664
rect 7745 5661 7757 5664
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 1765 5627 1823 5633
rect 1765 5593 1777 5627
rect 1811 5624 1823 5627
rect 2590 5624 2596 5636
rect 1811 5596 2596 5624
rect 1811 5593 1823 5596
rect 1765 5587 1823 5593
rect 2590 5584 2596 5596
rect 2648 5584 2654 5636
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 3878 5624 3884 5636
rect 2740 5596 3884 5624
rect 2740 5584 2746 5596
rect 3878 5584 3884 5596
rect 3936 5584 3942 5636
rect 7190 5584 7196 5636
rect 7248 5624 7254 5636
rect 8036 5624 8064 5655
rect 10502 5652 10508 5704
rect 10560 5692 10566 5704
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10560 5664 10701 5692
rect 10560 5652 10566 5664
rect 10689 5661 10701 5664
rect 10735 5692 10747 5695
rect 11054 5692 11060 5704
rect 10735 5664 11060 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13538 5692 13544 5704
rect 13127 5664 13544 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 13538 5652 13544 5664
rect 13596 5692 13602 5704
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 13596 5664 14657 5692
rect 13596 5652 13602 5664
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 15212 5692 15240 5732
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 18693 5763 18751 5769
rect 18693 5760 18705 5763
rect 17092 5732 18705 5760
rect 17092 5720 17098 5732
rect 18693 5729 18705 5732
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 25222 5720 25228 5772
rect 25280 5760 25286 5772
rect 26605 5763 26663 5769
rect 26605 5760 26617 5763
rect 25280 5732 26617 5760
rect 25280 5720 25286 5732
rect 26605 5729 26617 5732
rect 26651 5760 26663 5763
rect 27246 5760 27252 5772
rect 26651 5732 27252 5760
rect 26651 5729 26663 5732
rect 26605 5723 26663 5729
rect 27246 5720 27252 5732
rect 27304 5720 27310 5772
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 15212 5664 15393 5692
rect 14645 5655 14703 5661
rect 15381 5661 15393 5664
rect 15427 5692 15439 5695
rect 15562 5692 15568 5704
rect 15427 5664 15568 5692
rect 15427 5661 15439 5664
rect 15381 5655 15439 5661
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 15746 5652 15752 5664
rect 15804 5692 15810 5704
rect 16666 5692 16672 5704
rect 15804 5664 16672 5692
rect 15804 5652 15810 5664
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 20901 5695 20959 5701
rect 20901 5661 20913 5695
rect 20947 5692 20959 5695
rect 21358 5692 21364 5704
rect 20947 5664 21364 5692
rect 20947 5661 20959 5664
rect 20901 5655 20959 5661
rect 7248 5596 8064 5624
rect 12529 5627 12587 5633
rect 7248 5584 7254 5596
rect 12529 5593 12541 5627
rect 12575 5624 12587 5627
rect 12618 5624 12624 5636
rect 12575 5596 12624 5624
rect 12575 5593 12587 5596
rect 12529 5587 12587 5593
rect 12618 5584 12624 5596
rect 12676 5624 12682 5636
rect 13262 5624 13268 5636
rect 12676 5596 13268 5624
rect 12676 5584 12682 5596
rect 13262 5584 13268 5596
rect 13320 5584 13326 5636
rect 2130 5556 2136 5568
rect 2091 5528 2136 5556
rect 2130 5516 2136 5528
rect 2188 5516 2194 5568
rect 3513 5559 3571 5565
rect 3513 5525 3525 5559
rect 3559 5556 3571 5559
rect 3602 5556 3608 5568
rect 3559 5528 3608 5556
rect 3559 5525 3571 5528
rect 3513 5519 3571 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 4982 5556 4988 5568
rect 4943 5528 4988 5556
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 7561 5559 7619 5565
rect 7561 5525 7573 5559
rect 7607 5556 7619 5559
rect 8202 5556 8208 5568
rect 7607 5528 8208 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 14918 5516 14924 5568
rect 14976 5556 14982 5568
rect 15013 5559 15071 5565
rect 15013 5556 15025 5559
rect 14976 5528 15025 5556
rect 14976 5516 14982 5528
rect 15013 5525 15025 5528
rect 15059 5525 15071 5559
rect 15013 5519 15071 5525
rect 16761 5559 16819 5565
rect 16761 5525 16773 5559
rect 16807 5556 16819 5559
rect 16850 5556 16856 5568
rect 16807 5528 16856 5556
rect 16807 5525 16819 5528
rect 16761 5519 16819 5525
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 17512 5556 17540 5655
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 23017 5695 23075 5701
rect 23017 5661 23029 5695
rect 23063 5661 23075 5695
rect 23017 5655 23075 5661
rect 19886 5624 19892 5636
rect 19799 5596 19892 5624
rect 19886 5584 19892 5596
rect 19944 5624 19950 5636
rect 20622 5624 20628 5636
rect 19944 5596 20628 5624
rect 19944 5584 19950 5596
rect 20622 5584 20628 5596
rect 20680 5624 20686 5636
rect 23032 5624 23060 5655
rect 24026 5652 24032 5704
rect 24084 5692 24090 5704
rect 24486 5692 24492 5704
rect 24084 5664 24492 5692
rect 24084 5652 24090 5664
rect 24486 5652 24492 5664
rect 24544 5652 24550 5704
rect 26142 5652 26148 5704
rect 26200 5692 26206 5704
rect 26513 5695 26571 5701
rect 26513 5692 26525 5695
rect 26200 5664 26525 5692
rect 26200 5652 26206 5664
rect 26513 5661 26525 5664
rect 26559 5661 26571 5695
rect 26513 5655 26571 5661
rect 27617 5695 27675 5701
rect 27617 5661 27629 5695
rect 27663 5692 27675 5695
rect 27982 5692 27988 5704
rect 27663 5664 27988 5692
rect 27663 5661 27675 5664
rect 27617 5655 27675 5661
rect 27982 5652 27988 5664
rect 28040 5652 28046 5704
rect 25038 5624 25044 5636
rect 20680 5596 23060 5624
rect 24999 5596 25044 5624
rect 20680 5584 20686 5596
rect 25038 5584 25044 5596
rect 25096 5584 25102 5636
rect 17862 5556 17868 5568
rect 17451 5528 17868 5556
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 20346 5556 20352 5568
rect 20307 5528 20352 5556
rect 20346 5516 20352 5528
rect 20404 5516 20410 5568
rect 21818 5556 21824 5568
rect 21779 5528 21824 5556
rect 21818 5516 21824 5528
rect 21876 5516 21882 5568
rect 22094 5516 22100 5568
rect 22152 5556 22158 5568
rect 22152 5528 22197 5556
rect 22152 5516 22158 5528
rect 23382 5516 23388 5568
rect 23440 5556 23446 5568
rect 23661 5559 23719 5565
rect 23661 5556 23673 5559
rect 23440 5528 23673 5556
rect 23440 5516 23446 5528
rect 23661 5525 23673 5528
rect 23707 5525 23719 5559
rect 23661 5519 23719 5525
rect 24946 5516 24952 5568
rect 25004 5556 25010 5568
rect 25406 5556 25412 5568
rect 25004 5528 25412 5556
rect 25004 5516 25010 5528
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 27614 5516 27620 5568
rect 27672 5556 27678 5568
rect 27893 5559 27951 5565
rect 27893 5556 27905 5559
rect 27672 5528 27905 5556
rect 27672 5516 27678 5528
rect 27893 5525 27905 5528
rect 27939 5525 27951 5559
rect 27893 5519 27951 5525
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1452 5324 1593 5352
rect 1452 5312 1458 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 2406 5352 2412 5364
rect 2367 5324 2412 5352
rect 1581 5315 1639 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 6546 5352 6552 5364
rect 5951 5324 6552 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 7374 5352 7380 5364
rect 6840 5324 7380 5352
rect 2038 5216 2044 5228
rect 1412 5188 2044 5216
rect 1412 5157 1440 5188
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 2590 5176 2596 5228
rect 2648 5216 2654 5228
rect 6840 5225 6868 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 9122 5352 9128 5364
rect 8803 5324 9128 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 10468 5324 10517 5352
rect 10468 5312 10474 5324
rect 10505 5321 10517 5324
rect 10551 5352 10563 5355
rect 10781 5355 10839 5361
rect 10781 5352 10793 5355
rect 10551 5324 10793 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 10781 5321 10793 5324
rect 10827 5321 10839 5355
rect 10781 5315 10839 5321
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11149 5355 11207 5361
rect 11149 5352 11161 5355
rect 11112 5324 11161 5352
rect 11112 5312 11118 5324
rect 11149 5321 11161 5324
rect 11195 5321 11207 5355
rect 11149 5315 11207 5321
rect 11517 5355 11575 5361
rect 11517 5321 11529 5355
rect 11563 5352 11575 5355
rect 11609 5355 11667 5361
rect 11609 5352 11621 5355
rect 11563 5324 11621 5352
rect 11563 5321 11575 5324
rect 11517 5315 11575 5321
rect 11609 5321 11621 5324
rect 11655 5321 11667 5355
rect 11609 5315 11667 5321
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12894 5352 12900 5364
rect 12299 5324 12900 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 9493 5287 9551 5293
rect 9493 5253 9505 5287
rect 9539 5284 9551 5287
rect 12268 5284 12296 5315
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 15654 5352 15660 5364
rect 15615 5324 15660 5352
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 16025 5355 16083 5361
rect 16025 5352 16037 5355
rect 15804 5324 16037 5352
rect 15804 5312 15810 5324
rect 16025 5321 16037 5324
rect 16071 5352 16083 5355
rect 17034 5352 17040 5364
rect 16071 5324 17040 5352
rect 16071 5321 16083 5324
rect 16025 5315 16083 5321
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 18966 5352 18972 5364
rect 18927 5324 18972 5352
rect 18966 5312 18972 5324
rect 19024 5312 19030 5364
rect 20714 5352 20720 5364
rect 20627 5324 20720 5352
rect 20714 5312 20720 5324
rect 20772 5352 20778 5364
rect 22830 5352 22836 5364
rect 20772 5324 22836 5352
rect 20772 5312 20778 5324
rect 22830 5312 22836 5324
rect 22888 5352 22894 5364
rect 22925 5355 22983 5361
rect 22925 5352 22937 5355
rect 22888 5324 22937 5352
rect 22888 5312 22894 5324
rect 22925 5321 22937 5324
rect 22971 5321 22983 5355
rect 24210 5352 24216 5364
rect 24171 5324 24216 5352
rect 22925 5315 22983 5321
rect 24210 5312 24216 5324
rect 24268 5312 24274 5364
rect 24578 5352 24584 5364
rect 24539 5324 24584 5352
rect 24578 5312 24584 5324
rect 24636 5312 24642 5364
rect 27246 5352 27252 5364
rect 27207 5324 27252 5352
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 35066 5312 35072 5364
rect 35124 5352 35130 5364
rect 35621 5355 35679 5361
rect 35621 5352 35633 5355
rect 35124 5324 35633 5352
rect 35124 5312 35130 5324
rect 35621 5321 35633 5324
rect 35667 5321 35679 5355
rect 35621 5315 35679 5321
rect 9539 5256 12296 5284
rect 9539 5253 9551 5256
rect 9493 5247 9551 5253
rect 6825 5219 6883 5225
rect 2648 5188 3556 5216
rect 2648 5176 2654 5188
rect 3528 5160 3556 5188
rect 6825 5185 6837 5219
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5216 7895 5219
rect 8202 5216 8208 5228
rect 7883 5188 8208 5216
rect 7883 5185 7895 5188
rect 7837 5179 7895 5185
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 2130 5108 2136 5160
rect 2188 5148 2194 5160
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 2188 5120 2513 5148
rect 2188 5108 2194 5120
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5117 3295 5151
rect 3510 5148 3516 5160
rect 3471 5120 3516 5148
rect 3237 5111 3295 5117
rect 3252 5080 3280 5111
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 3786 5148 3792 5160
rect 3747 5120 3792 5148
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 5074 5148 5080 5160
rect 5031 5120 5080 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 9125 5151 9183 5157
rect 9125 5117 9137 5151
rect 9171 5148 9183 5151
rect 9582 5148 9588 5160
rect 9171 5120 9588 5148
rect 9171 5117 9183 5120
rect 9125 5111 9183 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 3602 5080 3608 5092
rect 3252 5052 3608 5080
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 4338 5080 4344 5092
rect 4251 5052 4344 5080
rect 4338 5040 4344 5052
rect 4396 5080 4402 5092
rect 4893 5083 4951 5089
rect 4893 5080 4905 5083
rect 4396 5052 4905 5080
rect 4396 5040 4402 5052
rect 4893 5049 4905 5052
rect 4939 5080 4951 5083
rect 5347 5083 5405 5089
rect 5347 5080 5359 5083
rect 4939 5052 5359 5080
rect 4939 5049 4951 5052
rect 4893 5043 4951 5049
rect 5347 5049 5359 5052
rect 5393 5080 5405 5083
rect 6270 5080 6276 5092
rect 5393 5052 6276 5080
rect 5393 5049 5405 5052
rect 5347 5043 5405 5049
rect 6270 5040 6276 5052
rect 6328 5080 6334 5092
rect 8202 5089 8208 5092
rect 7745 5083 7803 5089
rect 7745 5080 7757 5083
rect 6328 5052 7757 5080
rect 6328 5040 6334 5052
rect 7745 5049 7757 5052
rect 7791 5080 7803 5083
rect 8199 5080 8208 5089
rect 7791 5052 8208 5080
rect 7791 5049 7803 5052
rect 7745 5043 7803 5049
rect 8199 5043 8208 5052
rect 8260 5080 8266 5092
rect 9968 5089 9996 5256
rect 21542 5244 21548 5296
rect 21600 5244 21606 5296
rect 23799 5287 23857 5293
rect 23799 5253 23811 5287
rect 23845 5284 23857 5287
rect 24762 5284 24768 5296
rect 23845 5256 24768 5284
rect 23845 5253 23857 5256
rect 23799 5247 23857 5253
rect 24762 5244 24768 5256
rect 24820 5244 24826 5296
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 11609 5219 11667 5225
rect 11609 5216 11621 5219
rect 10192 5188 11621 5216
rect 10192 5176 10198 5188
rect 11609 5185 11621 5188
rect 11655 5216 11667 5219
rect 21560 5216 21588 5244
rect 21637 5219 21695 5225
rect 21637 5216 21649 5219
rect 11655 5188 13124 5216
rect 21560 5188 21649 5216
rect 11655 5185 11667 5188
rect 11609 5179 11667 5185
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 12526 5148 12532 5160
rect 11379 5120 11836 5148
rect 12487 5120 12532 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 9947 5083 10005 5089
rect 9947 5080 9959 5083
rect 8260 5052 9959 5080
rect 8202 5040 8208 5043
rect 8260 5040 8266 5052
rect 9947 5049 9959 5052
rect 9993 5049 10005 5083
rect 9947 5043 10005 5049
rect 11808 5024 11836 5120
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 13096 5157 13124 5188
rect 21637 5185 21649 5188
rect 21683 5185 21695 5219
rect 22278 5216 22284 5228
rect 22191 5188 22284 5216
rect 21637 5179 21695 5185
rect 22278 5176 22284 5188
rect 22336 5216 22342 5228
rect 23382 5216 23388 5228
rect 22336 5188 23388 5216
rect 22336 5176 22342 5188
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 25038 5216 25044 5228
rect 24999 5188 25044 5216
rect 25038 5176 25044 5188
rect 25096 5176 25102 5228
rect 27522 5216 27528 5228
rect 27483 5188 27528 5216
rect 27522 5176 27528 5188
rect 27580 5176 27586 5228
rect 13081 5151 13139 5157
rect 13081 5117 13093 5151
rect 13127 5117 13139 5151
rect 13262 5148 13268 5160
rect 13223 5120 13268 5148
rect 13081 5111 13139 5117
rect 13096 5080 13124 5111
rect 13262 5108 13268 5120
rect 13320 5108 13326 5160
rect 13722 5148 13728 5160
rect 13683 5120 13728 5148
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 13906 5108 13912 5160
rect 13964 5148 13970 5160
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 13964 5120 14749 5148
rect 13964 5108 13970 5120
rect 14737 5117 14749 5120
rect 14783 5148 14795 5151
rect 14918 5148 14924 5160
rect 14783 5120 14924 5148
rect 14783 5117 14795 5120
rect 14737 5111 14795 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 16574 5108 16580 5160
rect 16632 5148 16638 5160
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 16632 5120 16681 5148
rect 16632 5108 16638 5120
rect 16669 5117 16681 5120
rect 16715 5148 16727 5151
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 16715 5120 17325 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 17954 5108 17960 5160
rect 18012 5148 18018 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 18012 5120 18061 5148
rect 18012 5108 18018 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 19794 5148 19800 5160
rect 19755 5120 19800 5148
rect 18049 5111 18107 5117
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 23728 5151 23786 5157
rect 23728 5117 23740 5151
rect 23774 5148 23786 5151
rect 24210 5148 24216 5160
rect 23774 5120 24216 5148
rect 23774 5117 23786 5120
rect 23728 5111 23786 5117
rect 24210 5108 24216 5120
rect 24268 5108 24274 5160
rect 26326 5108 26332 5160
rect 26384 5148 26390 5160
rect 26456 5151 26514 5157
rect 26456 5148 26468 5151
rect 26384 5120 26468 5148
rect 26384 5108 26390 5120
rect 26456 5117 26468 5120
rect 26502 5148 26514 5151
rect 26878 5148 26884 5160
rect 26502 5120 26884 5148
rect 26502 5117 26514 5120
rect 26456 5111 26514 5117
rect 26878 5108 26884 5120
rect 26936 5108 26942 5160
rect 28994 5108 29000 5160
rect 29052 5148 29058 5160
rect 35437 5151 35495 5157
rect 35437 5148 35449 5151
rect 29052 5120 35449 5148
rect 29052 5108 29058 5120
rect 35437 5117 35449 5120
rect 35483 5148 35495 5151
rect 35989 5151 36047 5157
rect 35989 5148 36001 5151
rect 35483 5120 36001 5148
rect 35483 5117 35495 5120
rect 35437 5111 35495 5117
rect 35989 5117 36001 5120
rect 36035 5117 36047 5151
rect 35989 5111 36047 5117
rect 14185 5083 14243 5089
rect 14185 5080 14197 5083
rect 13096 5052 14197 5080
rect 14185 5049 14197 5052
rect 14231 5049 14243 5083
rect 14642 5080 14648 5092
rect 14555 5052 14648 5080
rect 14185 5043 14243 5049
rect 14642 5040 14648 5052
rect 14700 5080 14706 5092
rect 15102 5089 15108 5092
rect 15099 5080 15108 5089
rect 14700 5052 15108 5080
rect 14700 5040 14706 5052
rect 15099 5043 15108 5052
rect 15102 5040 15108 5043
rect 15160 5040 15166 5092
rect 15286 5040 15292 5092
rect 15344 5080 15350 5092
rect 16393 5083 16451 5089
rect 16393 5080 16405 5083
rect 15344 5052 16405 5080
rect 15344 5040 15350 5052
rect 16393 5049 16405 5052
rect 16439 5080 16451 5083
rect 16485 5083 16543 5089
rect 16485 5080 16497 5083
rect 16439 5052 16497 5080
rect 16439 5049 16451 5052
rect 16393 5043 16451 5049
rect 16485 5049 16497 5052
rect 16531 5049 16543 5083
rect 17034 5080 17040 5092
rect 16995 5052 17040 5080
rect 16485 5043 16543 5049
rect 17034 5040 17040 5052
rect 17092 5040 17098 5092
rect 17770 5040 17776 5092
rect 17828 5080 17834 5092
rect 17865 5083 17923 5089
rect 17865 5080 17877 5083
rect 17828 5052 17877 5080
rect 17828 5040 17834 5052
rect 17865 5049 17877 5052
rect 17911 5080 17923 5083
rect 18138 5080 18144 5092
rect 17911 5052 18144 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18138 5040 18144 5052
rect 18196 5080 18202 5092
rect 18411 5083 18469 5089
rect 18411 5080 18423 5083
rect 18196 5052 18423 5080
rect 18196 5040 18202 5052
rect 18411 5049 18423 5052
rect 18457 5080 18469 5083
rect 19705 5083 19763 5089
rect 19705 5080 19717 5083
rect 18457 5052 19717 5080
rect 18457 5049 18469 5052
rect 18411 5043 18469 5049
rect 19705 5049 19717 5052
rect 19751 5080 19763 5083
rect 20159 5083 20217 5089
rect 20159 5080 20171 5083
rect 19751 5052 20171 5080
rect 19751 5049 19763 5052
rect 19705 5043 19763 5049
rect 20159 5049 20171 5052
rect 20205 5080 20217 5083
rect 21266 5080 21272 5092
rect 20205 5052 21272 5080
rect 20205 5049 20217 5052
rect 20159 5043 20217 5049
rect 20916 5024 20944 5052
rect 21266 5040 21272 5052
rect 21324 5040 21330 5092
rect 21726 5040 21732 5092
rect 21784 5080 21790 5092
rect 22002 5080 22008 5092
rect 21784 5052 22008 5080
rect 21784 5040 21790 5052
rect 22002 5040 22008 5052
rect 22060 5040 22066 5092
rect 24762 5080 24768 5092
rect 24723 5052 24768 5080
rect 24762 5040 24768 5052
rect 24820 5040 24826 5092
rect 24857 5083 24915 5089
rect 24857 5049 24869 5083
rect 24903 5080 24915 5083
rect 25685 5083 25743 5089
rect 25685 5080 25697 5083
rect 24903 5052 25697 5080
rect 24903 5049 24915 5052
rect 24857 5043 24915 5049
rect 25685 5049 25697 5052
rect 25731 5049 25743 5083
rect 25685 5043 25743 5049
rect 27617 5083 27675 5089
rect 27617 5049 27629 5083
rect 27663 5080 27675 5083
rect 27982 5080 27988 5092
rect 27663 5052 27988 5080
rect 27663 5049 27675 5052
rect 27617 5043 27675 5049
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 6638 5012 6644 5024
rect 2832 4984 2877 5012
rect 6599 4984 6644 5012
rect 2832 4972 2838 4984
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 11790 5012 11796 5024
rect 11751 4984 11796 5012
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 13630 5012 13636 5024
rect 13591 4984 13636 5012
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 19334 5012 19340 5024
rect 19295 4984 19340 5012
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20956 4984 21005 5012
rect 20956 4972 20962 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 21358 5012 21364 5024
rect 21319 4984 21364 5012
rect 20993 4975 21051 4981
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 22649 5015 22707 5021
rect 22649 4981 22661 5015
rect 22695 5012 22707 5015
rect 23290 5012 23296 5024
rect 22695 4984 23296 5012
rect 22695 4981 22707 4984
rect 22649 4975 22707 4981
rect 23290 4972 23296 4984
rect 23348 4972 23354 5024
rect 23474 5012 23480 5024
rect 23435 4984 23480 5012
rect 23474 4972 23480 4984
rect 23532 4972 23538 5024
rect 24670 4972 24676 5024
rect 24728 5012 24734 5024
rect 24872 5012 24900 5043
rect 27982 5040 27988 5052
rect 28040 5040 28046 5092
rect 28169 5083 28227 5089
rect 28169 5049 28181 5083
rect 28215 5080 28227 5083
rect 28258 5080 28264 5092
rect 28215 5052 28264 5080
rect 28215 5049 28227 5052
rect 28169 5043 28227 5049
rect 28258 5040 28264 5052
rect 28316 5040 28322 5092
rect 24728 4984 24900 5012
rect 26559 5015 26617 5021
rect 24728 4972 24734 4984
rect 26559 4981 26571 5015
rect 26605 5012 26617 5015
rect 26786 5012 26792 5024
rect 26605 4984 26792 5012
rect 26605 4981 26617 4984
rect 26559 4975 26617 4981
rect 26786 4972 26792 4984
rect 26844 4972 26850 5024
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2222 4808 2228 4820
rect 1995 4780 2228 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2222 4768 2228 4780
rect 2280 4808 2286 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 2280 4780 3801 4808
rect 2280 4768 2286 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4203 4811 4261 4817
rect 4203 4808 4215 4811
rect 4028 4780 4215 4808
rect 4028 4768 4034 4780
rect 4203 4777 4215 4780
rect 4249 4777 4261 4811
rect 5074 4808 5080 4820
rect 4987 4780 5080 4808
rect 4203 4771 4261 4777
rect 5074 4768 5080 4780
rect 5132 4808 5138 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5132 4780 5273 4808
rect 5132 4768 5138 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 7653 4811 7711 4817
rect 7653 4808 7665 4811
rect 7524 4780 7665 4808
rect 7524 4768 7530 4780
rect 7653 4777 7665 4780
rect 7699 4777 7711 4811
rect 7653 4771 7711 4777
rect 8757 4811 8815 4817
rect 8757 4777 8769 4811
rect 8803 4808 8815 4811
rect 9490 4808 9496 4820
rect 8803 4780 9496 4808
rect 8803 4777 8815 4780
rect 8757 4771 8815 4777
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 9640 4780 9781 4808
rect 9640 4768 9646 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9769 4771 9827 4777
rect 15105 4811 15163 4817
rect 15105 4777 15117 4811
rect 15151 4808 15163 4811
rect 15746 4808 15752 4820
rect 15151 4780 15752 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 18049 4811 18107 4817
rect 18049 4777 18061 4811
rect 18095 4808 18107 4811
rect 18138 4808 18144 4820
rect 18095 4780 18144 4808
rect 18095 4777 18107 4780
rect 18049 4771 18107 4777
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 21266 4808 21272 4820
rect 20763 4780 21272 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 21266 4768 21272 4780
rect 21324 4808 21330 4820
rect 21818 4808 21824 4820
rect 21324 4780 21824 4808
rect 21324 4768 21330 4780
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 23474 4808 23480 4820
rect 23435 4780 23480 4808
rect 23474 4768 23480 4780
rect 23532 4768 23538 4820
rect 24486 4808 24492 4820
rect 24447 4780 24492 4808
rect 24486 4768 24492 4780
rect 24544 4768 24550 4820
rect 25222 4768 25228 4820
rect 25280 4808 25286 4820
rect 25501 4811 25559 4817
rect 25501 4808 25513 4811
rect 25280 4780 25513 4808
rect 25280 4768 25286 4780
rect 25501 4777 25513 4780
rect 25547 4777 25559 4811
rect 25501 4771 25559 4777
rect 26651 4811 26709 4817
rect 26651 4777 26663 4811
rect 26697 4808 26709 4811
rect 27522 4808 27528 4820
rect 26697 4780 27528 4808
rect 26697 4777 26709 4780
rect 26651 4771 26709 4777
rect 27522 4768 27528 4780
rect 27580 4768 27586 4820
rect 2130 4700 2136 4752
rect 2188 4740 2194 4752
rect 8202 4749 8208 4752
rect 8199 4740 8208 4749
rect 2188 4712 5212 4740
rect 8163 4712 8208 4740
rect 2188 4700 2194 4712
rect 5184 4684 5212 4712
rect 8199 4703 8208 4712
rect 8202 4700 8208 4703
rect 8260 4700 8266 4752
rect 12161 4743 12219 4749
rect 12161 4740 12173 4743
rect 10888 4712 12173 4740
rect 10888 4684 10916 4712
rect 12161 4709 12173 4712
rect 12207 4740 12219 4743
rect 12253 4743 12311 4749
rect 12253 4740 12265 4743
rect 12207 4712 12265 4740
rect 12207 4709 12219 4712
rect 12161 4703 12219 4709
rect 12253 4709 12265 4712
rect 12299 4709 12311 4743
rect 13906 4740 13912 4752
rect 13867 4712 13912 4740
rect 12253 4703 12311 4709
rect 13906 4700 13912 4712
rect 13964 4700 13970 4752
rect 16022 4700 16028 4752
rect 16080 4740 16086 4752
rect 16080 4712 17080 4740
rect 16080 4700 16086 4712
rect 1762 4672 1768 4684
rect 1723 4644 1768 4672
rect 1762 4632 1768 4644
rect 1820 4632 1826 4684
rect 2409 4675 2467 4681
rect 2409 4641 2421 4675
rect 2455 4641 2467 4675
rect 2682 4672 2688 4684
rect 2643 4644 2688 4672
rect 2409 4635 2467 4641
rect 2424 4604 2452 4635
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4672 3111 4675
rect 3099 4644 3556 4672
rect 3099 4641 3111 4644
rect 3053 4635 3111 4641
rect 2958 4604 2964 4616
rect 2424 4576 2964 4604
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 3528 4477 3556 4644
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 4132 4675 4190 4681
rect 4132 4672 4144 4675
rect 3752 4644 4144 4672
rect 3752 4632 3758 4644
rect 4132 4641 4144 4644
rect 4178 4672 4190 4675
rect 4246 4672 4252 4684
rect 4178 4644 4252 4672
rect 4178 4641 4190 4644
rect 4132 4635 4190 4641
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 5166 4672 5172 4684
rect 5079 4644 5172 4672
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5902 4672 5908 4684
rect 5863 4644 5908 4672
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4641 6239 4675
rect 6546 4672 6552 4684
rect 6507 4644 6552 4672
rect 6181 4635 6239 4641
rect 6196 4604 6224 4635
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4641 10011 4675
rect 10134 4672 10140 4684
rect 10095 4644 10140 4672
rect 9953 4635 10011 4641
rect 6454 4604 6460 4616
rect 6196 4576 6460 4604
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 8018 4604 8024 4616
rect 7883 4576 8024 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 9968 4604 9996 4635
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10226 4632 10232 4684
rect 10284 4672 10290 4684
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 10284 4644 10517 4672
rect 10284 4632 10290 4644
rect 10505 4641 10517 4644
rect 10551 4641 10563 4675
rect 10870 4672 10876 4684
rect 10831 4644 10876 4672
rect 10505 4635 10563 4641
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 11940 4644 12449 4672
rect 11940 4632 11946 4644
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 13078 4672 13084 4684
rect 13039 4644 13084 4672
rect 12437 4635 12495 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13170 4632 13176 4684
rect 13228 4672 13234 4684
rect 13265 4675 13323 4681
rect 13265 4672 13277 4675
rect 13228 4644 13277 4672
rect 13228 4632 13234 4644
rect 13265 4641 13277 4644
rect 13311 4641 13323 4675
rect 13630 4672 13636 4684
rect 13591 4644 13636 4672
rect 13265 4635 13323 4641
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 15470 4632 15476 4684
rect 15528 4672 15534 4684
rect 17052 4681 17080 4712
rect 17126 4700 17132 4752
rect 17184 4740 17190 4752
rect 17678 4740 17684 4752
rect 17184 4712 17448 4740
rect 17639 4712 17684 4740
rect 17184 4700 17190 4712
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 15528 4644 16221 4672
rect 15528 4632 15534 4644
rect 16209 4641 16221 4644
rect 16255 4641 16267 4675
rect 16209 4635 16267 4641
rect 16945 4675 17003 4681
rect 16945 4641 16957 4675
rect 16991 4641 17003 4675
rect 16945 4635 17003 4641
rect 17037 4675 17095 4681
rect 17037 4641 17049 4675
rect 17083 4672 17095 4675
rect 17310 4672 17316 4684
rect 17083 4644 17316 4672
rect 17083 4641 17095 4644
rect 17037 4635 17095 4641
rect 10594 4604 10600 4616
rect 9968 4576 10600 4604
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4604 12219 4607
rect 13648 4604 13676 4632
rect 12207 4576 13676 4604
rect 14277 4607 14335 4613
rect 12207 4573 12219 4576
rect 12161 4567 12219 4573
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 14323 4576 15761 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 15749 4573 15761 4576
rect 15795 4604 15807 4607
rect 16758 4604 16764 4616
rect 15795 4576 16764 4604
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 16758 4564 16764 4576
rect 16816 4604 16822 4616
rect 16960 4604 16988 4635
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17420 4681 17448 4712
rect 17678 4700 17684 4712
rect 17736 4700 17742 4752
rect 19794 4700 19800 4752
rect 19852 4740 19858 4752
rect 19981 4743 20039 4749
rect 19981 4740 19993 4743
rect 19852 4712 19993 4740
rect 19852 4700 19858 4712
rect 19981 4709 19993 4712
rect 20027 4740 20039 4743
rect 20257 4743 20315 4749
rect 20257 4740 20269 4743
rect 20027 4712 20269 4740
rect 20027 4709 20039 4712
rect 19981 4703 20039 4709
rect 20257 4709 20269 4712
rect 20303 4709 20315 4743
rect 20257 4703 20315 4709
rect 20806 4700 20812 4752
rect 20864 4740 20870 4752
rect 21039 4743 21097 4749
rect 21039 4740 21051 4743
rect 20864 4712 21051 4740
rect 20864 4700 20870 4712
rect 21039 4709 21051 4712
rect 21085 4709 21097 4743
rect 21358 4740 21364 4752
rect 21319 4712 21364 4740
rect 21039 4703 21097 4709
rect 21358 4700 21364 4712
rect 21416 4700 21422 4752
rect 24854 4700 24860 4752
rect 24912 4749 24918 4752
rect 24912 4743 24960 4749
rect 24912 4709 24914 4743
rect 24948 4709 24960 4743
rect 24912 4703 24960 4709
rect 24912 4700 24918 4703
rect 26786 4700 26792 4752
rect 26844 4740 26850 4752
rect 27614 4740 27620 4752
rect 26844 4712 27620 4740
rect 26844 4700 26850 4712
rect 27614 4700 27620 4712
rect 27672 4700 27678 4752
rect 27706 4700 27712 4752
rect 27764 4740 27770 4752
rect 28258 4740 28264 4752
rect 27764 4712 27809 4740
rect 28219 4712 28264 4740
rect 27764 4700 27770 4712
rect 28258 4700 28264 4712
rect 28316 4700 28322 4752
rect 17405 4675 17463 4681
rect 17405 4641 17417 4675
rect 17451 4641 17463 4675
rect 18506 4672 18512 4684
rect 18467 4644 18512 4672
rect 17405 4635 17463 4641
rect 18506 4632 18512 4644
rect 18564 4632 18570 4684
rect 18782 4632 18788 4684
rect 18840 4672 18846 4684
rect 18969 4675 19027 4681
rect 18969 4672 18981 4675
rect 18840 4644 18981 4672
rect 18840 4632 18846 4644
rect 18969 4641 18981 4644
rect 19015 4641 19027 4675
rect 19334 4672 19340 4684
rect 19295 4644 19340 4672
rect 18969 4635 19027 4641
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 19702 4672 19708 4684
rect 19663 4644 19708 4672
rect 19702 4632 19708 4644
rect 19760 4632 19766 4684
rect 20070 4632 20076 4684
rect 20128 4672 20134 4684
rect 20952 4675 21010 4681
rect 20952 4672 20964 4675
rect 20128 4644 20964 4672
rect 20128 4632 20134 4644
rect 20952 4641 20964 4644
rect 20998 4672 21010 4675
rect 21450 4672 21456 4684
rect 20998 4644 21456 4672
rect 20998 4641 21010 4644
rect 20952 4635 21010 4641
rect 21450 4632 21456 4644
rect 21508 4632 21514 4684
rect 22370 4672 22376 4684
rect 22331 4644 22376 4672
rect 22370 4632 22376 4644
rect 22428 4632 22434 4684
rect 22738 4672 22744 4684
rect 22699 4644 22744 4672
rect 22738 4632 22744 4644
rect 22796 4632 22802 4684
rect 23290 4672 23296 4684
rect 23251 4644 23296 4672
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 23566 4672 23572 4684
rect 23527 4644 23572 4672
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 26602 4681 26608 4684
rect 26580 4675 26608 4681
rect 26580 4641 26592 4675
rect 26580 4635 26608 4641
rect 26602 4632 26608 4635
rect 26660 4632 26666 4684
rect 29178 4672 29184 4684
rect 29139 4644 29184 4672
rect 29178 4632 29184 4644
rect 29236 4632 29242 4684
rect 30650 4632 30656 4684
rect 30708 4681 30714 4684
rect 30708 4675 30746 4681
rect 30734 4641 30746 4675
rect 30708 4635 30746 4641
rect 30708 4632 30714 4635
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 16816 4576 18429 4604
rect 16816 4564 16822 4576
rect 18417 4573 18429 4576
rect 18463 4604 18475 4607
rect 18800 4604 18828 4632
rect 18463 4576 18828 4604
rect 18463 4573 18475 4576
rect 18417 4567 18475 4573
rect 21910 4564 21916 4616
rect 21968 4604 21974 4616
rect 24029 4607 24087 4613
rect 24029 4604 24041 4607
rect 21968 4576 24041 4604
rect 21968 4564 21974 4576
rect 24029 4573 24041 4576
rect 24075 4604 24087 4607
rect 24118 4604 24124 4616
rect 24075 4576 24124 4604
rect 24075 4573 24087 4576
rect 24029 4567 24087 4573
rect 24118 4564 24124 4576
rect 24176 4564 24182 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 24762 4604 24768 4616
rect 24627 4576 24768 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 26510 4496 26516 4548
rect 26568 4536 26574 4548
rect 27341 4539 27399 4545
rect 27341 4536 27353 4539
rect 26568 4508 27353 4536
rect 26568 4496 26574 4508
rect 27341 4505 27353 4508
rect 27387 4505 27399 4539
rect 27341 4499 27399 4505
rect 3513 4471 3571 4477
rect 3513 4437 3525 4471
rect 3559 4468 3571 4471
rect 3786 4468 3792 4480
rect 3559 4440 3792 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4525 4471 4583 4477
rect 4525 4468 4537 4471
rect 4212 4440 4537 4468
rect 4212 4428 4218 4440
rect 4525 4437 4537 4440
rect 4571 4437 4583 4471
rect 4525 4431 4583 4437
rect 9125 4471 9183 4477
rect 9125 4437 9137 4471
rect 9171 4468 9183 4471
rect 9582 4468 9588 4480
rect 9171 4440 9588 4468
rect 9171 4437 9183 4440
rect 9125 4431 9183 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 11514 4468 11520 4480
rect 11475 4440 11520 4468
rect 11514 4428 11520 4440
rect 11572 4468 11578 4480
rect 11882 4468 11888 4480
rect 11572 4440 11888 4468
rect 11572 4428 11578 4440
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 14240 4440 14657 4468
rect 14240 4428 14246 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 16022 4468 16028 4480
rect 15983 4440 16028 4468
rect 14645 4431 14703 4437
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 21821 4471 21879 4477
rect 21821 4437 21833 4471
rect 21867 4468 21879 4471
rect 22002 4468 22008 4480
rect 21867 4440 22008 4468
rect 21867 4437 21879 4440
rect 21821 4431 21879 4437
rect 22002 4428 22008 4440
rect 22060 4428 22066 4480
rect 22189 4471 22247 4477
rect 22189 4437 22201 4471
rect 22235 4468 22247 4471
rect 22370 4468 22376 4480
rect 22235 4440 22376 4468
rect 22235 4437 22247 4440
rect 22189 4431 22247 4437
rect 22370 4428 22376 4440
rect 22428 4428 22434 4480
rect 26786 4428 26792 4480
rect 26844 4468 26850 4480
rect 26973 4471 27031 4477
rect 26973 4468 26985 4471
rect 26844 4440 26985 4468
rect 26844 4428 26850 4440
rect 26973 4437 26985 4440
rect 27019 4437 27031 4471
rect 29546 4468 29552 4480
rect 29507 4440 29552 4468
rect 26973 4431 27031 4437
rect 29546 4428 29552 4440
rect 29604 4428 29610 4480
rect 30558 4428 30564 4480
rect 30616 4468 30622 4480
rect 30791 4471 30849 4477
rect 30791 4468 30803 4471
rect 30616 4440 30803 4468
rect 30616 4428 30622 4440
rect 30791 4437 30803 4440
rect 30837 4437 30849 4471
rect 30791 4431 30849 4437
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 2130 4224 2136 4276
rect 2188 4264 2194 4276
rect 2225 4267 2283 4273
rect 2225 4264 2237 4267
rect 2188 4236 2237 4264
rect 2188 4224 2194 4236
rect 2225 4233 2237 4236
rect 2271 4233 2283 4267
rect 2225 4227 2283 4233
rect 7929 4267 7987 4273
rect 7929 4233 7941 4267
rect 7975 4264 7987 4267
rect 8202 4264 8208 4276
rect 7975 4236 8208 4264
rect 7975 4233 7987 4236
rect 7929 4227 7987 4233
rect 2240 4060 2268 4227
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 10594 4264 10600 4276
rect 10555 4236 10600 4264
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 15470 4264 15476 4276
rect 15431 4236 15476 4264
rect 15470 4224 15476 4236
rect 15528 4224 15534 4276
rect 21269 4267 21327 4273
rect 21269 4233 21281 4267
rect 21315 4264 21327 4267
rect 21726 4264 21732 4276
rect 21315 4236 21732 4264
rect 21315 4233 21327 4236
rect 21269 4227 21327 4233
rect 21726 4224 21732 4236
rect 21784 4224 21790 4276
rect 22649 4267 22707 4273
rect 22649 4233 22661 4267
rect 22695 4264 22707 4267
rect 22738 4264 22744 4276
rect 22695 4236 22744 4264
rect 22695 4233 22707 4236
rect 22649 4227 22707 4233
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 26421 4267 26479 4273
rect 26421 4233 26433 4267
rect 26467 4264 26479 4267
rect 26602 4264 26608 4276
rect 26467 4236 26608 4264
rect 26467 4233 26479 4236
rect 26421 4227 26479 4233
rect 26602 4224 26608 4236
rect 26660 4224 26666 4276
rect 27614 4224 27620 4276
rect 27672 4264 27678 4276
rect 28077 4267 28135 4273
rect 28077 4264 28089 4267
rect 27672 4236 28089 4264
rect 27672 4224 27678 4236
rect 28077 4233 28089 4236
rect 28123 4233 28135 4267
rect 28077 4227 28135 4233
rect 29089 4267 29147 4273
rect 29089 4233 29101 4267
rect 29135 4264 29147 4267
rect 29178 4264 29184 4276
rect 29135 4236 29184 4264
rect 29135 4233 29147 4236
rect 29089 4227 29147 4233
rect 29178 4224 29184 4236
rect 29236 4224 29242 4276
rect 30650 4224 30656 4276
rect 30708 4264 30714 4276
rect 31294 4264 31300 4276
rect 30708 4236 31300 4264
rect 30708 4224 30714 4236
rect 31294 4224 31300 4236
rect 31352 4224 31358 4276
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 3602 4196 3608 4208
rect 3016 4168 3608 4196
rect 3016 4156 3022 4168
rect 3068 4069 3096 4168
rect 3602 4156 3608 4168
rect 3660 4156 3666 4208
rect 11517 4199 11575 4205
rect 11517 4165 11529 4199
rect 11563 4165 11575 4199
rect 11517 4159 11575 4165
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 4488 4100 4813 4128
rect 4488 4088 4494 4100
rect 4801 4097 4813 4100
rect 4847 4128 4859 4131
rect 5074 4128 5080 4140
rect 4847 4100 5080 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5442 4128 5448 4140
rect 5403 4100 5448 4128
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 6052 4100 7573 4128
rect 6052 4088 6058 4100
rect 7561 4097 7573 4100
rect 7607 4128 7619 4131
rect 11532 4128 11560 4159
rect 17310 4156 17316 4208
rect 17368 4196 17374 4208
rect 23566 4196 23572 4208
rect 17368 4168 18092 4196
rect 17368 4156 17374 4168
rect 17129 4131 17187 4137
rect 7607 4100 9168 4128
rect 11532 4100 13124 4128
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2240 4032 2421 4060
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4029 3111 4063
rect 3418 4060 3424 4072
rect 3379 4032 3424 4060
rect 3053 4023 3111 4029
rect 3418 4020 3424 4032
rect 3476 4020 3482 4072
rect 3786 4060 3792 4072
rect 3747 4032 3792 4060
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 9140 4069 9168 4100
rect 13096 4072 13124 4100
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17954 4128 17960 4140
rect 17175 4100 17960 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18064 4128 18092 4168
rect 23400 4168 23572 4196
rect 19797 4131 19855 4137
rect 19797 4128 19809 4131
rect 18064 4100 19809 4128
rect 18892 4072 18920 4100
rect 19797 4097 19809 4100
rect 19843 4097 19855 4131
rect 19797 4091 19855 4097
rect 20438 4088 20444 4140
rect 20496 4128 20502 4140
rect 21634 4128 21640 4140
rect 20496 4100 21640 4128
rect 20496 4088 20502 4100
rect 21634 4088 21640 4100
rect 21692 4128 21698 4140
rect 21913 4131 21971 4137
rect 21913 4128 21925 4131
rect 21692 4100 21925 4128
rect 21692 4088 21698 4100
rect 21913 4097 21925 4100
rect 21959 4128 21971 4131
rect 22370 4128 22376 4140
rect 21959 4100 22376 4128
rect 21959 4097 21971 4100
rect 21913 4091 21971 4097
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22922 4088 22928 4140
rect 22980 4128 22986 4140
rect 23017 4131 23075 4137
rect 23017 4128 23029 4131
rect 22980 4100 23029 4128
rect 22980 4088 22986 4100
rect 23017 4097 23029 4100
rect 23063 4128 23075 4131
rect 23400 4128 23428 4168
rect 23566 4156 23572 4168
rect 23624 4156 23630 4208
rect 23063 4100 23428 4128
rect 23063 4097 23075 4100
rect 23017 4091 23075 4097
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 23661 4131 23719 4137
rect 23661 4128 23673 4131
rect 23532 4100 23673 4128
rect 23532 4088 23538 4100
rect 23661 4097 23673 4100
rect 23707 4097 23719 4131
rect 30101 4131 30159 4137
rect 30101 4128 30113 4131
rect 23661 4091 23719 4097
rect 27448 4100 30113 4128
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 8260 4032 8401 4060
rect 8260 4020 8266 4032
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4029 9459 4063
rect 9582 4060 9588 4072
rect 9543 4032 9588 4060
rect 9401 4023 9459 4029
rect 2682 3952 2688 4004
rect 2740 3992 2746 4004
rect 3436 3992 3464 4020
rect 2740 3964 3464 3992
rect 4893 3995 4951 4001
rect 2740 3952 2746 3964
rect 4893 3961 4905 3995
rect 4939 3992 4951 3995
rect 4982 3992 4988 4004
rect 4939 3964 4988 3992
rect 4939 3961 4951 3964
rect 4893 3955 4951 3961
rect 4982 3952 4988 3964
rect 5040 3952 5046 4004
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 5721 3995 5779 4001
rect 5721 3992 5733 3995
rect 5224 3964 5733 3992
rect 5224 3952 5230 3964
rect 5721 3961 5733 3964
rect 5767 3961 5779 3995
rect 5721 3955 5779 3961
rect 6181 3995 6239 4001
rect 6181 3961 6193 3995
rect 6227 3992 6239 3995
rect 6546 3992 6552 4004
rect 6227 3964 6552 3992
rect 6227 3961 6239 3964
rect 6181 3955 6239 3961
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 8018 3992 8024 4004
rect 7239 3964 8024 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 8018 3952 8024 3964
rect 8076 3992 8082 4004
rect 9140 3992 9168 4023
rect 9306 3992 9312 4004
rect 8076 3964 8524 3992
rect 9140 3964 9312 3992
rect 8076 3952 8082 3964
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 2498 3924 2504 3936
rect 2459 3896 2504 3924
rect 2498 3884 2504 3896
rect 2556 3884 2562 3936
rect 4246 3924 4252 3936
rect 4207 3896 4252 3924
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3924 4675 3927
rect 5994 3924 6000 3936
rect 4663 3896 6000 3924
rect 4663 3893 4675 3896
rect 4617 3887 4675 3893
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6454 3924 6460 3936
rect 6415 3896 6460 3924
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 8202 3924 8208 3936
rect 8163 3896 8208 3924
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8496 3933 8524 3964
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3893 8539 3927
rect 8481 3887 8539 3893
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 9416 3924 9444 4023
rect 9582 4020 9588 4032
rect 9640 4060 9646 4072
rect 10870 4060 10876 4072
rect 9640 4032 10876 4060
rect 9640 4020 9646 4032
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11379 4032 11836 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11808 3936 11836 4032
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 11940 4032 12449 4060
rect 11940 4020 11946 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 13078 4060 13084 4072
rect 12991 4032 13084 4060
rect 12437 4023 12495 4029
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13262 4060 13268 4072
rect 13223 4032 13268 4060
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13630 4060 13636 4072
rect 13591 4032 13636 4060
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15528 4032 15669 4060
rect 15528 4020 15534 4032
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 15657 4023 15715 4029
rect 16393 4063 16451 4069
rect 16393 4029 16405 4063
rect 16439 4029 16451 4063
rect 16666 4060 16672 4072
rect 16627 4032 16672 4060
rect 16393 4023 16451 4029
rect 13096 3992 13124 4020
rect 14829 3995 14887 4001
rect 14829 3992 14841 3995
rect 13096 3964 14841 3992
rect 14829 3961 14841 3964
rect 14875 3992 14887 3995
rect 16408 3992 16436 4023
rect 16666 4020 16672 4032
rect 16724 4020 16730 4072
rect 17034 4060 17040 4072
rect 16995 4032 17040 4060
rect 17034 4020 17040 4032
rect 17092 4020 17098 4072
rect 18141 4063 18199 4069
rect 18141 4060 18153 4063
rect 17788 4032 18153 4060
rect 16758 3992 16764 4004
rect 14875 3964 16764 3992
rect 14875 3961 14887 3964
rect 14829 3955 14887 3961
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 10226 3924 10232 3936
rect 9180 3896 10232 3924
rect 9180 3884 9186 3896
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 11790 3924 11796 3936
rect 11751 3896 11796 3924
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12250 3924 12256 3936
rect 12211 3896 12256 3924
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 13633 3927 13691 3933
rect 13633 3924 13645 3927
rect 13596 3896 13645 3924
rect 13596 3884 13602 3896
rect 13633 3893 13645 3896
rect 13679 3893 13691 3927
rect 13633 3887 13691 3893
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 14642 3924 14648 3936
rect 14507 3896 14648 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 15197 3927 15255 3933
rect 15197 3893 15209 3927
rect 15243 3924 15255 3927
rect 15378 3924 15384 3936
rect 15243 3896 15384 3924
rect 15243 3893 15255 3896
rect 15197 3887 15255 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 17402 3924 17408 3936
rect 17363 3896 17408 3924
rect 17402 3884 17408 3896
rect 17460 3924 17466 3936
rect 17788 3933 17816 4032
rect 18141 4029 18153 4032
rect 18187 4060 18199 4063
rect 18506 4060 18512 4072
rect 18187 4032 18512 4060
rect 18187 4029 18199 4032
rect 18141 4023 18199 4029
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 18782 4060 18788 4072
rect 18743 4032 18788 4060
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 18874 4020 18880 4072
rect 18932 4060 18938 4072
rect 19242 4060 19248 4072
rect 18932 4032 19025 4060
rect 19203 4032 19248 4060
rect 18932 4020 18938 4032
rect 19242 4020 19248 4032
rect 19300 4060 19306 4072
rect 19702 4060 19708 4072
rect 19300 4032 19708 4060
rect 19300 4020 19306 4032
rect 19702 4020 19708 4032
rect 19760 4020 19766 4072
rect 20346 4060 20352 4072
rect 20307 4032 20352 4060
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 22094 4020 22100 4072
rect 22152 4060 22158 4072
rect 24581 4063 24639 4069
rect 22152 4032 22197 4060
rect 22152 4020 22158 4032
rect 24581 4029 24593 4063
rect 24627 4060 24639 4063
rect 24670 4060 24676 4072
rect 24627 4032 24676 4060
rect 24627 4029 24639 4032
rect 24581 4023 24639 4029
rect 24670 4020 24676 4032
rect 24728 4020 24734 4072
rect 25314 4020 25320 4072
rect 25372 4060 25378 4072
rect 25498 4069 25504 4072
rect 25444 4063 25504 4069
rect 25444 4060 25456 4063
rect 25372 4032 25456 4060
rect 25372 4020 25378 4032
rect 25444 4029 25456 4032
rect 25490 4029 25504 4063
rect 25444 4023 25504 4029
rect 25498 4020 25504 4023
rect 25556 4060 25562 4072
rect 25869 4063 25927 4069
rect 25869 4060 25881 4063
rect 25556 4032 25881 4060
rect 25556 4020 25562 4032
rect 25869 4029 25881 4032
rect 25915 4029 25927 4063
rect 26510 4060 26516 4072
rect 26471 4032 26516 4060
rect 25869 4023 25927 4029
rect 26510 4020 26516 4032
rect 26568 4020 26574 4072
rect 27448 4069 27476 4100
rect 30101 4097 30113 4100
rect 30147 4128 30159 4131
rect 30466 4128 30472 4140
rect 30147 4100 30472 4128
rect 30147 4097 30159 4100
rect 30101 4091 30159 4097
rect 30466 4088 30472 4100
rect 30524 4088 30530 4140
rect 27433 4063 27491 4069
rect 27433 4029 27445 4063
rect 27479 4029 27491 4063
rect 27433 4023 27491 4029
rect 29086 4020 29092 4072
rect 29144 4060 29150 4072
rect 29308 4063 29366 4069
rect 29308 4060 29320 4063
rect 29144 4032 29320 4060
rect 29144 4020 29150 4032
rect 29308 4029 29320 4032
rect 29354 4060 29366 4063
rect 29730 4060 29736 4072
rect 29354 4032 29736 4060
rect 29354 4029 29366 4032
rect 29308 4023 29366 4029
rect 29730 4020 29736 4032
rect 29788 4020 29794 4072
rect 20257 3995 20315 4001
rect 20257 3961 20269 3995
rect 20303 3992 20315 3995
rect 20711 3995 20769 4001
rect 20711 3992 20723 3995
rect 20303 3964 20723 3992
rect 20303 3961 20315 3964
rect 20257 3955 20315 3961
rect 20711 3961 20723 3964
rect 20757 3992 20769 3995
rect 20806 3992 20812 4004
rect 20757 3964 20812 3992
rect 20757 3961 20769 3964
rect 20711 3955 20769 3961
rect 20806 3952 20812 3964
rect 20864 3952 20870 4004
rect 21450 3952 21456 4004
rect 21508 3992 21514 4004
rect 21637 3995 21695 4001
rect 21637 3992 21649 3995
rect 21508 3964 21649 3992
rect 21508 3952 21514 3964
rect 21637 3961 21649 3964
rect 21683 3992 21695 3995
rect 22830 3992 22836 4004
rect 21683 3964 22836 3992
rect 21683 3961 21695 3964
rect 21637 3955 21695 3961
rect 22830 3952 22836 3964
rect 22888 3952 22894 4004
rect 23982 3995 24040 4001
rect 23982 3992 23994 3995
rect 23492 3964 23994 3992
rect 23492 3936 23520 3964
rect 23982 3961 23994 3964
rect 24028 3992 24040 3995
rect 24028 3964 24716 3992
rect 24028 3961 24040 3964
rect 23982 3955 24040 3961
rect 17773 3927 17831 3933
rect 17773 3924 17785 3927
rect 17460 3896 17785 3924
rect 17460 3884 17466 3896
rect 17773 3893 17785 3896
rect 17819 3893 17831 3927
rect 17773 3887 17831 3893
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18141 3927 18199 3933
rect 18141 3924 18153 3927
rect 17920 3896 18153 3924
rect 17920 3884 17926 3896
rect 18141 3893 18153 3896
rect 18187 3893 18199 3927
rect 18141 3887 18199 3893
rect 22281 3927 22339 3933
rect 22281 3893 22293 3927
rect 22327 3924 22339 3927
rect 22554 3924 22560 3936
rect 22327 3896 22560 3924
rect 22327 3893 22339 3896
rect 22281 3887 22339 3893
rect 22554 3884 22560 3896
rect 22612 3924 22618 3936
rect 23290 3924 23296 3936
rect 22612 3896 23296 3924
rect 22612 3884 22618 3896
rect 23290 3884 23296 3896
rect 23348 3884 23354 3936
rect 23474 3924 23480 3936
rect 23435 3896 23480 3924
rect 23474 3884 23480 3896
rect 23532 3884 23538 3936
rect 24688 3924 24716 3964
rect 24762 3952 24768 4004
rect 24820 3992 24826 4004
rect 25225 3995 25283 4001
rect 25225 3992 25237 3995
rect 24820 3964 25237 3992
rect 24820 3952 24826 3964
rect 25225 3961 25237 3964
rect 25271 3961 25283 3995
rect 25225 3955 25283 3961
rect 26786 3952 26792 4004
rect 26844 4001 26850 4004
rect 26844 3995 26892 4001
rect 26844 3961 26846 3995
rect 26880 3961 26892 3995
rect 26844 3955 26892 3961
rect 26844 3952 26850 3955
rect 27706 3952 27712 4004
rect 27764 3952 27770 4004
rect 29411 3995 29469 4001
rect 29411 3961 29423 3995
rect 29457 3992 29469 3995
rect 30374 3992 30380 4004
rect 29457 3964 30380 3992
rect 29457 3961 29469 3964
rect 29411 3955 29469 3961
rect 30374 3952 30380 3964
rect 30432 3952 30438 4004
rect 30466 3952 30472 4004
rect 30524 3992 30530 4004
rect 31018 3992 31024 4004
rect 30524 3964 30569 3992
rect 30979 3964 31024 3992
rect 30524 3952 30530 3964
rect 31018 3952 31024 3964
rect 31076 3952 31082 4004
rect 24854 3924 24860 3936
rect 24688 3896 24860 3924
rect 24854 3884 24860 3896
rect 24912 3884 24918 3936
rect 25547 3927 25605 3933
rect 25547 3893 25559 3927
rect 25593 3924 25605 3927
rect 25866 3924 25872 3936
rect 25593 3896 25872 3924
rect 25593 3893 25605 3896
rect 25547 3887 25605 3893
rect 25866 3884 25872 3896
rect 25924 3884 25930 3936
rect 27724 3924 27752 3952
rect 27801 3927 27859 3933
rect 27801 3924 27813 3927
rect 27724 3896 27813 3924
rect 27801 3893 27813 3896
rect 27847 3924 27859 3927
rect 29270 3924 29276 3936
rect 27847 3896 29276 3924
rect 27847 3893 27859 3896
rect 27801 3887 27859 3893
rect 29270 3884 29276 3896
rect 29328 3884 29334 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 1765 3723 1823 3729
rect 1765 3689 1777 3723
rect 1811 3720 1823 3723
rect 1854 3720 1860 3732
rect 1811 3692 1860 3720
rect 1811 3689 1823 3692
rect 1765 3683 1823 3689
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 2590 3680 2596 3732
rect 2648 3729 2654 3732
rect 2648 3723 2697 3729
rect 2648 3689 2651 3723
rect 2685 3689 2697 3723
rect 2648 3683 2697 3689
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3418 3720 3424 3732
rect 3099 3692 3424 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 2648 3680 2654 3683
rect 2133 3655 2191 3661
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 3068 3652 3096 3683
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 4801 3723 4859 3729
rect 4801 3689 4813 3723
rect 4847 3720 4859 3723
rect 4982 3720 4988 3732
rect 4847 3692 4988 3720
rect 4847 3689 4859 3692
rect 4801 3683 4859 3689
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 6638 3720 6644 3732
rect 5132 3692 5177 3720
rect 6599 3692 6644 3720
rect 5132 3680 5138 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 9122 3720 9128 3732
rect 9083 3692 9128 3720
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3720 9919 3723
rect 11514 3720 11520 3732
rect 9907 3692 11520 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 12526 3720 12532 3732
rect 12439 3692 12532 3720
rect 12526 3680 12532 3692
rect 12584 3720 12590 3732
rect 13262 3720 13268 3732
rect 12584 3692 13268 3720
rect 12584 3680 12590 3692
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 15528 3692 16313 3720
rect 15528 3680 15534 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 16758 3720 16764 3732
rect 16719 3692 16764 3720
rect 16301 3683 16359 3689
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 18840 3692 19257 3720
rect 18840 3680 18846 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 19245 3683 19303 3689
rect 20257 3723 20315 3729
rect 20257 3689 20269 3723
rect 20303 3720 20315 3723
rect 21910 3720 21916 3732
rect 20303 3692 21916 3720
rect 20303 3689 20315 3692
rect 20257 3683 20315 3689
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 22005 3723 22063 3729
rect 22005 3689 22017 3723
rect 22051 3720 22063 3723
rect 22370 3720 22376 3732
rect 22051 3692 22376 3720
rect 22051 3689 22063 3692
rect 22005 3683 22063 3689
rect 22370 3680 22376 3692
rect 22428 3720 22434 3732
rect 25866 3720 25872 3732
rect 22428 3692 22692 3720
rect 22428 3680 22434 3692
rect 8754 3652 8760 3664
rect 2179 3624 3096 3652
rect 8667 3624 8760 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 8754 3612 8760 3624
rect 8812 3652 8818 3664
rect 10594 3652 10600 3664
rect 8812 3624 10600 3652
rect 8812 3612 8818 3624
rect 10594 3612 10600 3624
rect 10652 3612 10658 3664
rect 11532 3652 11560 3680
rect 15105 3655 15163 3661
rect 11532 3624 15056 3652
rect 2568 3587 2626 3593
rect 2568 3553 2580 3587
rect 2614 3584 2626 3587
rect 2774 3584 2780 3596
rect 2614 3556 2780 3584
rect 2614 3553 2626 3556
rect 2568 3547 2626 3553
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 3421 3587 3479 3593
rect 3421 3553 3433 3587
rect 3467 3584 3479 3587
rect 3602 3584 3608 3596
rect 3467 3556 3608 3584
rect 3467 3553 3479 3556
rect 3421 3547 3479 3553
rect 3602 3544 3608 3556
rect 3660 3544 3666 3596
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 5224 3556 5273 3584
rect 5224 3544 5230 3556
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5994 3584 6000 3596
rect 5955 3556 6000 3584
rect 5261 3547 5319 3553
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3553 6331 3587
rect 6638 3584 6644 3596
rect 6599 3556 6644 3584
rect 6273 3547 6331 3553
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 6288 3516 6316 3547
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 9030 3584 9036 3596
rect 8711 3556 9036 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 9030 3544 9036 3556
rect 9088 3584 9094 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9088 3556 9689 3584
rect 9088 3544 9094 3556
rect 9677 3553 9689 3556
rect 9723 3584 9735 3587
rect 9766 3584 9772 3596
rect 9723 3556 9772 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 10134 3584 10140 3596
rect 10095 3556 10140 3584
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 11790 3584 11796 3596
rect 11751 3556 11796 3584
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 14274 3584 14280 3596
rect 14235 3556 14280 3584
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 15028 3584 15056 3624
rect 15105 3621 15117 3655
rect 15151 3652 15163 3655
rect 15286 3652 15292 3664
rect 15151 3624 15292 3652
rect 15151 3621 15163 3624
rect 15105 3615 15163 3621
rect 15286 3612 15292 3624
rect 15344 3612 15350 3664
rect 16025 3655 16083 3661
rect 16025 3621 16037 3655
rect 16071 3652 16083 3655
rect 16482 3652 16488 3664
rect 16071 3624 16488 3652
rect 16071 3621 16083 3624
rect 16025 3615 16083 3621
rect 16482 3612 16488 3624
rect 16540 3612 16546 3664
rect 18969 3655 19027 3661
rect 18969 3621 18981 3655
rect 19015 3652 19027 3655
rect 20346 3652 20352 3664
rect 19015 3624 20352 3652
rect 19015 3621 19027 3624
rect 18969 3615 19027 3621
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 20993 3655 21051 3661
rect 20993 3652 21005 3655
rect 20680 3624 21005 3652
rect 20680 3612 20686 3624
rect 20993 3621 21005 3624
rect 21039 3621 21051 3655
rect 20993 3615 21051 3621
rect 21085 3655 21143 3661
rect 21085 3621 21097 3655
rect 21131 3652 21143 3655
rect 21266 3652 21272 3664
rect 21131 3624 21272 3652
rect 21131 3621 21143 3624
rect 21085 3615 21143 3621
rect 21266 3612 21272 3624
rect 21324 3612 21330 3664
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 15028 3556 17325 3584
rect 17313 3553 17325 3556
rect 17359 3584 17371 3587
rect 17402 3584 17408 3596
rect 17359 3556 17408 3584
rect 17359 3553 17371 3556
rect 17313 3547 17371 3553
rect 17402 3544 17408 3556
rect 17460 3584 17466 3596
rect 17497 3587 17555 3593
rect 17497 3584 17509 3587
rect 17460 3556 17509 3584
rect 17460 3544 17466 3556
rect 17497 3553 17509 3556
rect 17543 3553 17555 3587
rect 17954 3584 17960 3596
rect 17915 3556 17960 3584
rect 17497 3547 17555 3553
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 18322 3584 18328 3596
rect 18283 3556 18328 3584
rect 18322 3544 18328 3556
rect 18380 3544 18386 3596
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3584 18751 3587
rect 19242 3584 19248 3596
rect 18739 3556 19248 3584
rect 18739 3553 18751 3556
rect 18693 3547 18751 3553
rect 11882 3516 11888 3528
rect 5500 3488 7972 3516
rect 11843 3488 11888 3516
rect 5500 3476 5506 3488
rect 7944 3457 7972 3488
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 14550 3516 14556 3528
rect 14415 3488 14556 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 14550 3476 14556 3488
rect 14608 3516 14614 3528
rect 15654 3516 15660 3528
rect 14608 3488 15660 3516
rect 14608 3476 14614 3488
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 18708 3516 18736 3547
rect 19242 3544 19248 3556
rect 19300 3584 19306 3596
rect 22664 3593 22692 3692
rect 24964 3692 25872 3720
rect 23937 3655 23995 3661
rect 23937 3621 23949 3655
rect 23983 3652 23995 3655
rect 24762 3652 24768 3664
rect 23983 3624 24768 3652
rect 23983 3621 23995 3624
rect 23937 3615 23995 3621
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 24964 3661 24992 3692
rect 25866 3680 25872 3692
rect 25924 3680 25930 3732
rect 28169 3723 28227 3729
rect 28169 3689 28181 3723
rect 28215 3720 28227 3723
rect 28258 3720 28264 3732
rect 28215 3692 28264 3720
rect 28215 3689 28227 3692
rect 28169 3683 28227 3689
rect 28258 3680 28264 3692
rect 28316 3680 28322 3732
rect 30374 3720 30380 3732
rect 30335 3692 30380 3720
rect 30374 3680 30380 3692
rect 30432 3680 30438 3732
rect 30466 3680 30472 3732
rect 30524 3720 30530 3732
rect 30524 3692 32260 3720
rect 30524 3680 30530 3692
rect 24949 3655 25007 3661
rect 24949 3621 24961 3655
rect 24995 3621 25007 3655
rect 24949 3615 25007 3621
rect 25041 3655 25099 3661
rect 25041 3621 25053 3655
rect 25087 3652 25099 3655
rect 25406 3652 25412 3664
rect 25087 3624 25412 3652
rect 25087 3621 25099 3624
rect 25041 3615 25099 3621
rect 25406 3612 25412 3624
rect 25464 3652 25470 3664
rect 26142 3652 26148 3664
rect 25464 3624 26148 3652
rect 25464 3612 25470 3624
rect 26142 3612 26148 3624
rect 26200 3612 26206 3664
rect 26326 3612 26332 3664
rect 26384 3652 26390 3664
rect 26786 3652 26792 3664
rect 26384 3624 26792 3652
rect 26384 3612 26390 3624
rect 26786 3612 26792 3624
rect 26844 3661 26850 3664
rect 26844 3655 26892 3661
rect 26844 3621 26846 3655
rect 26880 3621 26892 3655
rect 28276 3652 28304 3680
rect 28353 3655 28411 3661
rect 28353 3652 28365 3655
rect 28276 3624 28365 3652
rect 26844 3615 26892 3621
rect 28353 3621 28365 3624
rect 28399 3621 28411 3655
rect 28353 3615 28411 3621
rect 28445 3655 28503 3661
rect 28445 3621 28457 3655
rect 28491 3652 28503 3655
rect 28534 3652 28540 3664
rect 28491 3624 28540 3652
rect 28491 3621 28503 3624
rect 28445 3615 28503 3621
rect 26844 3612 26850 3615
rect 28534 3612 28540 3624
rect 28592 3652 28598 3664
rect 29178 3652 29184 3664
rect 28592 3624 29184 3652
rect 28592 3612 28598 3624
rect 29178 3612 29184 3624
rect 29236 3612 29242 3664
rect 30009 3655 30067 3661
rect 30009 3621 30021 3655
rect 30055 3652 30067 3655
rect 30558 3652 30564 3664
rect 30055 3624 30564 3652
rect 30055 3621 30067 3624
rect 30009 3615 30067 3621
rect 30558 3612 30564 3624
rect 30616 3612 30622 3664
rect 30650 3612 30656 3664
rect 30708 3652 30714 3664
rect 32125 3655 32183 3661
rect 32125 3652 32137 3655
rect 30708 3624 32137 3652
rect 30708 3612 30714 3624
rect 32125 3621 32137 3624
rect 32171 3621 32183 3655
rect 32125 3615 32183 3621
rect 32232 3596 32260 3692
rect 19613 3587 19671 3593
rect 19613 3584 19625 3587
rect 19300 3556 19625 3584
rect 19300 3544 19306 3556
rect 19613 3553 19625 3556
rect 19659 3553 19671 3587
rect 19613 3547 19671 3553
rect 22649 3587 22707 3593
rect 22649 3553 22661 3587
rect 22695 3553 22707 3587
rect 22649 3547 22707 3553
rect 19794 3516 19800 3528
rect 17184 3488 18736 3516
rect 19755 3488 19800 3516
rect 17184 3476 17190 3488
rect 19794 3476 19800 3488
rect 19852 3476 19858 3528
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3485 21327 3519
rect 22664 3516 22692 3547
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 22925 3587 22983 3593
rect 22925 3584 22937 3587
rect 22796 3556 22937 3584
rect 22796 3544 22802 3556
rect 22925 3553 22937 3556
rect 22971 3553 22983 3587
rect 22925 3547 22983 3553
rect 23290 3544 23296 3596
rect 23348 3584 23354 3596
rect 23477 3587 23535 3593
rect 23477 3584 23489 3587
rect 23348 3556 23489 3584
rect 23348 3544 23354 3556
rect 23477 3553 23489 3556
rect 23523 3584 23535 3587
rect 23750 3584 23756 3596
rect 23523 3556 23612 3584
rect 23711 3556 23756 3584
rect 23523 3553 23535 3556
rect 23477 3547 23535 3553
rect 22664 3488 23520 3516
rect 21269 3479 21327 3485
rect 7929 3451 7987 3457
rect 7929 3417 7941 3451
rect 7975 3448 7987 3451
rect 9122 3448 9128 3460
rect 7975 3420 9128 3448
rect 7975 3417 7987 3420
rect 7929 3411 7987 3417
rect 9122 3408 9128 3420
rect 9180 3408 9186 3460
rect 11054 3448 11060 3460
rect 11015 3420 11060 3448
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 15378 3408 15384 3460
rect 15436 3457 15442 3460
rect 15436 3451 15485 3457
rect 15436 3417 15439 3451
rect 15473 3417 15485 3451
rect 15562 3448 15568 3460
rect 15523 3420 15568 3448
rect 15436 3411 15485 3417
rect 15436 3408 15442 3411
rect 15562 3408 15568 3420
rect 15620 3408 15626 3460
rect 20530 3408 20536 3460
rect 20588 3448 20594 3460
rect 21284 3448 21312 3479
rect 22278 3448 22284 3460
rect 20588 3420 22284 3448
rect 20588 3408 20594 3420
rect 22278 3408 22284 3420
rect 22336 3408 22342 3460
rect 12897 3383 12955 3389
rect 12897 3349 12909 3383
rect 12943 3380 12955 3383
rect 13265 3383 13323 3389
rect 13265 3380 13277 3383
rect 12943 3352 13277 3380
rect 12943 3349 12955 3352
rect 12897 3343 12955 3349
rect 13265 3349 13277 3352
rect 13311 3380 13323 3383
rect 13630 3380 13636 3392
rect 13311 3352 13636 3380
rect 13311 3349 13323 3352
rect 13265 3343 13323 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 14737 3383 14795 3389
rect 14737 3349 14749 3383
rect 14783 3380 14795 3383
rect 14918 3380 14924 3392
rect 14783 3352 14924 3380
rect 14783 3349 14795 3352
rect 14737 3343 14795 3349
rect 14918 3340 14924 3352
rect 14976 3380 14982 3392
rect 15580 3380 15608 3408
rect 23492 3392 23520 3488
rect 23584 3448 23612 3556
rect 23750 3544 23756 3556
rect 23808 3544 23814 3596
rect 32214 3584 32220 3596
rect 32175 3556 32220 3584
rect 32214 3544 32220 3556
rect 32272 3544 32278 3596
rect 24946 3476 24952 3528
rect 25004 3516 25010 3528
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 25004 3488 25237 3516
rect 25004 3476 25010 3488
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 26418 3476 26424 3528
rect 26476 3516 26482 3528
rect 26513 3519 26571 3525
rect 26513 3516 26525 3519
rect 26476 3488 26525 3516
rect 26476 3476 26482 3488
rect 26513 3485 26525 3488
rect 26559 3485 26571 3519
rect 28997 3519 29055 3525
rect 28997 3516 29009 3519
rect 26513 3479 26571 3485
rect 28920 3488 29009 3516
rect 28920 3460 28948 3488
rect 28997 3485 29009 3488
rect 29043 3516 29055 3519
rect 29273 3519 29331 3525
rect 29273 3516 29285 3519
rect 29043 3488 29285 3516
rect 29043 3485 29055 3488
rect 28997 3479 29055 3485
rect 29273 3485 29285 3488
rect 29319 3485 29331 3519
rect 31018 3516 31024 3528
rect 30979 3488 31024 3516
rect 29273 3479 29331 3485
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 23584 3420 24624 3448
rect 24596 3392 24624 3420
rect 28902 3408 28908 3460
rect 28960 3408 28966 3460
rect 14976 3352 15608 3380
rect 14976 3340 14982 3352
rect 20622 3340 20628 3392
rect 20680 3380 20686 3392
rect 20717 3383 20775 3389
rect 20717 3380 20729 3383
rect 20680 3352 20729 3380
rect 20680 3340 20686 3352
rect 20717 3349 20729 3352
rect 20763 3349 20775 3383
rect 20717 3343 20775 3349
rect 20806 3340 20812 3392
rect 20864 3380 20870 3392
rect 22370 3380 22376 3392
rect 20864 3352 22376 3380
rect 20864 3340 20870 3352
rect 22370 3340 22376 3352
rect 22428 3340 22434 3392
rect 23474 3340 23480 3392
rect 23532 3380 23538 3392
rect 24213 3383 24271 3389
rect 24213 3380 24225 3383
rect 23532 3352 24225 3380
rect 23532 3340 23538 3352
rect 24213 3349 24225 3352
rect 24259 3349 24271 3383
rect 24578 3380 24584 3392
rect 24539 3352 24584 3380
rect 24213 3343 24271 3349
rect 24578 3340 24584 3352
rect 24636 3340 24642 3392
rect 26234 3380 26240 3392
rect 26195 3352 26240 3380
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 27430 3380 27436 3392
rect 27391 3352 27436 3380
rect 27430 3340 27436 3352
rect 27488 3340 27494 3392
rect 32490 3340 32496 3392
rect 32548 3380 32554 3392
rect 33137 3383 33195 3389
rect 33137 3380 33149 3383
rect 32548 3352 33149 3380
rect 32548 3340 32554 3352
rect 33137 3349 33149 3352
rect 33183 3349 33195 3383
rect 33137 3343 33195 3349
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 1762 3176 1768 3188
rect 1723 3148 1768 3176
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 2593 3179 2651 3185
rect 2593 3145 2605 3179
rect 2639 3176 2651 3179
rect 2774 3176 2780 3188
rect 2639 3148 2780 3176
rect 2639 3145 2651 3148
rect 2593 3139 2651 3145
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 6638 3176 6644 3188
rect 4571 3148 6644 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 1854 3068 1860 3120
rect 1912 3108 1918 3120
rect 2133 3111 2191 3117
rect 2133 3108 2145 3111
rect 1912 3080 2145 3108
rect 1912 3068 1918 3080
rect 2133 3077 2145 3080
rect 2179 3077 2191 3111
rect 4062 3108 4068 3120
rect 4023 3080 4068 3108
rect 2133 3071 2191 3077
rect 2148 3040 2176 3071
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 2148 3012 3832 3040
rect 3804 2984 3832 3012
rect 1762 2932 1768 2984
rect 1820 2972 1826 2984
rect 2958 2972 2964 2984
rect 1820 2944 2964 2972
rect 1820 2932 1826 2944
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2941 3387 2975
rect 3510 2972 3516 2984
rect 3471 2944 3516 2972
rect 3329 2935 3387 2941
rect 3234 2864 3240 2916
rect 3292 2904 3298 2916
rect 3344 2904 3372 2935
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3786 2932 3792 2984
rect 3844 2972 3850 2984
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 3844 2944 4077 2972
rect 3844 2932 3850 2944
rect 4065 2941 4077 2944
rect 4111 2972 4123 2975
rect 4540 2972 4568 3139
rect 6638 3136 6644 3148
rect 6696 3176 6702 3188
rect 7193 3179 7251 3185
rect 7193 3176 7205 3179
rect 6696 3148 7205 3176
rect 6696 3136 6702 3148
rect 7193 3145 7205 3148
rect 7239 3145 7251 3179
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 7193 3139 7251 3145
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 13725 3179 13783 3185
rect 13725 3145 13737 3179
rect 13771 3176 13783 3179
rect 14274 3176 14280 3188
rect 13771 3148 14280 3176
rect 13771 3145 13783 3148
rect 13725 3139 13783 3145
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14550 3185 14556 3188
rect 14534 3179 14556 3185
rect 14534 3145 14546 3179
rect 14534 3139 14556 3145
rect 14550 3136 14556 3139
rect 14608 3136 14614 3188
rect 14645 3179 14703 3185
rect 14645 3145 14657 3179
rect 14691 3176 14703 3179
rect 15286 3176 15292 3188
rect 14691 3148 15292 3176
rect 14691 3145 14703 3148
rect 14645 3139 14703 3145
rect 5166 3068 5172 3120
rect 5224 3108 5230 3120
rect 5813 3111 5871 3117
rect 5813 3108 5825 3111
rect 5224 3080 5825 3108
rect 5224 3068 5230 3080
rect 5813 3077 5825 3080
rect 5859 3108 5871 3111
rect 7469 3111 7527 3117
rect 7469 3108 7481 3111
rect 5859 3080 7481 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 7469 3077 7481 3080
rect 7515 3077 7527 3111
rect 7469 3071 7527 3077
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 5994 3040 6000 3052
rect 4939 3012 6000 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 5994 3000 6000 3012
rect 6052 3000 6058 3052
rect 4111 2944 4568 2972
rect 4985 2975 5043 2981
rect 4111 2941 4123 2944
rect 4065 2935 4123 2941
rect 4985 2941 4997 2975
rect 5031 2972 5043 2975
rect 6641 2975 6699 2981
rect 5031 2944 5396 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 3602 2904 3608 2916
rect 3292 2876 3608 2904
rect 3292 2864 3298 2876
rect 3602 2864 3608 2876
rect 3660 2864 3666 2916
rect 5368 2848 5396 2944
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 7006 2972 7012 2984
rect 6687 2944 7012 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 7484 2972 7512 3071
rect 13998 3068 14004 3120
rect 14056 3108 14062 3120
rect 14660 3108 14688 3139
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 15473 3179 15531 3185
rect 15473 3145 15485 3179
rect 15519 3176 15531 3179
rect 15562 3176 15568 3188
rect 15519 3148 15568 3176
rect 15519 3145 15531 3148
rect 15473 3139 15531 3145
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 17126 3176 17132 3188
rect 17087 3148 17132 3176
rect 17126 3136 17132 3148
rect 17184 3176 17190 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 17184 3148 17509 3176
rect 17184 3136 17190 3148
rect 17497 3145 17509 3148
rect 17543 3176 17555 3179
rect 17954 3176 17960 3188
rect 17543 3148 17960 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 18506 3136 18512 3188
rect 18564 3176 18570 3188
rect 19797 3179 19855 3185
rect 19797 3176 19809 3179
rect 18564 3148 19809 3176
rect 18564 3136 18570 3148
rect 19797 3145 19809 3148
rect 19843 3145 19855 3179
rect 19797 3139 19855 3145
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 21085 3179 21143 3185
rect 21085 3176 21097 3179
rect 20864 3148 21097 3176
rect 20864 3136 20870 3148
rect 21085 3145 21097 3148
rect 21131 3145 21143 3179
rect 21085 3139 21143 3145
rect 22738 3136 22744 3188
rect 22796 3176 22802 3188
rect 23017 3179 23075 3185
rect 23017 3176 23029 3179
rect 22796 3148 23029 3176
rect 22796 3136 22802 3148
rect 23017 3145 23029 3148
rect 23063 3176 23075 3179
rect 23566 3176 23572 3188
rect 23063 3148 23572 3176
rect 23063 3145 23075 3148
rect 23017 3139 23075 3145
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 25406 3176 25412 3188
rect 25367 3148 25412 3176
rect 25406 3136 25412 3148
rect 25464 3136 25470 3188
rect 27157 3179 27215 3185
rect 27157 3145 27169 3179
rect 27203 3176 27215 3179
rect 28534 3176 28540 3188
rect 27203 3148 28540 3176
rect 27203 3145 27215 3148
rect 27157 3139 27215 3145
rect 28534 3136 28540 3148
rect 28592 3136 28598 3188
rect 30561 3179 30619 3185
rect 30561 3145 30573 3179
rect 30607 3176 30619 3179
rect 30650 3176 30656 3188
rect 30607 3148 30656 3176
rect 30607 3145 30619 3148
rect 30561 3139 30619 3145
rect 30650 3136 30656 3148
rect 30708 3136 30714 3188
rect 32214 3176 32220 3188
rect 32175 3148 32220 3176
rect 32214 3136 32220 3148
rect 32272 3136 32278 3188
rect 14056 3080 14688 3108
rect 14056 3068 14062 3080
rect 9306 3040 9312 3052
rect 8772 3012 9312 3040
rect 7834 2972 7840 2984
rect 7484 2944 7840 2972
rect 7834 2932 7840 2944
rect 7892 2972 7898 2984
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7892 2944 8033 2972
rect 7892 2932 7898 2944
rect 8021 2941 8033 2944
rect 8067 2972 8079 2975
rect 8202 2972 8208 2984
rect 8067 2944 8208 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 8772 2981 8800 3012
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 14737 3043 14795 3049
rect 12492 3012 12537 3040
rect 12492 3000 12498 3012
rect 14737 3009 14749 3043
rect 14783 3009 14795 3043
rect 14737 3003 14795 3009
rect 8757 2975 8815 2981
rect 8757 2972 8769 2975
rect 8628 2944 8769 2972
rect 8628 2932 8634 2944
rect 8757 2941 8769 2944
rect 8803 2941 8815 2975
rect 8757 2935 8815 2941
rect 9033 2975 9091 2981
rect 9033 2941 9045 2975
rect 9079 2972 9091 2975
rect 9122 2972 9128 2984
rect 9079 2944 9128 2972
rect 9079 2941 9091 2944
rect 9033 2935 9091 2941
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9582 2972 9588 2984
rect 9263 2944 9588 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 8110 2864 8116 2916
rect 8168 2904 8174 2916
rect 9232 2904 9260 2935
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 11149 2975 11207 2981
rect 11149 2972 11161 2975
rect 11112 2944 11161 2972
rect 11112 2932 11118 2944
rect 11149 2941 11161 2944
rect 11195 2941 11207 2975
rect 12250 2972 12256 2984
rect 12163 2944 12256 2972
rect 11149 2935 11207 2941
rect 12250 2932 12256 2944
rect 12308 2972 12314 2984
rect 12529 2975 12587 2981
rect 12529 2972 12541 2975
rect 12308 2944 12541 2972
rect 12308 2932 12314 2944
rect 12529 2941 12541 2944
rect 12575 2941 12587 2975
rect 12529 2935 12587 2941
rect 13722 2932 13728 2984
rect 13780 2972 13786 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 13780 2944 14289 2972
rect 13780 2932 13786 2944
rect 14277 2941 14289 2944
rect 14323 2972 14335 2975
rect 14752 2972 14780 3003
rect 15378 3000 15384 3052
rect 15436 3040 15442 3052
rect 15933 3043 15991 3049
rect 15933 3040 15945 3043
rect 15436 3012 15945 3040
rect 15436 3000 15442 3012
rect 15933 3009 15945 3012
rect 15979 3009 15991 3043
rect 17972 3040 18000 3136
rect 22646 3108 22652 3120
rect 22607 3080 22652 3108
rect 22646 3068 22652 3080
rect 22704 3068 22710 3120
rect 24854 3068 24860 3120
rect 24912 3108 24918 3120
rect 26053 3111 26111 3117
rect 26053 3108 26065 3111
rect 24912 3080 26065 3108
rect 24912 3068 24918 3080
rect 26053 3077 26065 3080
rect 26099 3108 26111 3111
rect 26326 3108 26332 3120
rect 26099 3080 26332 3108
rect 26099 3077 26111 3080
rect 26053 3071 26111 3077
rect 26326 3068 26332 3080
rect 26384 3068 26390 3120
rect 32232 3080 32812 3108
rect 17972 3012 18552 3040
rect 15933 3003 15991 3009
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 14323 2944 15853 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 15841 2941 15853 2944
rect 15887 2972 15899 2975
rect 16298 2972 16304 2984
rect 15887 2944 16304 2972
rect 15887 2941 15899 2944
rect 15841 2935 15899 2941
rect 16298 2932 16304 2944
rect 16356 2972 16362 2984
rect 16574 2972 16580 2984
rect 16356 2944 16580 2972
rect 16356 2932 16362 2944
rect 16574 2932 16580 2944
rect 16632 2932 16638 2984
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 18524 2981 18552 3012
rect 22370 3000 22376 3052
rect 22428 3040 22434 3052
rect 23477 3043 23535 3049
rect 23477 3040 23489 3043
rect 22428 3012 23489 3040
rect 22428 3000 22434 3012
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17460 2944 18061 2972
rect 17460 2932 17466 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2941 18567 2975
rect 18874 2972 18880 2984
rect 18835 2944 18880 2972
rect 18509 2935 18567 2941
rect 18874 2932 18880 2944
rect 18932 2932 18938 2984
rect 19242 2972 19248 2984
rect 19203 2944 19248 2972
rect 19242 2932 19248 2944
rect 19300 2972 19306 2984
rect 20165 2975 20223 2981
rect 20165 2972 20177 2975
rect 19300 2944 20177 2972
rect 19300 2932 19306 2944
rect 20165 2941 20177 2944
rect 20211 2972 20223 2975
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 20211 2944 20545 2972
rect 20211 2941 20223 2944
rect 20165 2935 20223 2941
rect 20533 2941 20545 2944
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 21545 2975 21603 2981
rect 21545 2941 21557 2975
rect 21591 2972 21603 2975
rect 21634 2972 21640 2984
rect 21591 2944 21640 2972
rect 21591 2941 21603 2944
rect 21545 2935 21603 2941
rect 21634 2932 21640 2944
rect 21692 2932 21698 2984
rect 21910 2972 21916 2984
rect 21871 2944 21916 2972
rect 21910 2932 21916 2944
rect 21968 2972 21974 2984
rect 22094 2972 22100 2984
rect 21968 2944 22100 2972
rect 21968 2932 21974 2944
rect 22094 2932 22100 2944
rect 22152 2932 22158 2984
rect 22281 2975 22339 2981
rect 22281 2941 22293 2975
rect 22327 2972 22339 2975
rect 22462 2972 22468 2984
rect 22327 2944 22468 2972
rect 22327 2941 22339 2944
rect 22281 2935 22339 2941
rect 22462 2932 22468 2944
rect 22520 2932 22526 2984
rect 22664 2981 22692 3012
rect 23477 3009 23489 3012
rect 23523 3040 23535 3043
rect 23750 3040 23756 3052
rect 23523 3012 23756 3040
rect 23523 3009 23535 3012
rect 23477 3003 23535 3009
rect 23750 3000 23756 3012
rect 23808 3040 23814 3052
rect 26234 3040 26240 3052
rect 23808 3012 24900 3040
rect 26195 3012 26240 3040
rect 23808 3000 23814 3012
rect 22649 2975 22707 2981
rect 22649 2941 22661 2975
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 23661 2975 23719 2981
rect 23661 2941 23673 2975
rect 23707 2941 23719 2975
rect 24118 2972 24124 2984
rect 24079 2944 24124 2972
rect 23661 2935 23719 2941
rect 8168 2876 9260 2904
rect 10873 2907 10931 2913
rect 8168 2864 8174 2876
rect 10873 2873 10885 2907
rect 10919 2904 10931 2907
rect 10962 2904 10968 2916
rect 10919 2876 10968 2904
rect 10919 2873 10931 2876
rect 10873 2867 10931 2873
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 11790 2864 11796 2916
rect 11848 2904 11854 2916
rect 11885 2907 11943 2913
rect 11885 2904 11897 2907
rect 11848 2876 11897 2904
rect 11848 2864 11854 2876
rect 11885 2873 11897 2876
rect 11931 2904 11943 2907
rect 12618 2904 12624 2916
rect 11931 2876 12624 2904
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 12618 2864 12624 2876
rect 12676 2864 12682 2916
rect 14369 2907 14427 2913
rect 14369 2873 14381 2907
rect 14415 2904 14427 2907
rect 14918 2904 14924 2916
rect 14415 2876 14924 2904
rect 14415 2873 14427 2876
rect 14369 2867 14427 2873
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 15102 2904 15108 2916
rect 15063 2876 15108 2904
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 18892 2904 18920 2932
rect 19518 2904 19524 2916
rect 18892 2876 19524 2904
rect 19518 2864 19524 2876
rect 19576 2864 19582 2916
rect 20714 2864 20720 2916
rect 20772 2904 20778 2916
rect 22370 2904 22376 2916
rect 20772 2876 22376 2904
rect 20772 2864 20778 2876
rect 22370 2864 22376 2876
rect 22428 2904 22434 2916
rect 22554 2904 22560 2916
rect 22428 2876 22560 2904
rect 22428 2864 22434 2876
rect 22554 2864 22560 2876
rect 22612 2864 22618 2916
rect 23474 2864 23480 2916
rect 23532 2904 23538 2916
rect 23676 2904 23704 2935
rect 24118 2932 24124 2944
rect 24176 2932 24182 2984
rect 24578 2972 24584 2984
rect 24539 2944 24584 2972
rect 24578 2932 24584 2944
rect 24636 2932 24642 2984
rect 24872 2981 24900 3012
rect 26234 3000 26240 3012
rect 26292 3000 26298 3052
rect 29270 3040 29276 3052
rect 29231 3012 29276 3040
rect 29270 3000 29276 3012
rect 29328 3000 29334 3052
rect 30929 3043 30987 3049
rect 30929 3009 30941 3043
rect 30975 3040 30987 3043
rect 31294 3040 31300 3052
rect 30975 3012 31300 3040
rect 30975 3009 30987 3012
rect 30929 3003 30987 3009
rect 31294 3000 31300 3012
rect 31352 3000 31358 3052
rect 31573 3043 31631 3049
rect 31573 3009 31585 3043
rect 31619 3040 31631 3043
rect 32030 3040 32036 3052
rect 31619 3012 32036 3040
rect 31619 3009 31631 3012
rect 31573 3003 31631 3009
rect 32030 3000 32036 3012
rect 32088 3040 32094 3052
rect 32232 3040 32260 3080
rect 32490 3040 32496 3052
rect 32088 3012 32260 3040
rect 32324 3012 32496 3040
rect 32088 3000 32094 3012
rect 24857 2975 24915 2981
rect 24857 2941 24869 2975
rect 24903 2941 24915 2975
rect 24857 2935 24915 2941
rect 25133 2975 25191 2981
rect 25133 2941 25145 2975
rect 25179 2972 25191 2975
rect 26418 2972 26424 2984
rect 25179 2944 26424 2972
rect 25179 2941 25191 2944
rect 25133 2935 25191 2941
rect 26418 2932 26424 2944
rect 26476 2972 26482 2984
rect 27801 2975 27859 2981
rect 27801 2972 27813 2975
rect 26476 2944 27813 2972
rect 26476 2932 26482 2944
rect 27801 2941 27813 2944
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 28077 2975 28135 2981
rect 28077 2941 28089 2975
rect 28123 2972 28135 2975
rect 28994 2972 29000 2984
rect 28123 2944 29000 2972
rect 28123 2941 28135 2944
rect 28077 2935 28135 2941
rect 28994 2932 29000 2944
rect 29052 2932 29058 2984
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 29365 2975 29423 2981
rect 29365 2972 29377 2975
rect 29144 2944 29377 2972
rect 29144 2932 29150 2944
rect 29365 2941 29377 2944
rect 29411 2941 29423 2975
rect 29365 2935 29423 2941
rect 23532 2876 23704 2904
rect 23532 2864 23538 2876
rect 26326 2864 26332 2916
rect 26384 2904 26390 2916
rect 26558 2907 26616 2913
rect 26558 2904 26570 2907
rect 26384 2876 26570 2904
rect 26384 2864 26390 2876
rect 26558 2873 26570 2876
rect 26604 2873 26616 2907
rect 26558 2867 26616 2873
rect 30926 2864 30932 2916
rect 30984 2904 30990 2916
rect 31021 2907 31079 2913
rect 31021 2904 31033 2907
rect 30984 2876 31033 2904
rect 30984 2864 30990 2876
rect 31021 2873 31033 2876
rect 31067 2873 31079 2907
rect 31021 2867 31079 2873
rect 31202 2864 31208 2916
rect 31260 2904 31266 2916
rect 32324 2904 32352 3012
rect 32490 3000 32496 3012
rect 32548 3000 32554 3052
rect 32784 3049 32812 3080
rect 32769 3043 32827 3049
rect 32769 3009 32781 3043
rect 32815 3009 32827 3043
rect 32769 3003 32827 3009
rect 32582 2904 32588 2916
rect 31260 2876 32352 2904
rect 32495 2876 32588 2904
rect 31260 2864 31266 2876
rect 32582 2864 32588 2876
rect 32640 2904 32646 2916
rect 33413 2907 33471 2913
rect 33413 2904 33425 2907
rect 32640 2876 33425 2904
rect 32640 2864 32646 2876
rect 33413 2873 33425 2876
rect 33459 2873 33471 2907
rect 33413 2867 33471 2873
rect 5169 2839 5227 2845
rect 5169 2805 5181 2839
rect 5215 2836 5227 2839
rect 5258 2836 5264 2848
rect 5215 2808 5264 2836
rect 5215 2805 5227 2808
rect 5169 2799 5227 2805
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 5534 2836 5540 2848
rect 5408 2808 5540 2836
rect 5408 2796 5414 2808
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 7926 2836 7932 2848
rect 7887 2808 7932 2836
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 8294 2836 8300 2848
rect 8255 2808 8300 2836
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 18322 2836 18328 2848
rect 18235 2808 18328 2836
rect 18322 2796 18328 2808
rect 18380 2836 18386 2848
rect 18690 2836 18696 2848
rect 18380 2808 18696 2836
rect 18380 2796 18386 2808
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 27430 2836 27436 2848
rect 27391 2808 27436 2836
rect 27430 2796 27436 2808
rect 27488 2796 27494 2848
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 3016 2604 3065 2632
rect 3016 2592 3022 2604
rect 3053 2601 3065 2604
rect 3099 2601 3111 2635
rect 3053 2595 3111 2601
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 3421 2635 3479 2641
rect 3421 2632 3433 2635
rect 3292 2604 3433 2632
rect 3292 2592 3298 2604
rect 3421 2601 3433 2604
rect 3467 2601 3479 2635
rect 7834 2632 7840 2644
rect 7795 2604 7840 2632
rect 3421 2595 3479 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8570 2632 8576 2644
rect 8531 2604 8576 2632
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 8846 2632 8852 2644
rect 8807 2604 8852 2632
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12802 2632 12808 2644
rect 12492 2604 12537 2632
rect 12763 2604 12808 2632
rect 12492 2592 12498 2604
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 13722 2632 13728 2644
rect 13683 2604 13728 2632
rect 13722 2592 13728 2604
rect 13780 2632 13786 2644
rect 13906 2632 13912 2644
rect 13780 2604 13912 2632
rect 13780 2592 13786 2604
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 14918 2632 14924 2644
rect 14879 2604 14924 2632
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 15654 2592 15660 2644
rect 15712 2632 15718 2644
rect 16301 2635 16359 2641
rect 16301 2632 16313 2635
rect 15712 2604 16313 2632
rect 15712 2592 15718 2604
rect 16301 2601 16313 2604
rect 16347 2601 16359 2635
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 16301 2595 16359 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 20254 2641 20260 2644
rect 19889 2635 19947 2641
rect 19889 2632 19901 2635
rect 19392 2604 19901 2632
rect 19392 2592 19398 2604
rect 19889 2601 19901 2604
rect 19935 2601 19947 2635
rect 19889 2595 19947 2601
rect 20211 2635 20260 2641
rect 20211 2601 20223 2635
rect 20257 2601 20260 2635
rect 20211 2595 20260 2601
rect 20254 2592 20260 2595
rect 20312 2592 20318 2644
rect 20622 2632 20628 2644
rect 20583 2604 20628 2632
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 28994 2592 29000 2644
rect 29052 2632 29058 2644
rect 29089 2635 29147 2641
rect 29089 2632 29101 2635
rect 29052 2604 29101 2632
rect 29052 2592 29058 2604
rect 29089 2601 29101 2604
rect 29135 2601 29147 2635
rect 29546 2632 29552 2644
rect 29507 2604 29552 2632
rect 29089 2595 29147 2601
rect 2777 2567 2835 2573
rect 2777 2533 2789 2567
rect 2823 2564 2835 2567
rect 3510 2564 3516 2576
rect 2823 2536 3516 2564
rect 2823 2533 2835 2536
rect 2777 2527 2835 2533
rect 3510 2524 3516 2536
rect 3568 2564 3574 2576
rect 5261 2567 5319 2573
rect 5261 2564 5273 2567
rect 3568 2536 5273 2564
rect 3568 2524 3574 2536
rect 5261 2533 5273 2536
rect 5307 2564 5319 2567
rect 5442 2564 5448 2576
rect 5307 2536 5448 2564
rect 5307 2533 5319 2536
rect 5261 2527 5319 2533
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 7561 2567 7619 2573
rect 7561 2533 7573 2567
rect 7607 2564 7619 2567
rect 8110 2564 8116 2576
rect 7607 2536 8116 2564
rect 7607 2533 7619 2536
rect 7561 2527 7619 2533
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 10962 2524 10968 2576
rect 11020 2564 11026 2576
rect 11422 2564 11428 2576
rect 11020 2536 11428 2564
rect 11020 2524 11026 2536
rect 11422 2524 11428 2536
rect 11480 2524 11486 2576
rect 1765 2499 1823 2505
rect 1765 2465 1777 2499
rect 1811 2496 1823 2499
rect 3234 2496 3240 2508
rect 1811 2468 3240 2496
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 3234 2456 3240 2468
rect 3292 2456 3298 2508
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 7926 2496 7932 2508
rect 7699 2468 7932 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 7926 2456 7932 2468
rect 7984 2496 7990 2508
rect 8662 2496 8668 2508
rect 7984 2468 8248 2496
rect 8623 2468 8668 2496
rect 7984 2456 7990 2468
rect 8220 2369 8248 2468
rect 8662 2456 8668 2468
rect 8720 2496 8726 2508
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8720 2468 9137 2496
rect 8720 2456 8726 2468
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 9125 2459 9183 2465
rect 10520 2468 10793 2496
rect 10520 2372 10548 2468
rect 10781 2465 10793 2468
rect 10827 2465 10839 2499
rect 12452 2496 12480 2592
rect 16850 2564 16856 2576
rect 16763 2536 16856 2564
rect 16850 2524 16856 2536
rect 16908 2564 16914 2576
rect 18156 2564 18184 2592
rect 18646 2567 18704 2573
rect 18646 2564 18658 2567
rect 16908 2536 17724 2564
rect 18156 2536 18658 2564
rect 16908 2524 16914 2536
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12452 2468 12633 2496
rect 10781 2459 10839 2465
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 13722 2456 13728 2508
rect 13780 2496 13786 2508
rect 13817 2499 13875 2505
rect 13817 2496 13829 2499
rect 13780 2468 13829 2496
rect 13780 2456 13786 2468
rect 13817 2465 13829 2468
rect 13863 2465 13875 2499
rect 13817 2459 13875 2465
rect 13906 2456 13912 2508
rect 13964 2505 13970 2508
rect 13964 2499 14022 2505
rect 13964 2465 13976 2499
rect 14010 2465 14022 2499
rect 13964 2459 14022 2465
rect 13964 2456 13970 2459
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15160 2468 15485 2496
rect 15160 2456 15166 2468
rect 15473 2465 15485 2468
rect 15519 2496 15531 2499
rect 15519 2468 16160 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 12066 2428 12072 2440
rect 12027 2400 12072 2428
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2428 13415 2431
rect 14182 2428 14188 2440
rect 13403 2400 14188 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 15286 2428 15292 2440
rect 15199 2400 15292 2428
rect 15286 2388 15292 2400
rect 15344 2428 15350 2440
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 15344 2400 15945 2428
rect 15344 2388 15350 2400
rect 15933 2397 15945 2400
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 8205 2363 8263 2369
rect 8205 2329 8217 2363
rect 8251 2360 8263 2363
rect 9030 2360 9036 2372
rect 8251 2332 9036 2360
rect 8251 2329 8263 2332
rect 8205 2323 8263 2329
rect 9030 2320 9036 2332
rect 9088 2320 9094 2372
rect 10502 2360 10508 2372
rect 10463 2332 10508 2360
rect 10502 2320 10508 2332
rect 10560 2320 10566 2372
rect 14093 2363 14151 2369
rect 14093 2329 14105 2363
rect 14139 2360 14151 2363
rect 14918 2360 14924 2372
rect 14139 2332 14924 2360
rect 14139 2329 14151 2332
rect 14093 2323 14151 2329
rect 14918 2320 14924 2332
rect 14976 2320 14982 2372
rect 15654 2360 15660 2372
rect 15615 2332 15660 2360
rect 15654 2320 15660 2332
rect 15712 2320 15718 2372
rect 16132 2360 16160 2468
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 17460 2468 17505 2496
rect 17460 2456 17466 2468
rect 16758 2428 16764 2440
rect 16719 2400 16764 2428
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 17696 2428 17724 2536
rect 18646 2533 18658 2536
rect 18692 2533 18704 2567
rect 19518 2564 19524 2576
rect 19479 2536 19524 2564
rect 18646 2527 18704 2533
rect 19518 2524 19524 2536
rect 19576 2564 19582 2576
rect 21453 2567 21511 2573
rect 21453 2564 21465 2567
rect 19576 2536 21465 2564
rect 19576 2524 19582 2536
rect 21453 2533 21465 2536
rect 21499 2564 21511 2567
rect 23106 2564 23112 2576
rect 21499 2536 21772 2564
rect 23067 2536 23112 2564
rect 21499 2533 21511 2536
rect 21453 2527 21511 2533
rect 18322 2496 18328 2508
rect 18283 2468 18328 2496
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 20070 2456 20076 2508
rect 20128 2505 20134 2508
rect 20128 2499 20166 2505
rect 20154 2496 20166 2499
rect 20530 2496 20536 2508
rect 20154 2468 20536 2496
rect 20154 2465 20166 2468
rect 20128 2459 20166 2465
rect 20128 2456 20134 2459
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 20993 2499 21051 2505
rect 20993 2465 21005 2499
rect 21039 2496 21051 2499
rect 21542 2496 21548 2508
rect 21039 2468 21548 2496
rect 21039 2465 21051 2468
rect 20993 2459 21051 2465
rect 21542 2456 21548 2468
rect 21600 2496 21606 2508
rect 21637 2499 21695 2505
rect 21637 2496 21649 2499
rect 21600 2468 21649 2496
rect 21600 2456 21606 2468
rect 21637 2465 21649 2468
rect 21683 2465 21695 2499
rect 21637 2459 21695 2465
rect 21744 2428 21772 2536
rect 23106 2524 23112 2536
rect 23164 2524 23170 2576
rect 23845 2567 23903 2573
rect 23845 2564 23857 2567
rect 23216 2536 23857 2564
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22152 2468 22197 2496
rect 22152 2456 22158 2468
rect 22370 2456 22376 2508
rect 22428 2496 22434 2508
rect 22465 2499 22523 2505
rect 22465 2496 22477 2499
rect 22428 2468 22477 2496
rect 22428 2456 22434 2468
rect 22465 2465 22477 2468
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 22922 2456 22928 2508
rect 22980 2496 22986 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22980 2468 23029 2496
rect 22980 2456 22986 2468
rect 23017 2465 23029 2468
rect 23063 2496 23075 2499
rect 23216 2496 23244 2536
rect 23845 2533 23857 2536
rect 23891 2564 23903 2567
rect 26237 2567 26295 2573
rect 23891 2536 25268 2564
rect 23891 2533 23903 2536
rect 23845 2527 23903 2533
rect 23474 2496 23480 2508
rect 23063 2468 23244 2496
rect 23387 2468 23480 2496
rect 23063 2465 23075 2468
rect 23017 2459 23075 2465
rect 23474 2456 23480 2468
rect 23532 2496 23538 2508
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 23532 2468 24041 2496
rect 23532 2456 23538 2468
rect 24029 2465 24041 2468
rect 24075 2465 24087 2499
rect 24029 2459 24087 2465
rect 24118 2456 24124 2508
rect 24176 2496 24182 2508
rect 24765 2499 24823 2505
rect 24765 2496 24777 2499
rect 24176 2468 24777 2496
rect 24176 2456 24182 2468
rect 24765 2465 24777 2468
rect 24811 2465 24823 2499
rect 25038 2496 25044 2508
rect 24999 2468 25044 2496
rect 24765 2459 24823 2465
rect 22940 2428 22968 2456
rect 17696 2400 19288 2428
rect 21744 2400 22968 2428
rect 24780 2428 24808 2459
rect 25038 2456 25044 2468
rect 25096 2456 25102 2508
rect 25240 2505 25268 2536
rect 26237 2533 26249 2567
rect 26283 2564 26295 2567
rect 26326 2564 26332 2576
rect 26283 2536 26332 2564
rect 26283 2533 26295 2536
rect 26237 2527 26295 2533
rect 26326 2524 26332 2536
rect 26384 2564 26390 2576
rect 26605 2567 26663 2573
rect 26605 2564 26617 2567
rect 26384 2536 26617 2564
rect 26384 2524 26390 2536
rect 26605 2533 26617 2536
rect 26651 2564 26663 2567
rect 27154 2564 27160 2576
rect 26651 2536 27160 2564
rect 26651 2533 26663 2536
rect 26605 2527 26663 2533
rect 27154 2524 27160 2536
rect 27212 2573 27218 2576
rect 27212 2567 27260 2573
rect 27212 2533 27214 2567
rect 27248 2533 27260 2567
rect 27212 2527 27260 2533
rect 27212 2524 27218 2527
rect 27614 2524 27620 2576
rect 27672 2564 27678 2576
rect 28445 2567 28503 2573
rect 28445 2564 28457 2567
rect 27672 2536 28457 2564
rect 27672 2524 27678 2536
rect 28445 2533 28457 2536
rect 28491 2533 28503 2567
rect 29104 2564 29132 2595
rect 29546 2592 29552 2604
rect 29604 2632 29610 2644
rect 30926 2632 30932 2644
rect 29604 2604 29960 2632
rect 30887 2604 30932 2632
rect 29604 2592 29610 2604
rect 29932 2573 29960 2604
rect 30926 2592 30932 2604
rect 30984 2592 30990 2644
rect 31294 2632 31300 2644
rect 31255 2604 31300 2632
rect 31294 2592 31300 2604
rect 31352 2592 31358 2644
rect 31662 2641 31668 2644
rect 31619 2635 31668 2641
rect 31619 2601 31631 2635
rect 31665 2601 31668 2635
rect 31619 2595 31668 2601
rect 31662 2592 31668 2595
rect 31720 2592 31726 2644
rect 32030 2632 32036 2644
rect 31991 2604 32036 2632
rect 32030 2592 32036 2604
rect 32088 2592 32094 2644
rect 29825 2567 29883 2573
rect 29825 2564 29837 2567
rect 29104 2536 29837 2564
rect 28445 2527 28503 2533
rect 29825 2533 29837 2536
rect 29871 2533 29883 2567
rect 29825 2527 29883 2533
rect 29917 2567 29975 2573
rect 29917 2533 29929 2567
rect 29963 2533 29975 2567
rect 29917 2527 29975 2533
rect 25225 2499 25283 2505
rect 25225 2465 25237 2499
rect 25271 2465 25283 2499
rect 25225 2459 25283 2465
rect 25501 2499 25559 2505
rect 25501 2465 25513 2499
rect 25547 2496 25559 2499
rect 26881 2499 26939 2505
rect 26881 2496 26893 2499
rect 25547 2468 26893 2496
rect 25547 2465 25559 2468
rect 25501 2459 25559 2465
rect 26881 2465 26893 2468
rect 26927 2496 26939 2499
rect 27430 2496 27436 2508
rect 26927 2468 27436 2496
rect 26927 2465 26939 2468
rect 26881 2459 26939 2465
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 27798 2496 27804 2508
rect 27759 2468 27804 2496
rect 27798 2456 27804 2468
rect 27856 2456 27862 2508
rect 28696 2499 28754 2505
rect 28696 2465 28708 2499
rect 28742 2496 28754 2499
rect 28902 2496 28908 2508
rect 28742 2468 28908 2496
rect 28742 2465 28754 2468
rect 28696 2459 28754 2465
rect 28902 2456 28908 2468
rect 28960 2456 28966 2508
rect 31548 2499 31606 2505
rect 31548 2465 31560 2499
rect 31594 2496 31606 2499
rect 32048 2496 32076 2592
rect 32582 2524 32588 2576
rect 32640 2524 32646 2576
rect 31594 2468 32076 2496
rect 32401 2499 32459 2505
rect 31594 2465 31606 2468
rect 31548 2459 31606 2465
rect 32401 2465 32413 2499
rect 32447 2496 32459 2499
rect 32600 2496 32628 2524
rect 32677 2499 32735 2505
rect 32677 2496 32689 2499
rect 32447 2468 32689 2496
rect 32447 2465 32459 2468
rect 32401 2459 32459 2465
rect 32677 2465 32689 2468
rect 32723 2465 32735 2499
rect 32677 2459 32735 2465
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 24780 2400 25881 2428
rect 19260 2369 19288 2400
rect 25869 2397 25881 2400
rect 25915 2428 25927 2431
rect 28077 2431 28135 2437
rect 28077 2428 28089 2431
rect 25915 2400 28089 2428
rect 25915 2397 25927 2400
rect 25869 2391 25927 2397
rect 28077 2397 28089 2400
rect 28123 2397 28135 2431
rect 28920 2428 28948 2456
rect 30101 2431 30159 2437
rect 30101 2428 30113 2431
rect 28920 2400 30113 2428
rect 28077 2391 28135 2397
rect 30101 2397 30113 2400
rect 30147 2397 30159 2431
rect 30101 2391 30159 2397
rect 30926 2388 30932 2440
rect 30984 2428 30990 2440
rect 32585 2431 32643 2437
rect 32585 2428 32597 2431
rect 30984 2400 32597 2428
rect 30984 2388 30990 2400
rect 32585 2397 32597 2400
rect 32631 2397 32643 2431
rect 32585 2391 32643 2397
rect 34149 2431 34207 2437
rect 34149 2397 34161 2431
rect 34195 2397 34207 2431
rect 34149 2391 34207 2397
rect 17681 2363 17739 2369
rect 17681 2360 17693 2363
rect 16132 2332 17693 2360
rect 17681 2329 17693 2332
rect 17727 2329 17739 2363
rect 17681 2323 17739 2329
rect 19245 2363 19303 2369
rect 19245 2329 19257 2363
rect 19291 2329 19303 2363
rect 19245 2323 19303 2329
rect 28767 2363 28825 2369
rect 28767 2329 28779 2363
rect 28813 2360 28825 2363
rect 28902 2360 28908 2372
rect 28813 2332 28908 2360
rect 28813 2329 28825 2332
rect 28767 2323 28825 2329
rect 28902 2320 28908 2332
rect 28960 2320 28966 2372
rect 31294 2320 31300 2372
rect 31352 2360 31358 2372
rect 34164 2360 34192 2391
rect 31352 2332 34192 2360
rect 31352 2320 31358 2332
rect 13814 2252 13820 2304
rect 13872 2292 13878 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13872 2264 14289 2292
rect 13872 2252 13878 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
rect 19334 8 19340 60
rect 19392 48 19398 60
rect 28902 48 28908 60
rect 19392 20 28908 48
rect 19392 8 19398 20
rect 28902 8 28908 20
rect 28960 8 28966 60
<< via1 >>
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 35624 11339 35676 11348
rect 35624 11305 35633 11339
rect 35633 11305 35667 11339
rect 35667 11305 35676 11339
rect 35624 11296 35676 11305
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 35440 11203 35492 11212
rect 35440 11169 35449 11203
rect 35449 11169 35483 11203
rect 35483 11169 35492 11203
rect 35440 11160 35492 11169
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 1400 10752 1452 10804
rect 2688 10752 2740 10804
rect 35440 10455 35492 10464
rect 35440 10421 35449 10455
rect 35449 10421 35483 10455
rect 35483 10421 35492 10455
rect 35440 10412 35492 10421
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 35624 10251 35676 10260
rect 35624 10217 35633 10251
rect 35633 10217 35667 10251
rect 35667 10217 35676 10251
rect 35624 10208 35676 10217
rect 1676 10072 1728 10124
rect 35440 10115 35492 10124
rect 35440 10081 35449 10115
rect 35449 10081 35483 10115
rect 35483 10081 35492 10115
rect 35440 10072 35492 10081
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 35440 9503 35492 9512
rect 35440 9469 35449 9503
rect 35449 9469 35483 9503
rect 35483 9469 35492 9503
rect 35440 9460 35492 9469
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 1492 9120 1544 9172
rect 35716 9120 35768 9172
rect 2044 8984 2096 9036
rect 2688 8984 2740 9036
rect 3424 8984 3476 9036
rect 35440 9027 35492 9036
rect 35440 8993 35449 9027
rect 35449 8993 35483 9027
rect 35483 8993 35492 9027
rect 35440 8984 35492 8993
rect 2688 8780 2740 8832
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 1768 8576 1820 8628
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 3424 8619 3476 8628
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 35440 8576 35492 8628
rect 35624 8619 35676 8628
rect 35624 8585 35633 8619
rect 35633 8585 35667 8619
rect 35667 8585 35676 8619
rect 35624 8576 35676 8585
rect 2596 8508 2648 8560
rect 5448 8508 5500 8560
rect 3976 8483 4028 8492
rect 2872 8372 2924 8424
rect 3056 8415 3108 8424
rect 3056 8381 3065 8415
rect 3065 8381 3099 8415
rect 3099 8381 3108 8415
rect 3056 8372 3108 8381
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 4068 8372 4120 8424
rect 35440 8415 35492 8424
rect 35440 8381 35449 8415
rect 35449 8381 35483 8415
rect 35483 8381 35492 8415
rect 35440 8372 35492 8381
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 2504 8032 2556 8084
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 6644 8032 6696 8084
rect 35532 8032 35584 8084
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 2044 7896 2096 7948
rect 2504 7939 2556 7948
rect 2504 7905 2513 7939
rect 2513 7905 2547 7939
rect 2547 7905 2556 7939
rect 2504 7896 2556 7905
rect 5908 7896 5960 7948
rect 9864 7939 9916 7948
rect 9864 7905 9908 7939
rect 9908 7905 9916 7939
rect 9864 7896 9916 7905
rect 14188 7939 14240 7948
rect 14188 7905 14232 7939
rect 14232 7905 14240 7939
rect 19156 7939 19208 7948
rect 14188 7896 14240 7905
rect 19156 7905 19165 7939
rect 19165 7905 19199 7939
rect 19199 7905 19208 7939
rect 19156 7896 19208 7905
rect 35440 7939 35492 7948
rect 35440 7905 35449 7939
rect 35449 7905 35483 7939
rect 35483 7905 35492 7939
rect 35440 7896 35492 7905
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 5172 7828 5224 7880
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 10324 7692 10376 7744
rect 14464 7692 14516 7744
rect 20444 7692 20496 7744
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 1860 7488 1912 7540
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 4160 7488 4212 7540
rect 2504 7420 2556 7472
rect 3700 7420 3752 7472
rect 3240 7352 3292 7404
rect 4252 7352 4304 7404
rect 5080 7420 5132 7472
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 1676 7284 1728 7336
rect 4436 7284 4488 7336
rect 3148 7259 3200 7268
rect 3148 7225 3157 7259
rect 3157 7225 3191 7259
rect 3191 7225 3200 7259
rect 3148 7216 3200 7225
rect 3240 7259 3292 7268
rect 3240 7225 3249 7259
rect 3249 7225 3283 7259
rect 3283 7225 3292 7259
rect 3240 7216 3292 7225
rect 3976 7148 4028 7200
rect 4160 7148 4212 7200
rect 13084 7284 13136 7336
rect 14372 7488 14424 7540
rect 16672 7488 16724 7540
rect 19156 7488 19208 7540
rect 19800 7488 19852 7540
rect 35440 7488 35492 7540
rect 35808 7488 35860 7540
rect 36728 7531 36780 7540
rect 36728 7497 36737 7531
rect 36737 7497 36771 7531
rect 36771 7497 36780 7531
rect 36728 7488 36780 7497
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 16672 7284 16724 7336
rect 19064 7327 19116 7336
rect 19064 7293 19108 7327
rect 19108 7293 19116 7327
rect 19892 7327 19944 7336
rect 19064 7284 19116 7293
rect 19892 7293 19901 7327
rect 19901 7293 19935 7327
rect 19935 7293 19944 7327
rect 19892 7284 19944 7293
rect 19984 7284 20036 7336
rect 21640 7327 21692 7336
rect 13728 7216 13780 7268
rect 14832 7216 14884 7268
rect 21640 7293 21649 7327
rect 21649 7293 21683 7327
rect 21683 7293 21692 7327
rect 21640 7284 21692 7293
rect 34980 7284 35032 7336
rect 36544 7327 36596 7336
rect 36544 7293 36553 7327
rect 36553 7293 36587 7327
rect 36587 7293 36596 7327
rect 36544 7284 36596 7293
rect 5908 7148 5960 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 10508 7148 10560 7200
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 14188 7148 14240 7200
rect 15016 7148 15068 7200
rect 23020 7216 23072 7268
rect 15568 7148 15620 7200
rect 18972 7191 19024 7200
rect 18972 7157 18981 7191
rect 18981 7157 19015 7191
rect 19015 7157 19024 7191
rect 18972 7148 19024 7157
rect 19248 7148 19300 7200
rect 20168 7148 20220 7200
rect 20904 7191 20956 7200
rect 20904 7157 20913 7191
rect 20913 7157 20947 7191
rect 20947 7157 20956 7191
rect 20904 7148 20956 7157
rect 21916 7148 21968 7200
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 9496 6944 9548 6996
rect 9680 6944 9732 6996
rect 4252 6919 4304 6928
rect 2412 6808 2464 6860
rect 4252 6885 4261 6919
rect 4261 6885 4295 6919
rect 4295 6885 4304 6919
rect 4252 6876 4304 6885
rect 5172 6876 5224 6928
rect 5816 6919 5868 6928
rect 5816 6885 5825 6919
rect 5825 6885 5859 6919
rect 5859 6885 5868 6919
rect 5816 6876 5868 6885
rect 10324 6919 10376 6928
rect 10324 6885 10333 6919
rect 10333 6885 10367 6919
rect 10367 6885 10376 6919
rect 10324 6876 10376 6885
rect 10416 6919 10468 6928
rect 10416 6885 10425 6919
rect 10425 6885 10459 6919
rect 10459 6885 10468 6919
rect 10416 6876 10468 6885
rect 15476 6919 15528 6928
rect 3884 6740 3936 6792
rect 4344 6740 4396 6792
rect 2780 6672 2832 6724
rect 4436 6672 4488 6724
rect 12992 6808 13044 6860
rect 15476 6885 15485 6919
rect 15485 6885 15519 6919
rect 15519 6885 15528 6919
rect 15476 6876 15528 6885
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6920 6740 6972 6792
rect 8760 6740 8812 6792
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 14096 6740 14148 6792
rect 16580 6808 16632 6860
rect 23388 6944 23440 6996
rect 18236 6851 18288 6860
rect 18236 6817 18280 6851
rect 18280 6817 18288 6851
rect 18236 6808 18288 6817
rect 19064 6808 19116 6860
rect 20720 6808 20772 6860
rect 23480 6808 23532 6860
rect 24492 6851 24544 6860
rect 24492 6817 24501 6851
rect 24501 6817 24535 6851
rect 24535 6817 24544 6851
rect 24492 6808 24544 6817
rect 35440 6851 35492 6860
rect 35440 6817 35449 6851
rect 35449 6817 35483 6851
rect 35483 6817 35492 6851
rect 35440 6808 35492 6817
rect 15384 6783 15436 6792
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 15568 6740 15620 6792
rect 18604 6740 18656 6792
rect 20812 6740 20864 6792
rect 2504 6604 2556 6656
rect 4068 6604 4120 6656
rect 10600 6604 10652 6656
rect 18972 6672 19024 6724
rect 19892 6715 19944 6724
rect 19892 6681 19901 6715
rect 19901 6681 19935 6715
rect 19935 6681 19944 6715
rect 19892 6672 19944 6681
rect 20904 6672 20956 6724
rect 21548 6715 21600 6724
rect 21548 6681 21557 6715
rect 21557 6681 21591 6715
rect 21591 6681 21600 6715
rect 21548 6672 21600 6681
rect 35256 6672 35308 6724
rect 11336 6647 11388 6656
rect 11336 6613 11345 6647
rect 11345 6613 11379 6647
rect 11379 6613 11388 6647
rect 11336 6604 11388 6613
rect 13636 6604 13688 6656
rect 14832 6604 14884 6656
rect 15108 6647 15160 6656
rect 15108 6613 15117 6647
rect 15117 6613 15151 6647
rect 15151 6613 15160 6647
rect 15108 6604 15160 6613
rect 17040 6647 17092 6656
rect 17040 6613 17049 6647
rect 17049 6613 17083 6647
rect 17083 6613 17092 6647
rect 17040 6604 17092 6613
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 19064 6647 19116 6656
rect 19064 6613 19073 6647
rect 19073 6613 19107 6647
rect 19107 6613 19116 6647
rect 19064 6604 19116 6613
rect 19340 6604 19392 6656
rect 20168 6604 20220 6656
rect 24584 6647 24636 6656
rect 24584 6613 24593 6647
rect 24593 6613 24627 6647
rect 24627 6613 24636 6647
rect 24584 6604 24636 6613
rect 24860 6604 24912 6656
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 1952 6400 2004 6452
rect 3240 6400 3292 6452
rect 4068 6443 4120 6452
rect 4068 6409 4077 6443
rect 4077 6409 4111 6443
rect 4111 6409 4120 6443
rect 4068 6400 4120 6409
rect 5724 6400 5776 6452
rect 8760 6443 8812 6452
rect 8760 6409 8769 6443
rect 8769 6409 8803 6443
rect 8803 6409 8812 6443
rect 8760 6400 8812 6409
rect 10416 6400 10468 6452
rect 12992 6443 13044 6452
rect 12992 6409 13001 6443
rect 13001 6409 13035 6443
rect 13035 6409 13044 6443
rect 12992 6400 13044 6409
rect 15476 6400 15528 6452
rect 18236 6443 18288 6452
rect 18236 6409 18245 6443
rect 18245 6409 18279 6443
rect 18279 6409 18288 6443
rect 18236 6400 18288 6409
rect 18604 6400 18656 6452
rect 21272 6400 21324 6452
rect 2412 6375 2464 6384
rect 2412 6341 2421 6375
rect 2421 6341 2455 6375
rect 2455 6341 2464 6375
rect 2412 6332 2464 6341
rect 4252 6332 4304 6384
rect 5816 6332 5868 6384
rect 2780 6264 2832 6316
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 4436 6264 4488 6316
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 11152 6375 11204 6384
rect 11152 6341 11161 6375
rect 11161 6341 11195 6375
rect 11195 6341 11204 6375
rect 11152 6332 11204 6341
rect 14004 6332 14056 6384
rect 21548 6332 21600 6384
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 15108 6264 15160 6316
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 18972 6264 19024 6316
rect 20812 6264 20864 6316
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 13636 6239 13688 6248
rect 12440 6196 12492 6205
rect 13636 6205 13645 6239
rect 13645 6205 13679 6239
rect 13679 6205 13688 6239
rect 13636 6196 13688 6205
rect 18420 6239 18472 6248
rect 18420 6205 18464 6239
rect 18464 6205 18472 6239
rect 18880 6239 18932 6248
rect 18420 6196 18472 6205
rect 18880 6205 18889 6239
rect 18889 6205 18923 6239
rect 18923 6205 18932 6239
rect 18880 6196 18932 6205
rect 23296 6400 23348 6452
rect 24492 6443 24544 6452
rect 24492 6409 24501 6443
rect 24501 6409 24535 6443
rect 24535 6409 24544 6443
rect 24492 6400 24544 6409
rect 24676 6400 24728 6452
rect 25228 6332 25280 6384
rect 35440 6375 35492 6384
rect 35440 6341 35449 6375
rect 35449 6341 35483 6375
rect 35483 6341 35492 6375
rect 35440 6332 35492 6341
rect 24860 6264 24912 6316
rect 25412 6307 25464 6316
rect 25412 6273 25421 6307
rect 25421 6273 25455 6307
rect 25455 6273 25464 6307
rect 25412 6264 25464 6273
rect 2320 6128 2372 6180
rect 4344 6128 4396 6180
rect 9128 6171 9180 6180
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 4068 6060 4120 6112
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 9128 6137 9137 6171
rect 9137 6137 9171 6171
rect 9171 6137 9180 6171
rect 9128 6128 9180 6137
rect 9680 6128 9732 6180
rect 13544 6171 13596 6180
rect 13544 6137 13553 6171
rect 13553 6137 13587 6171
rect 13587 6137 13596 6171
rect 13544 6128 13596 6137
rect 14648 6128 14700 6180
rect 14832 6128 14884 6180
rect 15660 6128 15712 6180
rect 12624 6103 12676 6112
rect 6552 6060 6604 6069
rect 12624 6069 12633 6103
rect 12633 6069 12667 6103
rect 12667 6069 12676 6103
rect 12624 6060 12676 6069
rect 14740 6060 14792 6112
rect 15384 6060 15436 6112
rect 16580 6060 16632 6112
rect 17868 6103 17920 6112
rect 17868 6069 17877 6103
rect 17877 6069 17911 6103
rect 17911 6069 17920 6103
rect 17868 6060 17920 6069
rect 18972 6060 19024 6112
rect 19708 6128 19760 6180
rect 21088 6171 21140 6180
rect 20720 6060 20772 6112
rect 21088 6137 21097 6171
rect 21097 6137 21131 6171
rect 21131 6137 21140 6171
rect 21088 6128 21140 6137
rect 23480 6171 23532 6180
rect 23480 6137 23489 6171
rect 23489 6137 23523 6171
rect 23523 6137 23532 6171
rect 25228 6171 25280 6180
rect 23480 6128 23532 6137
rect 25228 6137 25237 6171
rect 25237 6137 25271 6171
rect 25271 6137 25280 6171
rect 25228 6128 25280 6137
rect 22744 6060 22796 6112
rect 24032 6103 24084 6112
rect 24032 6069 24041 6103
rect 24041 6069 24075 6103
rect 24075 6069 24084 6103
rect 24032 6060 24084 6069
rect 25044 6060 25096 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 2412 5788 2464 5840
rect 3884 5831 3936 5840
rect 3884 5797 3893 5831
rect 3893 5797 3927 5831
rect 3927 5797 3936 5831
rect 3884 5788 3936 5797
rect 4344 5788 4396 5840
rect 6276 5831 6328 5840
rect 6276 5797 6279 5831
rect 6279 5797 6313 5831
rect 6313 5797 6328 5831
rect 6276 5788 6328 5797
rect 9128 5856 9180 5908
rect 10324 5899 10376 5908
rect 10324 5865 10333 5899
rect 10333 5865 10367 5899
rect 10367 5865 10376 5899
rect 10324 5856 10376 5865
rect 14096 5856 14148 5908
rect 7472 5788 7524 5840
rect 10416 5788 10468 5840
rect 12532 5788 12584 5840
rect 12900 5788 12952 5840
rect 13544 5788 13596 5840
rect 14740 5788 14792 5840
rect 17776 5788 17828 5840
rect 19340 5831 19392 5840
rect 19340 5797 19349 5831
rect 19349 5797 19383 5831
rect 19383 5797 19392 5831
rect 19340 5788 19392 5797
rect 19708 5788 19760 5840
rect 21272 5831 21324 5840
rect 21272 5797 21275 5831
rect 21275 5797 21309 5831
rect 21309 5797 21324 5831
rect 21272 5788 21324 5797
rect 22744 5831 22796 5840
rect 22744 5797 22753 5831
rect 22753 5797 22787 5831
rect 22787 5797 22796 5831
rect 22744 5788 22796 5797
rect 22836 5831 22888 5840
rect 22836 5797 22845 5831
rect 22845 5797 22879 5831
rect 22879 5797 22888 5831
rect 24584 5831 24636 5840
rect 22836 5788 22888 5797
rect 24584 5797 24593 5831
rect 24593 5797 24627 5831
rect 24627 5797 24636 5831
rect 24584 5788 24636 5797
rect 4252 5720 4304 5772
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 6644 5652 6696 5704
rect 7380 5652 7432 5704
rect 2596 5584 2648 5636
rect 2688 5584 2740 5636
rect 3884 5584 3936 5636
rect 7196 5584 7248 5636
rect 10508 5652 10560 5704
rect 11060 5652 11112 5704
rect 13544 5652 13596 5704
rect 17040 5720 17092 5772
rect 25228 5720 25280 5772
rect 27252 5720 27304 5772
rect 15568 5652 15620 5704
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 16672 5652 16724 5704
rect 12624 5584 12676 5636
rect 13268 5584 13320 5636
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 3608 5516 3660 5568
rect 4988 5559 5040 5568
rect 4988 5525 4997 5559
rect 4997 5525 5031 5559
rect 5031 5525 5040 5559
rect 4988 5516 5040 5525
rect 8208 5516 8260 5568
rect 14924 5516 14976 5568
rect 16856 5516 16908 5568
rect 21364 5652 21416 5704
rect 19892 5627 19944 5636
rect 19892 5593 19901 5627
rect 19901 5593 19935 5627
rect 19935 5593 19944 5627
rect 19892 5584 19944 5593
rect 20628 5584 20680 5636
rect 24032 5652 24084 5704
rect 24492 5695 24544 5704
rect 24492 5661 24501 5695
rect 24501 5661 24535 5695
rect 24535 5661 24544 5695
rect 24492 5652 24544 5661
rect 26148 5652 26200 5704
rect 27988 5652 28040 5704
rect 25044 5627 25096 5636
rect 25044 5593 25053 5627
rect 25053 5593 25087 5627
rect 25087 5593 25096 5627
rect 25044 5584 25096 5593
rect 17868 5516 17920 5568
rect 20352 5559 20404 5568
rect 20352 5525 20361 5559
rect 20361 5525 20395 5559
rect 20395 5525 20404 5559
rect 20352 5516 20404 5525
rect 21824 5559 21876 5568
rect 21824 5525 21833 5559
rect 21833 5525 21867 5559
rect 21867 5525 21876 5559
rect 21824 5516 21876 5525
rect 22100 5559 22152 5568
rect 22100 5525 22109 5559
rect 22109 5525 22143 5559
rect 22143 5525 22152 5559
rect 22100 5516 22152 5525
rect 23388 5516 23440 5568
rect 24952 5516 25004 5568
rect 25412 5559 25464 5568
rect 25412 5525 25421 5559
rect 25421 5525 25455 5559
rect 25455 5525 25464 5559
rect 25412 5516 25464 5525
rect 27620 5516 27672 5568
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 1400 5312 1452 5364
rect 2412 5355 2464 5364
rect 2412 5321 2421 5355
rect 2421 5321 2455 5355
rect 2455 5321 2464 5355
rect 2412 5312 2464 5321
rect 6552 5312 6604 5364
rect 7380 5355 7432 5364
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 2596 5176 2648 5228
rect 7380 5321 7389 5355
rect 7389 5321 7423 5355
rect 7423 5321 7432 5355
rect 7380 5312 7432 5321
rect 9128 5312 9180 5364
rect 10416 5312 10468 5364
rect 11060 5312 11112 5364
rect 12900 5312 12952 5364
rect 15660 5355 15712 5364
rect 15660 5321 15669 5355
rect 15669 5321 15703 5355
rect 15703 5321 15712 5355
rect 15660 5312 15712 5321
rect 15752 5312 15804 5364
rect 17040 5312 17092 5364
rect 18972 5355 19024 5364
rect 18972 5321 18981 5355
rect 18981 5321 19015 5355
rect 19015 5321 19024 5355
rect 18972 5312 19024 5321
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 20720 5312 20772 5321
rect 22836 5312 22888 5364
rect 24216 5355 24268 5364
rect 24216 5321 24225 5355
rect 24225 5321 24259 5355
rect 24259 5321 24268 5355
rect 24216 5312 24268 5321
rect 24584 5355 24636 5364
rect 24584 5321 24593 5355
rect 24593 5321 24627 5355
rect 24627 5321 24636 5355
rect 24584 5312 24636 5321
rect 27252 5355 27304 5364
rect 27252 5321 27261 5355
rect 27261 5321 27295 5355
rect 27295 5321 27304 5355
rect 27252 5312 27304 5321
rect 35072 5312 35124 5364
rect 8208 5176 8260 5228
rect 2136 5108 2188 5160
rect 3516 5151 3568 5160
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 3792 5151 3844 5160
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 5080 5108 5132 5160
rect 9588 5151 9640 5160
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 3608 5040 3660 5092
rect 4344 5083 4396 5092
rect 4344 5049 4353 5083
rect 4353 5049 4387 5083
rect 4387 5049 4396 5083
rect 4344 5040 4396 5049
rect 6276 5083 6328 5092
rect 6276 5049 6285 5083
rect 6285 5049 6319 5083
rect 6319 5049 6328 5083
rect 6276 5040 6328 5049
rect 8208 5083 8260 5092
rect 8208 5049 8211 5083
rect 8211 5049 8245 5083
rect 8245 5049 8260 5083
rect 21548 5244 21600 5296
rect 24768 5244 24820 5296
rect 10140 5176 10192 5228
rect 12532 5151 12584 5160
rect 8208 5040 8260 5049
rect 12532 5117 12541 5151
rect 12541 5117 12575 5151
rect 12575 5117 12584 5151
rect 12532 5108 12584 5117
rect 22284 5219 22336 5228
rect 22284 5185 22293 5219
rect 22293 5185 22327 5219
rect 22327 5185 22336 5219
rect 22284 5176 22336 5185
rect 23388 5176 23440 5228
rect 25044 5219 25096 5228
rect 25044 5185 25053 5219
rect 25053 5185 25087 5219
rect 25087 5185 25096 5219
rect 25044 5176 25096 5185
rect 27528 5219 27580 5228
rect 27528 5185 27537 5219
rect 27537 5185 27571 5219
rect 27571 5185 27580 5219
rect 27528 5176 27580 5185
rect 13268 5151 13320 5160
rect 13268 5117 13277 5151
rect 13277 5117 13311 5151
rect 13311 5117 13320 5151
rect 13268 5108 13320 5117
rect 13728 5151 13780 5160
rect 13728 5117 13737 5151
rect 13737 5117 13771 5151
rect 13771 5117 13780 5151
rect 13728 5108 13780 5117
rect 13912 5108 13964 5160
rect 14924 5108 14976 5160
rect 16580 5108 16632 5160
rect 17960 5108 18012 5160
rect 19800 5151 19852 5160
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 24216 5108 24268 5160
rect 26332 5108 26384 5160
rect 26884 5151 26936 5160
rect 26884 5117 26893 5151
rect 26893 5117 26927 5151
rect 26927 5117 26936 5151
rect 26884 5108 26936 5117
rect 29000 5108 29052 5160
rect 14648 5083 14700 5092
rect 14648 5049 14657 5083
rect 14657 5049 14691 5083
rect 14691 5049 14700 5083
rect 15108 5083 15160 5092
rect 14648 5040 14700 5049
rect 15108 5049 15111 5083
rect 15111 5049 15145 5083
rect 15145 5049 15160 5083
rect 15108 5040 15160 5049
rect 15292 5040 15344 5092
rect 17040 5083 17092 5092
rect 17040 5049 17049 5083
rect 17049 5049 17083 5083
rect 17083 5049 17092 5083
rect 17040 5040 17092 5049
rect 17776 5040 17828 5092
rect 18144 5040 18196 5092
rect 21272 5040 21324 5092
rect 21732 5083 21784 5092
rect 21732 5049 21741 5083
rect 21741 5049 21775 5083
rect 21775 5049 21784 5083
rect 21732 5040 21784 5049
rect 22008 5040 22060 5092
rect 24768 5083 24820 5092
rect 24768 5049 24777 5083
rect 24777 5049 24811 5083
rect 24811 5049 24820 5083
rect 24768 5040 24820 5049
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 6644 5015 6696 5024
rect 2780 4972 2832 4981
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 19340 5015 19392 5024
rect 19340 4981 19349 5015
rect 19349 4981 19383 5015
rect 19383 4981 19392 5015
rect 19340 4972 19392 4981
rect 20904 4972 20956 5024
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 23296 4972 23348 5024
rect 23480 5015 23532 5024
rect 23480 4981 23489 5015
rect 23489 4981 23523 5015
rect 23523 4981 23532 5015
rect 23480 4972 23532 4981
rect 24676 4972 24728 5024
rect 27988 5040 28040 5092
rect 28264 5040 28316 5092
rect 26792 4972 26844 5024
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 2228 4768 2280 4820
rect 3976 4768 4028 4820
rect 5080 4811 5132 4820
rect 5080 4777 5089 4811
rect 5089 4777 5123 4811
rect 5123 4777 5132 4811
rect 5080 4768 5132 4777
rect 7472 4768 7524 4820
rect 9496 4768 9548 4820
rect 9588 4768 9640 4820
rect 15752 4768 15804 4820
rect 18144 4768 18196 4820
rect 21272 4768 21324 4820
rect 21824 4768 21876 4820
rect 23480 4811 23532 4820
rect 23480 4777 23489 4811
rect 23489 4777 23523 4811
rect 23523 4777 23532 4811
rect 23480 4768 23532 4777
rect 24492 4811 24544 4820
rect 24492 4777 24501 4811
rect 24501 4777 24535 4811
rect 24535 4777 24544 4811
rect 24492 4768 24544 4777
rect 25228 4768 25280 4820
rect 27528 4768 27580 4820
rect 2136 4700 2188 4752
rect 8208 4743 8260 4752
rect 8208 4709 8211 4743
rect 8211 4709 8245 4743
rect 8245 4709 8260 4743
rect 8208 4700 8260 4709
rect 13912 4743 13964 4752
rect 13912 4709 13921 4743
rect 13921 4709 13955 4743
rect 13955 4709 13964 4743
rect 13912 4700 13964 4709
rect 16028 4700 16080 4752
rect 1768 4675 1820 4684
rect 1768 4641 1777 4675
rect 1777 4641 1811 4675
rect 1811 4641 1820 4675
rect 1768 4632 1820 4641
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 2688 4632 2740 4641
rect 2964 4564 3016 4616
rect 3700 4632 3752 4684
rect 4252 4632 4304 4684
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 5908 4675 5960 4684
rect 5908 4641 5917 4675
rect 5917 4641 5951 4675
rect 5951 4641 5960 4675
rect 5908 4632 5960 4641
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 10140 4675 10192 4684
rect 6460 4564 6512 4616
rect 8024 4564 8076 4616
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 10232 4632 10284 4684
rect 10876 4675 10928 4684
rect 10876 4641 10885 4675
rect 10885 4641 10919 4675
rect 10919 4641 10928 4675
rect 10876 4632 10928 4641
rect 11888 4632 11940 4684
rect 13084 4675 13136 4684
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 13176 4632 13228 4684
rect 13636 4675 13688 4684
rect 13636 4641 13645 4675
rect 13645 4641 13679 4675
rect 13679 4641 13688 4675
rect 13636 4632 13688 4641
rect 15476 4632 15528 4684
rect 17132 4700 17184 4752
rect 17684 4743 17736 4752
rect 10600 4564 10652 4616
rect 16764 4564 16816 4616
rect 17316 4632 17368 4684
rect 17684 4709 17693 4743
rect 17693 4709 17727 4743
rect 17727 4709 17736 4743
rect 17684 4700 17736 4709
rect 19800 4700 19852 4752
rect 20812 4700 20864 4752
rect 21364 4743 21416 4752
rect 21364 4709 21373 4743
rect 21373 4709 21407 4743
rect 21407 4709 21416 4743
rect 21364 4700 21416 4709
rect 24860 4700 24912 4752
rect 26792 4700 26844 4752
rect 27620 4743 27672 4752
rect 27620 4709 27629 4743
rect 27629 4709 27663 4743
rect 27663 4709 27672 4743
rect 27620 4700 27672 4709
rect 27712 4743 27764 4752
rect 27712 4709 27721 4743
rect 27721 4709 27755 4743
rect 27755 4709 27764 4743
rect 28264 4743 28316 4752
rect 27712 4700 27764 4709
rect 28264 4709 28273 4743
rect 28273 4709 28307 4743
rect 28307 4709 28316 4743
rect 28264 4700 28316 4709
rect 18512 4675 18564 4684
rect 18512 4641 18521 4675
rect 18521 4641 18555 4675
rect 18555 4641 18564 4675
rect 18512 4632 18564 4641
rect 18788 4632 18840 4684
rect 19340 4675 19392 4684
rect 19340 4641 19349 4675
rect 19349 4641 19383 4675
rect 19383 4641 19392 4675
rect 19340 4632 19392 4641
rect 19708 4675 19760 4684
rect 19708 4641 19717 4675
rect 19717 4641 19751 4675
rect 19751 4641 19760 4675
rect 19708 4632 19760 4641
rect 20076 4632 20128 4684
rect 21456 4632 21508 4684
rect 22376 4675 22428 4684
rect 22376 4641 22385 4675
rect 22385 4641 22419 4675
rect 22419 4641 22428 4675
rect 22376 4632 22428 4641
rect 22744 4675 22796 4684
rect 22744 4641 22753 4675
rect 22753 4641 22787 4675
rect 22787 4641 22796 4675
rect 22744 4632 22796 4641
rect 23296 4675 23348 4684
rect 23296 4641 23305 4675
rect 23305 4641 23339 4675
rect 23339 4641 23348 4675
rect 23296 4632 23348 4641
rect 23572 4675 23624 4684
rect 23572 4641 23581 4675
rect 23581 4641 23615 4675
rect 23615 4641 23624 4675
rect 23572 4632 23624 4641
rect 26608 4675 26660 4684
rect 26608 4641 26626 4675
rect 26626 4641 26660 4675
rect 26608 4632 26660 4641
rect 29184 4675 29236 4684
rect 29184 4641 29193 4675
rect 29193 4641 29227 4675
rect 29227 4641 29236 4675
rect 29184 4632 29236 4641
rect 30656 4675 30708 4684
rect 30656 4641 30700 4675
rect 30700 4641 30708 4675
rect 30656 4632 30708 4641
rect 21916 4564 21968 4616
rect 24124 4564 24176 4616
rect 24768 4564 24820 4616
rect 26516 4496 26568 4548
rect 3792 4428 3844 4480
rect 4160 4428 4212 4480
rect 9588 4428 9640 4480
rect 11520 4471 11572 4480
rect 11520 4437 11529 4471
rect 11529 4437 11563 4471
rect 11563 4437 11572 4471
rect 11888 4471 11940 4480
rect 11520 4428 11572 4437
rect 11888 4437 11897 4471
rect 11897 4437 11931 4471
rect 11931 4437 11940 4471
rect 11888 4428 11940 4437
rect 14188 4428 14240 4480
rect 16028 4471 16080 4480
rect 16028 4437 16037 4471
rect 16037 4437 16071 4471
rect 16071 4437 16080 4471
rect 16028 4428 16080 4437
rect 22008 4428 22060 4480
rect 22376 4428 22428 4480
rect 26792 4428 26844 4480
rect 29552 4471 29604 4480
rect 29552 4437 29561 4471
rect 29561 4437 29595 4471
rect 29595 4437 29604 4471
rect 29552 4428 29604 4437
rect 30564 4428 30616 4480
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 2136 4224 2188 4276
rect 8208 4224 8260 4276
rect 10600 4267 10652 4276
rect 10600 4233 10609 4267
rect 10609 4233 10643 4267
rect 10643 4233 10652 4267
rect 10600 4224 10652 4233
rect 15476 4267 15528 4276
rect 15476 4233 15485 4267
rect 15485 4233 15519 4267
rect 15519 4233 15528 4267
rect 15476 4224 15528 4233
rect 21732 4224 21784 4276
rect 22744 4224 22796 4276
rect 26608 4224 26660 4276
rect 27620 4224 27672 4276
rect 29184 4224 29236 4276
rect 30656 4224 30708 4276
rect 31300 4267 31352 4276
rect 31300 4233 31309 4267
rect 31309 4233 31343 4267
rect 31343 4233 31352 4267
rect 31300 4224 31352 4233
rect 2964 4156 3016 4208
rect 3608 4156 3660 4208
rect 4436 4088 4488 4140
rect 5080 4088 5132 4140
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 6000 4088 6052 4140
rect 17316 4156 17368 4208
rect 3424 4063 3476 4072
rect 3424 4029 3433 4063
rect 3433 4029 3467 4063
rect 3467 4029 3476 4063
rect 3424 4020 3476 4029
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 8208 4020 8260 4072
rect 17960 4088 18012 4140
rect 20444 4088 20496 4140
rect 21640 4088 21692 4140
rect 22376 4088 22428 4140
rect 22928 4088 22980 4140
rect 23572 4156 23624 4208
rect 23480 4088 23532 4140
rect 9588 4063 9640 4072
rect 2688 3952 2740 4004
rect 4988 3952 5040 4004
rect 5172 3952 5224 4004
rect 6552 3952 6604 4004
rect 8024 3952 8076 4004
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 2504 3927 2556 3936
rect 2504 3893 2513 3927
rect 2513 3893 2547 3927
rect 2547 3893 2556 3927
rect 2504 3884 2556 3893
rect 4252 3927 4304 3936
rect 4252 3893 4261 3927
rect 4261 3893 4295 3927
rect 4295 3893 4304 3927
rect 4252 3884 4304 3893
rect 6000 3884 6052 3936
rect 6460 3927 6512 3936
rect 6460 3893 6469 3927
rect 6469 3893 6503 3927
rect 6503 3893 6512 3927
rect 6460 3884 6512 3893
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 9312 3952 9364 4004
rect 9128 3884 9180 3936
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 10876 4063 10928 4072
rect 9588 4020 9640 4029
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 10876 4020 10928 4029
rect 11888 4020 11940 4072
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 13268 4063 13320 4072
rect 13268 4029 13277 4063
rect 13277 4029 13311 4063
rect 13311 4029 13320 4063
rect 13268 4020 13320 4029
rect 13636 4063 13688 4072
rect 13636 4029 13645 4063
rect 13645 4029 13679 4063
rect 13679 4029 13688 4063
rect 13636 4020 13688 4029
rect 15476 4020 15528 4072
rect 16672 4063 16724 4072
rect 16672 4029 16681 4063
rect 16681 4029 16715 4063
rect 16715 4029 16724 4063
rect 16672 4020 16724 4029
rect 17040 4063 17092 4072
rect 17040 4029 17049 4063
rect 17049 4029 17083 4063
rect 17083 4029 17092 4063
rect 17040 4020 17092 4029
rect 16764 3952 16816 4004
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 12256 3927 12308 3936
rect 12256 3893 12265 3927
rect 12265 3893 12299 3927
rect 12299 3893 12308 3927
rect 12256 3884 12308 3893
rect 13544 3884 13596 3936
rect 14648 3884 14700 3936
rect 15384 3884 15436 3936
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 18512 4020 18564 4072
rect 18788 4063 18840 4072
rect 18788 4029 18797 4063
rect 18797 4029 18831 4063
rect 18831 4029 18840 4063
rect 18788 4020 18840 4029
rect 18880 4063 18932 4072
rect 18880 4029 18889 4063
rect 18889 4029 18923 4063
rect 18923 4029 18932 4063
rect 19248 4063 19300 4072
rect 18880 4020 18932 4029
rect 19248 4029 19257 4063
rect 19257 4029 19291 4063
rect 19291 4029 19300 4063
rect 19248 4020 19300 4029
rect 19708 4020 19760 4072
rect 20352 4063 20404 4072
rect 20352 4029 20361 4063
rect 20361 4029 20395 4063
rect 20395 4029 20404 4063
rect 20352 4020 20404 4029
rect 22100 4063 22152 4072
rect 22100 4029 22109 4063
rect 22109 4029 22143 4063
rect 22143 4029 22152 4063
rect 22100 4020 22152 4029
rect 24676 4020 24728 4072
rect 25320 4020 25372 4072
rect 25504 4020 25556 4072
rect 26516 4063 26568 4072
rect 26516 4029 26525 4063
rect 26525 4029 26559 4063
rect 26559 4029 26568 4063
rect 26516 4020 26568 4029
rect 30472 4088 30524 4140
rect 29092 4020 29144 4072
rect 29736 4063 29788 4072
rect 29736 4029 29745 4063
rect 29745 4029 29779 4063
rect 29779 4029 29788 4063
rect 29736 4020 29788 4029
rect 20812 3952 20864 4004
rect 21456 3952 21508 4004
rect 22836 3952 22888 4004
rect 17408 3884 17460 3893
rect 17868 3884 17920 3936
rect 22560 3884 22612 3936
rect 23296 3884 23348 3936
rect 23480 3927 23532 3936
rect 23480 3893 23489 3927
rect 23489 3893 23523 3927
rect 23523 3893 23532 3927
rect 23480 3884 23532 3893
rect 24768 3952 24820 4004
rect 26792 3952 26844 4004
rect 27712 3952 27764 4004
rect 30380 3995 30432 4004
rect 30380 3961 30389 3995
rect 30389 3961 30423 3995
rect 30423 3961 30432 3995
rect 30380 3952 30432 3961
rect 30472 3995 30524 4004
rect 30472 3961 30481 3995
rect 30481 3961 30515 3995
rect 30515 3961 30524 3995
rect 31024 3995 31076 4004
rect 30472 3952 30524 3961
rect 31024 3961 31033 3995
rect 31033 3961 31067 3995
rect 31067 3961 31076 3995
rect 31024 3952 31076 3961
rect 24860 3927 24912 3936
rect 24860 3893 24869 3927
rect 24869 3893 24903 3927
rect 24903 3893 24912 3927
rect 24860 3884 24912 3893
rect 25872 3884 25924 3936
rect 29276 3884 29328 3936
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 1860 3680 1912 3732
rect 2596 3680 2648 3732
rect 3424 3680 3476 3732
rect 4988 3680 5040 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 6644 3723 6696 3732
rect 5080 3680 5132 3689
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 11520 3680 11572 3732
rect 12532 3723 12584 3732
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 13268 3680 13320 3732
rect 15476 3680 15528 3732
rect 16764 3723 16816 3732
rect 16764 3689 16773 3723
rect 16773 3689 16807 3723
rect 16807 3689 16816 3723
rect 16764 3680 16816 3689
rect 18788 3680 18840 3732
rect 21916 3680 21968 3732
rect 22376 3680 22428 3732
rect 25872 3723 25924 3732
rect 8760 3655 8812 3664
rect 8760 3621 8769 3655
rect 8769 3621 8803 3655
rect 8803 3621 8812 3655
rect 8760 3612 8812 3621
rect 10600 3612 10652 3664
rect 2780 3544 2832 3596
rect 3608 3544 3660 3596
rect 5172 3544 5224 3596
rect 6000 3587 6052 3596
rect 6000 3553 6009 3587
rect 6009 3553 6043 3587
rect 6043 3553 6052 3587
rect 6000 3544 6052 3553
rect 6644 3587 6696 3596
rect 5448 3476 5500 3528
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 9036 3544 9088 3596
rect 9772 3544 9824 3596
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 11796 3587 11848 3596
rect 11796 3553 11805 3587
rect 11805 3553 11839 3587
rect 11839 3553 11848 3587
rect 11796 3544 11848 3553
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 14280 3544 14332 3553
rect 15292 3655 15344 3664
rect 15292 3621 15301 3655
rect 15301 3621 15335 3655
rect 15335 3621 15344 3655
rect 15292 3612 15344 3621
rect 16488 3612 16540 3664
rect 20352 3612 20404 3664
rect 20628 3612 20680 3664
rect 21272 3612 21324 3664
rect 17408 3544 17460 3596
rect 17960 3587 18012 3596
rect 17960 3553 17969 3587
rect 17969 3553 18003 3587
rect 18003 3553 18012 3587
rect 17960 3544 18012 3553
rect 18328 3587 18380 3596
rect 18328 3553 18337 3587
rect 18337 3553 18371 3587
rect 18371 3553 18380 3587
rect 18328 3544 18380 3553
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 14556 3476 14608 3528
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 17132 3476 17184 3528
rect 19248 3544 19300 3596
rect 24768 3612 24820 3664
rect 25872 3689 25881 3723
rect 25881 3689 25915 3723
rect 25915 3689 25924 3723
rect 25872 3680 25924 3689
rect 28264 3680 28316 3732
rect 30380 3723 30432 3732
rect 30380 3689 30389 3723
rect 30389 3689 30423 3723
rect 30423 3689 30432 3723
rect 30380 3680 30432 3689
rect 30472 3680 30524 3732
rect 25412 3612 25464 3664
rect 26148 3612 26200 3664
rect 26332 3612 26384 3664
rect 26792 3612 26844 3664
rect 28540 3612 28592 3664
rect 29184 3612 29236 3664
rect 30564 3655 30616 3664
rect 30564 3621 30573 3655
rect 30573 3621 30607 3655
rect 30607 3621 30616 3655
rect 30564 3612 30616 3621
rect 30656 3655 30708 3664
rect 30656 3621 30665 3655
rect 30665 3621 30699 3655
rect 30699 3621 30708 3655
rect 30656 3612 30708 3621
rect 19800 3519 19852 3528
rect 19800 3485 19809 3519
rect 19809 3485 19843 3519
rect 19843 3485 19852 3519
rect 19800 3476 19852 3485
rect 22744 3544 22796 3596
rect 23296 3544 23348 3596
rect 23756 3587 23808 3596
rect 9128 3408 9180 3460
rect 11060 3451 11112 3460
rect 11060 3417 11069 3451
rect 11069 3417 11103 3451
rect 11103 3417 11112 3451
rect 11060 3408 11112 3417
rect 15384 3408 15436 3460
rect 15568 3451 15620 3460
rect 15568 3417 15577 3451
rect 15577 3417 15611 3451
rect 15611 3417 15620 3451
rect 15568 3408 15620 3417
rect 20536 3408 20588 3460
rect 22284 3408 22336 3460
rect 13636 3340 13688 3392
rect 14924 3340 14976 3392
rect 23756 3553 23765 3587
rect 23765 3553 23799 3587
rect 23799 3553 23808 3587
rect 23756 3544 23808 3553
rect 32220 3587 32272 3596
rect 32220 3553 32229 3587
rect 32229 3553 32263 3587
rect 32263 3553 32272 3587
rect 32220 3544 32272 3553
rect 24952 3476 25004 3528
rect 26424 3476 26476 3528
rect 31024 3519 31076 3528
rect 31024 3485 31033 3519
rect 31033 3485 31067 3519
rect 31067 3485 31076 3519
rect 31024 3476 31076 3485
rect 28908 3408 28960 3460
rect 20628 3340 20680 3392
rect 20812 3340 20864 3392
rect 22376 3383 22428 3392
rect 22376 3349 22385 3383
rect 22385 3349 22419 3383
rect 22419 3349 22428 3383
rect 22376 3340 22428 3349
rect 23480 3340 23532 3392
rect 24584 3383 24636 3392
rect 24584 3349 24593 3383
rect 24593 3349 24627 3383
rect 24627 3349 24636 3383
rect 24584 3340 24636 3349
rect 26240 3383 26292 3392
rect 26240 3349 26249 3383
rect 26249 3349 26283 3383
rect 26283 3349 26292 3383
rect 26240 3340 26292 3349
rect 27436 3383 27488 3392
rect 27436 3349 27445 3383
rect 27445 3349 27479 3383
rect 27479 3349 27488 3383
rect 27436 3340 27488 3349
rect 32496 3340 32548 3392
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 1768 3179 1820 3188
rect 1768 3145 1777 3179
rect 1777 3145 1811 3179
rect 1811 3145 1820 3179
rect 1768 3136 1820 3145
rect 2780 3136 2832 3188
rect 1860 3068 1912 3120
rect 4068 3111 4120 3120
rect 4068 3077 4077 3111
rect 4077 3077 4111 3111
rect 4111 3077 4120 3111
rect 4068 3068 4120 3077
rect 1768 2932 1820 2984
rect 2964 2975 3016 2984
rect 2964 2941 2973 2975
rect 2973 2941 3007 2975
rect 3007 2941 3016 2975
rect 2964 2932 3016 2941
rect 3516 2975 3568 2984
rect 3240 2864 3292 2916
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 3792 2932 3844 2984
rect 6644 3136 6696 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 14280 3136 14332 3188
rect 14556 3179 14608 3188
rect 14556 3145 14580 3179
rect 14580 3145 14608 3179
rect 14556 3136 14608 3145
rect 5172 3068 5224 3120
rect 6000 3000 6052 3052
rect 3608 2864 3660 2916
rect 7012 2975 7064 2984
rect 7012 2941 7021 2975
rect 7021 2941 7055 2975
rect 7055 2941 7064 2975
rect 7012 2932 7064 2941
rect 14004 3068 14056 3120
rect 15292 3136 15344 3188
rect 15568 3136 15620 3188
rect 17132 3179 17184 3188
rect 17132 3145 17141 3179
rect 17141 3145 17175 3179
rect 17175 3145 17184 3179
rect 17132 3136 17184 3145
rect 17960 3136 18012 3188
rect 18512 3136 18564 3188
rect 20812 3136 20864 3188
rect 22744 3136 22796 3188
rect 23572 3136 23624 3188
rect 25412 3179 25464 3188
rect 25412 3145 25421 3179
rect 25421 3145 25455 3179
rect 25455 3145 25464 3179
rect 25412 3136 25464 3145
rect 28540 3179 28592 3188
rect 28540 3145 28549 3179
rect 28549 3145 28583 3179
rect 28583 3145 28592 3179
rect 28540 3136 28592 3145
rect 30656 3136 30708 3188
rect 32220 3179 32272 3188
rect 32220 3145 32229 3179
rect 32229 3145 32263 3179
rect 32263 3145 32272 3179
rect 32220 3136 32272 3145
rect 7840 2932 7892 2984
rect 8208 2932 8260 2984
rect 8576 2932 8628 2984
rect 9312 3000 9364 3052
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 9128 2932 9180 2984
rect 8116 2864 8168 2916
rect 9588 2932 9640 2984
rect 11060 2932 11112 2984
rect 12256 2975 12308 2984
rect 12256 2941 12265 2975
rect 12265 2941 12299 2975
rect 12299 2941 12308 2975
rect 12256 2932 12308 2941
rect 13728 2932 13780 2984
rect 15384 3000 15436 3052
rect 22652 3111 22704 3120
rect 22652 3077 22661 3111
rect 22661 3077 22695 3111
rect 22695 3077 22704 3111
rect 22652 3068 22704 3077
rect 24860 3068 24912 3120
rect 26332 3068 26384 3120
rect 16304 2932 16356 2984
rect 16580 2975 16632 2984
rect 16580 2941 16589 2975
rect 16589 2941 16623 2975
rect 16623 2941 16632 2975
rect 16580 2932 16632 2941
rect 17408 2932 17460 2984
rect 22376 3000 22428 3052
rect 18880 2975 18932 2984
rect 18880 2941 18889 2975
rect 18889 2941 18923 2975
rect 18923 2941 18932 2975
rect 18880 2932 18932 2941
rect 19248 2975 19300 2984
rect 19248 2941 19257 2975
rect 19257 2941 19291 2975
rect 19291 2941 19300 2975
rect 19248 2932 19300 2941
rect 21640 2932 21692 2984
rect 21916 2975 21968 2984
rect 21916 2941 21925 2975
rect 21925 2941 21959 2975
rect 21959 2941 21968 2975
rect 21916 2932 21968 2941
rect 22100 2932 22152 2984
rect 22468 2932 22520 2984
rect 23756 3000 23808 3052
rect 26240 3043 26292 3052
rect 24124 2975 24176 2984
rect 10968 2907 11020 2916
rect 10968 2873 10977 2907
rect 10977 2873 11011 2907
rect 11011 2873 11020 2907
rect 10968 2864 11020 2873
rect 11796 2864 11848 2916
rect 12624 2864 12676 2916
rect 14924 2864 14976 2916
rect 15108 2907 15160 2916
rect 15108 2873 15117 2907
rect 15117 2873 15151 2907
rect 15151 2873 15160 2907
rect 15108 2864 15160 2873
rect 19524 2864 19576 2916
rect 20720 2864 20772 2916
rect 22376 2864 22428 2916
rect 22560 2864 22612 2916
rect 23480 2864 23532 2916
rect 24124 2941 24133 2975
rect 24133 2941 24167 2975
rect 24167 2941 24176 2975
rect 24124 2932 24176 2941
rect 24584 2975 24636 2984
rect 24584 2941 24593 2975
rect 24593 2941 24627 2975
rect 24627 2941 24636 2975
rect 24584 2932 24636 2941
rect 26240 3009 26249 3043
rect 26249 3009 26283 3043
rect 26283 3009 26292 3043
rect 26240 3000 26292 3009
rect 29276 3043 29328 3052
rect 29276 3009 29285 3043
rect 29285 3009 29319 3043
rect 29319 3009 29328 3043
rect 29276 3000 29328 3009
rect 31300 3000 31352 3052
rect 32036 3000 32088 3052
rect 32496 3043 32548 3052
rect 26424 2932 26476 2984
rect 29000 2932 29052 2984
rect 29092 2975 29144 2984
rect 29092 2941 29101 2975
rect 29101 2941 29135 2975
rect 29135 2941 29144 2975
rect 29092 2932 29144 2941
rect 26332 2864 26384 2916
rect 30932 2864 30984 2916
rect 31208 2864 31260 2916
rect 32496 3009 32505 3043
rect 32505 3009 32539 3043
rect 32539 3009 32548 3043
rect 32496 3000 32548 3009
rect 32588 2907 32640 2916
rect 32588 2873 32597 2907
rect 32597 2873 32631 2907
rect 32631 2873 32640 2907
rect 32588 2864 32640 2873
rect 5264 2796 5316 2848
rect 5356 2796 5408 2848
rect 5540 2839 5592 2848
rect 5540 2805 5549 2839
rect 5549 2805 5583 2839
rect 5583 2805 5592 2839
rect 5540 2796 5592 2805
rect 7932 2839 7984 2848
rect 7932 2805 7941 2839
rect 7941 2805 7975 2839
rect 7975 2805 7984 2839
rect 7932 2796 7984 2805
rect 8300 2839 8352 2848
rect 8300 2805 8309 2839
rect 8309 2805 8343 2839
rect 8343 2805 8352 2839
rect 8300 2796 8352 2805
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 18696 2796 18748 2848
rect 27436 2839 27488 2848
rect 27436 2805 27445 2839
rect 27445 2805 27479 2839
rect 27479 2805 27488 2839
rect 27436 2796 27488 2805
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 2964 2592 3016 2644
rect 3240 2592 3292 2644
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 8576 2635 8628 2644
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 8852 2635 8904 2644
rect 8852 2601 8861 2635
rect 8861 2601 8895 2635
rect 8895 2601 8904 2635
rect 8852 2592 8904 2601
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12808 2635 12860 2644
rect 12440 2592 12492 2601
rect 12808 2601 12817 2635
rect 12817 2601 12851 2635
rect 12851 2601 12860 2635
rect 12808 2592 12860 2601
rect 13728 2635 13780 2644
rect 13728 2601 13737 2635
rect 13737 2601 13771 2635
rect 13771 2601 13780 2635
rect 13728 2592 13780 2601
rect 13912 2592 13964 2644
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 15660 2592 15712 2644
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 19340 2592 19392 2644
rect 20260 2592 20312 2644
rect 20628 2635 20680 2644
rect 20628 2601 20637 2635
rect 20637 2601 20671 2635
rect 20671 2601 20680 2635
rect 20628 2592 20680 2601
rect 29000 2592 29052 2644
rect 29552 2635 29604 2644
rect 3516 2524 3568 2576
rect 5448 2524 5500 2576
rect 8116 2524 8168 2576
rect 10968 2524 11020 2576
rect 11428 2567 11480 2576
rect 11428 2533 11437 2567
rect 11437 2533 11471 2567
rect 11471 2533 11480 2567
rect 11428 2524 11480 2533
rect 3240 2456 3292 2508
rect 7932 2456 7984 2508
rect 8668 2499 8720 2508
rect 8668 2465 8677 2499
rect 8677 2465 8711 2499
rect 8711 2465 8720 2499
rect 8668 2456 8720 2465
rect 16856 2567 16908 2576
rect 16856 2533 16865 2567
rect 16865 2533 16899 2567
rect 16899 2533 16908 2567
rect 16856 2524 16908 2533
rect 13728 2456 13780 2508
rect 13912 2456 13964 2508
rect 15108 2456 15160 2508
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 14188 2388 14240 2397
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 9036 2320 9088 2372
rect 10508 2363 10560 2372
rect 10508 2329 10517 2363
rect 10517 2329 10551 2363
rect 10551 2329 10560 2363
rect 10508 2320 10560 2329
rect 14924 2320 14976 2372
rect 15660 2363 15712 2372
rect 15660 2329 15669 2363
rect 15669 2329 15703 2363
rect 15703 2329 15712 2363
rect 15660 2320 15712 2329
rect 17408 2499 17460 2508
rect 17408 2465 17417 2499
rect 17417 2465 17451 2499
rect 17451 2465 17460 2499
rect 17408 2456 17460 2465
rect 16764 2431 16816 2440
rect 16764 2397 16773 2431
rect 16773 2397 16807 2431
rect 16807 2397 16816 2431
rect 16764 2388 16816 2397
rect 19524 2567 19576 2576
rect 19524 2533 19533 2567
rect 19533 2533 19567 2567
rect 19567 2533 19576 2567
rect 19524 2524 19576 2533
rect 23112 2567 23164 2576
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 20076 2499 20128 2508
rect 20076 2465 20120 2499
rect 20120 2465 20128 2499
rect 20076 2456 20128 2465
rect 20536 2456 20588 2508
rect 21548 2456 21600 2508
rect 23112 2533 23121 2567
rect 23121 2533 23155 2567
rect 23155 2533 23164 2567
rect 23112 2524 23164 2533
rect 22100 2499 22152 2508
rect 22100 2465 22109 2499
rect 22109 2465 22143 2499
rect 22143 2465 22152 2499
rect 22100 2456 22152 2465
rect 22376 2456 22428 2508
rect 22928 2456 22980 2508
rect 23480 2499 23532 2508
rect 23480 2465 23489 2499
rect 23489 2465 23523 2499
rect 23523 2465 23532 2499
rect 23480 2456 23532 2465
rect 24124 2456 24176 2508
rect 25044 2499 25096 2508
rect 25044 2465 25053 2499
rect 25053 2465 25087 2499
rect 25087 2465 25096 2499
rect 25044 2456 25096 2465
rect 26332 2524 26384 2576
rect 27160 2524 27212 2576
rect 27620 2524 27672 2576
rect 29552 2601 29561 2635
rect 29561 2601 29595 2635
rect 29595 2601 29604 2635
rect 30932 2635 30984 2644
rect 29552 2592 29604 2601
rect 30932 2601 30941 2635
rect 30941 2601 30975 2635
rect 30975 2601 30984 2635
rect 30932 2592 30984 2601
rect 31300 2635 31352 2644
rect 31300 2601 31309 2635
rect 31309 2601 31343 2635
rect 31343 2601 31352 2635
rect 31300 2592 31352 2601
rect 31668 2592 31720 2644
rect 32036 2635 32088 2644
rect 32036 2601 32045 2635
rect 32045 2601 32079 2635
rect 32079 2601 32088 2635
rect 32036 2592 32088 2601
rect 27436 2456 27488 2508
rect 27804 2499 27856 2508
rect 27804 2465 27813 2499
rect 27813 2465 27847 2499
rect 27847 2465 27856 2499
rect 27804 2456 27856 2465
rect 28908 2456 28960 2508
rect 32588 2524 32640 2576
rect 30932 2388 30984 2440
rect 28908 2320 28960 2372
rect 31300 2320 31352 2372
rect 13820 2252 13872 2304
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
rect 19340 8 19392 60
rect 28908 8 28960 60
<< metal2 >>
rect 1766 15600 1822 15609
rect 1766 15535 1822 15544
rect 1490 12880 1546 12889
rect 1490 12815 1546 12824
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10810 1440 11154
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1504 10418 1532 12815
rect 1582 12064 1638 12073
rect 1582 11999 1638 12008
rect 1596 11354 1624 11999
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1582 11112 1638 11121
rect 1582 11047 1638 11056
rect 1412 10390 1532 10418
rect 1412 5370 1440 10390
rect 1490 10296 1546 10305
rect 1596 10266 1624 11047
rect 1490 10231 1546 10240
rect 1584 10260 1636 10266
rect 1504 9178 1532 10231
rect 1584 10202 1636 10208
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1688 9382 1716 10066
rect 1676 9376 1728 9382
rect 1582 9344 1638 9353
rect 1676 9318 1728 9324
rect 1582 9279 1638 9288
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1596 8090 1624 9279
rect 1688 8945 1716 9318
rect 1674 8936 1730 8945
rect 1674 8871 1730 8880
rect 1780 8634 1808 15535
rect 6642 15520 6698 16000
rect 19982 15520 20038 16000
rect 33322 15520 33378 16000
rect 35530 15600 35586 15609
rect 35530 15535 35586 15544
rect 1858 14648 1914 14657
rect 1858 14583 1914 14592
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1872 7546 1900 14583
rect 1950 13832 2006 13841
rect 1950 13767 2006 13776
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1688 7002 1716 7278
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1964 6458 1992 13767
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2042 9072 2098 9081
rect 2700 9042 2728 10746
rect 3422 9616 3478 9625
rect 3422 9551 3478 9560
rect 3436 9042 3464 9551
rect 2042 9007 2044 9016
rect 2096 9007 2098 9016
rect 2688 9036 2740 9042
rect 2044 8978 2096 8984
rect 2688 8978 2740 8984
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 2056 8634 2084 8978
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2596 8560 2648 8566
rect 2502 8528 2558 8537
rect 2596 8502 2648 8508
rect 2502 8463 2558 8472
rect 2516 8090 2544 8463
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2056 7857 2084 7890
rect 2042 7848 2098 7857
rect 2042 7783 2098 7792
rect 2056 7546 2084 7783
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2516 7478 2544 7890
rect 2608 7585 2636 8502
rect 2700 8129 2728 8774
rect 3436 8634 3464 8978
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 5448 8560 5500 8566
rect 5078 8528 5134 8537
rect 3976 8492 4028 8498
rect 5448 8502 5500 8508
rect 5078 8463 5080 8472
rect 3976 8434 4028 8440
rect 5132 8463 5134 8472
rect 5080 8434 5132 8440
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2686 8120 2742 8129
rect 2686 8055 2742 8064
rect 2594 7576 2650 7585
rect 2594 7511 2650 7520
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 2424 6390 2452 6802
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2424 6202 2452 6326
rect 2332 6186 2452 6202
rect 2320 6180 2452 6186
rect 2372 6174 2452 6180
rect 2320 6122 2372 6128
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2056 5953 2084 6054
rect 2042 5944 2098 5953
rect 2042 5879 2098 5888
rect 2424 5846 2452 6174
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 2042 5264 2098 5273
rect 2042 5199 2044 5208
rect 2096 5199 2098 5208
rect 2044 5170 2096 5176
rect 2148 5166 2176 5510
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2148 4758 2176 5102
rect 2240 4826 2268 5646
rect 2424 5370 2452 5782
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1780 3194 1808 4626
rect 2148 4282 2176 4694
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2516 3942 2544 6598
rect 2792 6322 2820 6666
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2596 5636 2648 5642
rect 2596 5578 2648 5584
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2608 5234 2636 5578
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2700 4842 2728 5578
rect 2792 5030 2820 6258
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2608 4814 2728 4842
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 1872 3738 1900 3878
rect 2608 3738 2636 4814
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2700 4010 2728 4626
rect 2778 4040 2834 4049
rect 2688 4004 2740 4010
rect 2778 3975 2834 3984
rect 2688 3946 2740 3952
rect 2792 3777 2820 3975
rect 2778 3768 2834 3777
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2596 3732 2648 3738
rect 2778 3703 2834 3712
rect 2596 3674 2648 3680
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1780 2990 1808 3130
rect 1872 3126 1900 3674
rect 2792 3602 2820 3703
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2792 3194 2820 3538
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1766 2408 1822 2417
rect 1766 2343 1822 2352
rect 1780 480 1808 2343
rect 2884 513 2912 8366
rect 3068 8265 3096 8366
rect 3054 8256 3110 8265
rect 3054 8191 3110 8200
rect 3148 7744 3200 7750
rect 3988 7721 4016 8434
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4080 8242 4108 8366
rect 4080 8214 4200 8242
rect 4172 7886 4200 8214
rect 5078 8120 5134 8129
rect 5078 8055 5080 8064
rect 5132 8055 5134 8064
rect 5080 8026 5132 8032
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3148 7686 3200 7692
rect 3974 7712 4030 7721
rect 3160 7274 3188 7686
rect 3974 7647 4030 7656
rect 4172 7546 4200 7822
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3700 7472 3752 7478
rect 3700 7414 3752 7420
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3252 7274 3280 7346
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 6458 3280 7210
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2976 4214 3004 4558
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3436 3913 3464 4014
rect 3422 3904 3478 3913
rect 3422 3839 3478 3848
rect 3436 3738 3464 3839
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 2962 3496 3018 3505
rect 2962 3431 3018 3440
rect 2976 2990 3004 3431
rect 3528 2990 3556 5102
rect 3620 5098 3648 5510
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3620 4593 3648 5034
rect 3712 4690 3740 7414
rect 4264 7410 4292 7958
rect 4342 7576 4398 7585
rect 4342 7511 4398 7520
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 5846 3924 6734
rect 3884 5840 3936 5846
rect 3884 5782 3936 5788
rect 3896 5642 3924 5782
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3606 4584 3662 4593
rect 3606 4519 3662 4528
rect 3620 4214 3648 4519
rect 3804 4486 3832 5102
rect 3988 4826 4016 7142
rect 4172 6882 4200 7142
rect 4080 6854 4200 6882
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4080 6662 4108 6854
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6458 4108 6598
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4080 6118 4108 6394
rect 4264 6390 4292 6870
rect 4356 6798 4384 7511
rect 5092 7478 5120 8026
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 5184 7410 5212 7822
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4264 5778 4292 6326
rect 4356 6322 4384 6734
rect 4448 6730 4476 7278
rect 5184 6934 5212 7346
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5460 6882 5488 8502
rect 5630 8120 5686 8129
rect 6656 8090 6684 15520
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 16670 11656 16726 11665
rect 16670 11591 16726 11600
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 12990 9072 13046 9081
rect 12990 9007 13046 9016
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 13004 8401 13032 9007
rect 12990 8392 13046 8401
rect 12990 8327 13046 8336
rect 5630 8055 5686 8064
rect 6644 8084 6696 8090
rect 5644 7721 5672 8055
rect 6644 8026 6696 8032
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 5630 7712 5686 7721
rect 5630 7647 5686 7656
rect 5920 7206 5948 7890
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 6826 7440 6882 7449
rect 6826 7375 6882 7384
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5816 6928 5868 6934
rect 5460 6854 5764 6882
rect 5816 6870 5868 6876
rect 5736 6798 5764 6854
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4448 6322 4476 6666
rect 5736 6458 5764 6734
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5828 6390 5856 6870
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4356 5846 4384 6122
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 4080 4434 4108 5646
rect 4356 5098 4384 5782
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4160 4480 4212 4486
rect 4080 4428 4160 4434
rect 4080 4422 4212 4428
rect 3608 4208 3660 4214
rect 3608 4150 3660 4156
rect 3620 3602 3648 4150
rect 3804 4078 3832 4422
rect 4080 4406 4200 4422
rect 3974 4176 4030 4185
rect 3974 4111 4030 4120
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 2976 2650 3004 2926
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 3252 2650 3280 2858
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3252 2514 3280 2586
rect 3528 2582 3556 2926
rect 3620 2922 3648 3538
rect 3804 2990 3832 4014
rect 3988 3097 4016 4111
rect 4080 3126 4108 4406
rect 4264 3942 4292 4626
rect 4448 4146 4476 6258
rect 5920 6225 5948 7142
rect 6840 6633 6868 7375
rect 9876 7206 9904 7890
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10690 7712 10746 7721
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9508 6882 9536 6938
rect 9692 6882 9720 6938
rect 9508 6854 9720 6882
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 6826 6624 6882 6633
rect 6826 6559 6882 6568
rect 6932 6322 6960 6734
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8772 6458 8800 6734
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 6225 7236 6258
rect 9876 6225 9904 7142
rect 10336 6934 10364 7686
rect 10690 7647 10746 7656
rect 10704 7206 10732 7647
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 5906 6216 5962 6225
rect 5460 6174 5906 6202
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 5000 4010 5028 5510
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5092 4826 5120 5102
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4068 3120 4120 3126
rect 3974 3088 4030 3097
rect 4068 3062 4120 3068
rect 3974 3023 4030 3032
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3516 2576 3568 2582
rect 3516 2518 3568 2524
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 2870 504 2926 513
rect 1766 0 1822 480
rect 2870 439 2926 448
rect 4264 241 4292 3878
rect 5000 3738 5028 3946
rect 5092 3738 5120 4082
rect 5184 4010 5212 4626
rect 5460 4146 5488 6174
rect 5906 6151 5962 6160
rect 7194 6216 7250 6225
rect 9862 6216 9918 6225
rect 7194 6151 7250 6160
rect 9128 6180 9180 6186
rect 5920 6091 5948 6151
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6288 5098 6316 5782
rect 6564 5370 6592 6054
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6656 5030 6684 5646
rect 7208 5642 7236 6151
rect 9680 6180 9732 6186
rect 9128 6122 9180 6128
rect 9508 6140 9680 6168
rect 9140 5914 9168 6122
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7392 5370 7420 5646
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 5908 4684 5960 4690
rect 6552 4684 6604 4690
rect 5960 4644 6040 4672
rect 5908 4626 5960 4632
rect 6012 4146 6040 4644
rect 6552 4626 6604 4632
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5184 3602 5212 3946
rect 6012 3942 6040 4082
rect 6472 3942 6500 4558
rect 6564 4010 6592 4626
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6000 3936 6052 3942
rect 5262 3904 5318 3913
rect 6460 3936 6512 3942
rect 6000 3878 6052 3884
rect 6458 3904 6460 3913
rect 6512 3904 6514 3913
rect 5262 3839 5318 3848
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5184 3126 5212 3538
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5276 2854 5304 3839
rect 6012 3602 6040 3878
rect 6458 3839 6514 3848
rect 6000 3596 6052 3602
rect 6564 3584 6592 3946
rect 6656 3738 6684 4966
rect 7484 4826 7512 5782
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 8220 5234 8248 5510
rect 9140 5370 9168 5850
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 8208 5228 8260 5234
rect 8260 5188 8340 5216
rect 8208 5170 8260 5176
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 8220 4758 8248 5034
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 8036 4010 8064 4558
rect 8220 4282 8248 4694
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 8220 3942 8248 4014
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6644 3596 6696 3602
rect 6564 3556 6644 3584
rect 6000 3538 6052 3544
rect 6644 3538 6696 3544
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5368 480 5396 2790
rect 5460 2582 5488 3470
rect 6012 3058 6040 3538
rect 6656 3194 6684 3538
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 8220 2990 8248 3878
rect 7012 2984 7064 2990
rect 7010 2952 7012 2961
rect 7840 2984 7892 2990
rect 7064 2952 7066 2961
rect 7840 2926 7892 2932
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 7010 2887 7066 2896
rect 5540 2848 5592 2854
rect 5538 2816 5540 2825
rect 5592 2816 5594 2825
rect 5538 2751 5594 2760
rect 7852 2650 7880 2926
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 7944 2514 7972 2790
rect 8128 2582 8156 2858
rect 8312 2854 8340 5188
rect 9508 4826 9536 6140
rect 9862 6151 9918 6160
rect 9680 6122 9732 6128
rect 9876 5953 9904 6151
rect 9862 5944 9918 5953
rect 10336 5914 10364 6870
rect 10428 6458 10456 6870
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 9862 5879 9918 5888
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10428 5846 10456 6394
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10428 5370 10456 5782
rect 10520 5710 10548 7142
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6322 10640 6598
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9600 4826 9628 5102
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 10152 4690 10180 5170
rect 10598 4992 10654 5001
rect 10598 4927 10654 4936
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10152 4593 10180 4626
rect 10138 4584 10194 4593
rect 10138 4519 10194 4528
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 4078 9628 4422
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9128 3936 9180 3942
rect 9126 3904 9128 3913
rect 9180 3904 9182 3913
rect 9126 3839 9182 3848
rect 9140 3738 9168 3839
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 9126 3632 9182 3641
rect 8772 3505 8800 3606
rect 9036 3596 9088 3602
rect 9126 3567 9182 3576
rect 9036 3538 9088 3544
rect 8758 3496 8814 3505
rect 8758 3431 8814 3440
rect 8850 3360 8906 3369
rect 8850 3295 8906 3304
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8588 2650 8616 2926
rect 8666 2816 8722 2825
rect 8666 2751 8722 2760
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 8680 2514 8708 2751
rect 8864 2650 8892 3295
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 9048 2378 9076 3538
rect 9140 3466 9168 3567
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 9140 2990 9168 3402
rect 9324 3233 9352 3946
rect 9310 3224 9366 3233
rect 9310 3159 9366 3168
rect 9324 3058 9352 3159
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9600 2990 9628 4014
rect 10152 3602 10180 4519
rect 10244 3942 10272 4626
rect 10612 4622 10640 4927
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10612 4282 10640 4558
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10244 3777 10272 3878
rect 10230 3768 10286 3777
rect 10230 3703 10286 3712
rect 10612 3670 10640 4218
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 9784 3194 9812 3538
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 10704 2689 10732 7142
rect 13004 6866 13032 8327
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 7585 14228 7890
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14186 7576 14242 7585
rect 14186 7511 14242 7520
rect 14370 7576 14426 7585
rect 14370 7511 14372 7520
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 13726 7304 13782 7313
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 11336 6656 11388 6662
rect 11334 6624 11336 6633
rect 11388 6624 11390 6633
rect 11334 6559 11390 6568
rect 13004 6458 13032 6802
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 11164 5817 11192 6326
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 11150 5808 11206 5817
rect 11150 5743 11206 5752
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5370 11100 5646
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10888 4078 10916 4626
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 11532 3738 11560 4422
rect 11808 3942 11836 4966
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11900 4486 11928 4626
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4078 11928 4422
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11808 3602 11836 3878
rect 12268 3641 12296 3878
rect 12254 3632 12310 3641
rect 11796 3596 11848 3602
rect 12254 3567 12310 3576
rect 11796 3538 11848 3544
rect 11058 3496 11114 3505
rect 11058 3431 11060 3440
rect 11112 3431 11114 3440
rect 11060 3402 11112 3408
rect 11072 2990 11100 3402
rect 11518 3088 11574 3097
rect 11518 3023 11520 3032
rect 11572 3023 11574 3032
rect 11520 2994 11572 3000
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11808 2922 11836 3538
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 3233 11928 3470
rect 11886 3224 11942 3233
rect 11886 3159 11942 3168
rect 12452 3058 12480 6190
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12544 5166 12572 5782
rect 12636 5642 12664 6054
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12912 5370 12940 5782
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12544 5001 12572 5102
rect 12530 4992 12586 5001
rect 12530 4927 12586 4936
rect 12544 4321 12572 4927
rect 13096 4842 13124 7278
rect 13726 7239 13728 7248
rect 13780 7239 13782 7248
rect 13728 7210 13780 7216
rect 14200 7206 14228 7511
rect 14424 7511 14426 7520
rect 14372 7482 14424 7488
rect 14476 7410 14504 7686
rect 16684 7546 16712 11591
rect 19996 10713 20024 15520
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 33336 11665 33364 15520
rect 35254 13832 35310 13841
rect 35254 13767 35310 13776
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 35070 12880 35126 12889
rect 35070 12815 35126 12824
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 33322 11656 33378 11665
rect 33322 11591 33378 11600
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 19982 10704 20038 10713
rect 19982 10639 20038 10648
rect 23386 10704 23442 10713
rect 23386 10639 23442 10648
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 18878 9480 18934 9489
rect 18878 9415 18934 9424
rect 17222 7712 17278 7721
rect 17222 7647 17278 7656
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 16672 7336 16724 7342
rect 15382 7304 15438 7313
rect 14832 7268 14884 7274
rect 16672 7278 16724 7284
rect 15382 7239 15438 7248
rect 14832 7210 14884 7216
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 13636 6656 13688 6662
rect 14016 6633 14044 6734
rect 13636 6598 13688 6604
rect 14002 6624 14058 6633
rect 13648 6254 13676 6598
rect 14002 6559 14058 6568
rect 14016 6390 14044 6559
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 13556 5846 13584 6122
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13280 5166 13308 5578
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13004 4814 13124 4842
rect 12806 4448 12862 4457
rect 12806 4383 12862 4392
rect 12530 4312 12586 4321
rect 12530 4247 12586 4256
rect 12530 3768 12586 3777
rect 12530 3703 12532 3712
rect 12584 3703 12586 3712
rect 12532 3674 12584 3680
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 10690 2680 10746 2689
rect 10690 2615 10746 2624
rect 10980 2582 11008 2858
rect 12268 2825 12296 2926
rect 12254 2816 12310 2825
rect 12254 2751 12310 2760
rect 12452 2650 12480 2994
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 10968 2576 11020 2582
rect 11428 2576 11480 2582
rect 10968 2518 11020 2524
rect 11426 2544 11428 2553
rect 11480 2544 11482 2553
rect 11426 2479 11482 2488
rect 12072 2440 12124 2446
rect 10506 2408 10562 2417
rect 9036 2372 9088 2378
rect 10506 2343 10508 2352
rect 9036 2314 9088 2320
rect 10560 2343 10562 2352
rect 12070 2408 12072 2417
rect 12124 2408 12126 2417
rect 12070 2343 12126 2352
rect 10508 2314 10560 2320
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 9048 480 9076 2314
rect 12636 480 12664 2858
rect 12820 2650 12848 4383
rect 13004 2802 13032 4814
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13176 4684 13228 4690
rect 13280 4672 13308 5102
rect 13228 4644 13308 4672
rect 13176 4626 13228 4632
rect 13096 4078 13124 4626
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13188 3641 13216 4626
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13280 3738 13308 4014
rect 13556 3942 13584 5646
rect 13648 5030 13676 6190
rect 14108 5914 14136 6734
rect 14844 6662 14872 7210
rect 15016 7200 15068 7206
rect 15068 7148 15240 7154
rect 15016 7142 15240 7148
rect 15028 7126 15240 7142
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 14844 6186 14872 6598
rect 15120 6322 15148 6598
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13636 4684 13688 4690
rect 13740 4672 13768 5102
rect 13924 4758 13952 5102
rect 14660 5098 14688 6122
rect 14740 6112 14792 6118
rect 15212 6089 15240 7126
rect 15396 6798 15424 7239
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15396 6118 15424 6734
rect 15488 6458 15516 6870
rect 15580 6798 15608 7142
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15384 6112 15436 6118
rect 14740 6054 14792 6060
rect 15198 6080 15254 6089
rect 14752 5846 14780 6054
rect 15384 6054 15436 6060
rect 15198 6015 15254 6024
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 15580 5710 15608 6734
rect 16394 6216 16450 6225
rect 15660 6180 15712 6186
rect 16394 6151 16450 6160
rect 15660 6122 15712 6128
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14936 5166 14964 5510
rect 15672 5370 15700 6122
rect 15752 5704 15804 5710
rect 15750 5672 15752 5681
rect 15804 5672 15806 5681
rect 15750 5607 15806 5616
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15106 5128 15162 5137
rect 14648 5092 14700 5098
rect 15106 5063 15108 5072
rect 14648 5034 14700 5040
rect 15160 5063 15162 5072
rect 15292 5092 15344 5098
rect 15108 5034 15160 5040
rect 15292 5034 15344 5040
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 13688 4644 13768 4672
rect 13636 4626 13688 4632
rect 13648 4078 13676 4626
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13174 3632 13230 3641
rect 13174 3567 13230 3576
rect 13648 3398 13676 4014
rect 13636 3392 13688 3398
rect 14200 3369 14228 4422
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14660 3720 14688 3878
rect 14568 3692 14688 3720
rect 14278 3632 14334 3641
rect 14278 3567 14280 3576
rect 14332 3567 14334 3576
rect 14280 3538 14332 3544
rect 13636 3334 13688 3340
rect 14186 3360 14242 3369
rect 13004 2774 13216 2802
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13188 1329 13216 2774
rect 13648 2417 13676 3334
rect 14186 3295 14242 3304
rect 14292 3194 14320 3538
rect 14568 3534 14596 3692
rect 15304 3670 15332 5034
rect 15764 4826 15792 5306
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15488 4321 15516 4626
rect 15566 4584 15622 4593
rect 15566 4519 15622 4528
rect 15474 4312 15530 4321
rect 15474 4247 15476 4256
rect 15528 4247 15530 4256
rect 15476 4218 15528 4224
rect 15488 4078 15516 4218
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14568 3194 14596 3470
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14280 3188 14332 3194
rect 14200 3148 14280 3176
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13818 2952 13874 2961
rect 13740 2650 13768 2926
rect 13818 2887 13874 2896
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13726 2544 13782 2553
rect 13726 2479 13728 2488
rect 13780 2479 13782 2488
rect 13728 2450 13780 2456
rect 13634 2408 13690 2417
rect 13634 2343 13690 2352
rect 13832 2310 13860 2887
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 13924 2514 13952 2586
rect 14016 2553 14044 3062
rect 14002 2544 14058 2553
rect 13912 2508 13964 2514
rect 14002 2479 14058 2488
rect 13912 2450 13964 2456
rect 14200 2446 14228 3148
rect 14280 3130 14332 3136
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14936 2922 14964 3334
rect 15304 3194 15332 3606
rect 15396 3505 15424 3878
rect 15488 3738 15516 4014
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15382 3496 15438 3505
rect 15580 3466 15608 4519
rect 16040 4486 16068 4694
rect 16028 4480 16080 4486
rect 16026 4448 16028 4457
rect 16080 4448 16082 4457
rect 16026 4383 16082 4392
rect 16408 4185 16436 6151
rect 16592 6118 16620 6802
rect 16580 6112 16632 6118
rect 16500 6060 16580 6066
rect 16500 6054 16632 6060
rect 16500 6038 16620 6054
rect 16394 4176 16450 4185
rect 16394 4111 16450 4120
rect 16500 3670 16528 6038
rect 16684 5710 16712 7278
rect 17236 7177 17264 7647
rect 17222 7168 17278 7177
rect 17222 7103 17278 7112
rect 18234 6896 18290 6905
rect 18234 6831 18236 6840
rect 18288 6831 18290 6840
rect 18236 6802 18288 6808
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17052 5778 17080 6598
rect 18248 6458 18276 6802
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18616 6458 18644 6734
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 17498 6352 17554 6361
rect 17498 6287 17500 6296
rect 17552 6287 17554 6296
rect 17500 6258 17552 6264
rect 18420 6248 18472 6254
rect 18418 6216 18420 6225
rect 18472 6216 18474 6225
rect 18418 6151 18474 6160
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15382 3431 15384 3440
rect 15436 3431 15438 3440
rect 15568 3460 15620 3466
rect 15384 3402 15436 3408
rect 15568 3402 15620 3408
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 14936 2650 14964 2858
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14936 2378 14964 2586
rect 15120 2514 15148 2858
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15304 2446 15332 3130
rect 15396 3058 15424 3402
rect 15580 3194 15608 3402
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15672 2650 15700 3470
rect 16592 2990 16620 5102
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16684 3369 16712 4014
rect 16776 4010 16804 4558
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16776 3738 16804 3946
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16670 3360 16726 3369
rect 16670 3295 16726 3304
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15658 2408 15714 2417
rect 14924 2372 14976 2378
rect 15658 2343 15660 2352
rect 14924 2314 14976 2320
rect 15712 2343 15714 2352
rect 15660 2314 15712 2320
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13174 1320 13230 1329
rect 13174 1255 13230 1264
rect 16316 480 16344 2926
rect 16868 2582 16896 5510
rect 17052 5370 17080 5714
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 17052 5250 17080 5306
rect 17052 5222 17172 5250
rect 17040 5092 17092 5098
rect 17040 5034 17092 5040
rect 17052 4865 17080 5034
rect 17038 4856 17094 4865
rect 17038 4791 17094 4800
rect 17144 4758 17172 5222
rect 17788 5137 17816 5782
rect 17880 5658 17908 6054
rect 17880 5630 18000 5658
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17774 5128 17830 5137
rect 17774 5063 17776 5072
rect 17828 5063 17830 5072
rect 17776 5034 17828 5040
rect 17788 5003 17816 5034
rect 17682 4992 17738 5001
rect 17682 4927 17738 4936
rect 17696 4758 17724 4927
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 17040 4072 17092 4078
rect 17144 4060 17172 4694
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17328 4214 17356 4626
rect 17316 4208 17368 4214
rect 17316 4150 17368 4156
rect 17092 4032 17172 4060
rect 17040 4014 17092 4020
rect 17144 3534 17172 4032
rect 17880 3942 17908 5510
rect 17972 5166 18000 5630
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17972 4146 18000 5102
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18156 4826 18184 5034
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17420 3602 17448 3878
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17130 3224 17186 3233
rect 17130 3159 17132 3168
rect 17184 3159 17186 3168
rect 17132 3130 17184 3136
rect 17420 2990 17448 3538
rect 17972 3194 18000 3538
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 18156 2650 18184 4762
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18524 4078 18552 4626
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18340 3369 18368 3538
rect 18326 3360 18382 3369
rect 18326 3295 18382 3304
rect 18524 3194 18552 4014
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18708 2854 18736 6598
rect 18892 6254 18920 9415
rect 23294 9072 23350 9081
rect 23294 9007 23350 9016
rect 20074 8936 20130 8945
rect 20074 8871 20130 8880
rect 19982 8256 20038 8265
rect 19982 8191 20038 8200
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19168 7546 19196 7890
rect 19890 7848 19946 7857
rect 19890 7783 19946 7792
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 18984 6730 19012 7142
rect 19076 7041 19104 7278
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19062 7032 19118 7041
rect 19062 6967 19118 6976
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 18984 6322 19012 6666
rect 19076 6662 19104 6802
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18880 6248 18932 6254
rect 19076 6202 19104 6598
rect 19260 6225 19288 7142
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 18880 6190 18932 6196
rect 18984 6174 19104 6202
rect 19246 6216 19302 6225
rect 18984 6118 19012 6174
rect 19246 6151 19302 6160
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18984 5370 19012 6054
rect 19352 5846 19380 6598
rect 19708 6180 19760 6186
rect 19708 6122 19760 6128
rect 19720 5846 19748 6122
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 19708 5840 19760 5846
rect 19708 5782 19760 5788
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 19812 5250 19840 7482
rect 19904 7342 19932 7783
rect 19996 7342 20024 8191
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19904 5642 19932 6666
rect 19892 5636 19944 5642
rect 19892 5578 19944 5584
rect 19812 5222 19932 5250
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19352 4690 19380 4966
rect 19812 4758 19840 5102
rect 19800 4752 19852 4758
rect 19800 4694 19852 4700
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 18800 4078 18828 4626
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 18800 3738 18828 4014
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18892 2990 18920 4014
rect 19260 3602 19288 4014
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19260 2990 19288 3538
rect 19352 3369 19380 4626
rect 19720 4078 19748 4626
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19904 3641 19932 5222
rect 20088 4690 20116 8871
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20180 6662 20208 7142
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20364 4078 20392 5510
rect 20456 4146 20484 7686
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20732 6118 20760 6802
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20824 6322 20852 6734
rect 20916 6730 20944 7142
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20628 5636 20680 5642
rect 20628 5578 20680 5584
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20364 3670 20392 4014
rect 20640 3670 20668 5578
rect 20732 5370 20760 6054
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20824 4758 20852 6258
rect 21086 6216 21142 6225
rect 21284 6202 21312 6394
rect 21560 6390 21588 6666
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21142 6174 21312 6202
rect 21086 6151 21088 6160
rect 21140 6151 21142 6160
rect 21088 6122 21140 6128
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 21284 5098 21312 5782
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21272 5092 21324 5098
rect 21272 5034 21324 5040
rect 21376 5030 21404 5646
rect 21560 5302 21588 6326
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 20904 5024 20956 5030
rect 21364 5024 21416 5030
rect 20904 4966 20956 4972
rect 21362 4992 21364 5001
rect 21652 5001 21680 7278
rect 23020 7268 23072 7274
rect 23020 7210 23072 7216
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21824 5568 21876 5574
rect 21824 5510 21876 5516
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21416 4992 21418 5001
rect 20812 4752 20864 4758
rect 20812 4694 20864 4700
rect 20916 4570 20944 4966
rect 21362 4927 21418 4936
rect 21638 4992 21694 5001
rect 21638 4927 21694 4936
rect 21362 4856 21418 4865
rect 21272 4820 21324 4826
rect 21362 4791 21418 4800
rect 21272 4762 21324 4768
rect 20824 4542 20944 4570
rect 20824 4010 20852 4542
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20824 3913 20852 3946
rect 20810 3904 20866 3913
rect 20810 3839 20866 3848
rect 21284 3670 21312 4762
rect 21376 4758 21404 4791
rect 21364 4752 21416 4758
rect 21364 4694 21416 4700
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 21468 4010 21496 4626
rect 21652 4593 21680 4927
rect 21638 4584 21694 4593
rect 21638 4519 21694 4528
rect 21744 4282 21772 5034
rect 21836 4826 21864 5510
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 21928 4622 21956 7142
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22756 5846 22784 6054
rect 22744 5840 22796 5846
rect 22744 5782 22796 5788
rect 22836 5840 22888 5846
rect 22836 5782 22888 5788
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22112 5114 22140 5510
rect 22848 5370 22876 5782
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22020 5098 22140 5114
rect 22008 5092 22140 5098
rect 22060 5086 22140 5092
rect 22008 5034 22060 5040
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 21732 4276 21784 4282
rect 21732 4218 21784 4224
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 20352 3664 20404 3670
rect 19890 3632 19946 3641
rect 19890 3567 19946 3576
rect 20258 3632 20314 3641
rect 20352 3606 20404 3612
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 21272 3664 21324 3670
rect 21272 3606 21324 3612
rect 20258 3567 20314 3576
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19338 3360 19394 3369
rect 19338 3295 19394 3304
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 17406 2544 17462 2553
rect 18340 2514 18368 2790
rect 19352 2650 19380 3295
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19536 2582 19564 2858
rect 19524 2576 19576 2582
rect 19524 2518 19576 2524
rect 17406 2479 17408 2488
rect 17460 2479 17462 2488
rect 18328 2508 18380 2514
rect 17408 2450 17460 2456
rect 18328 2450 18380 2456
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16776 2145 16804 2382
rect 19812 2145 19840 3470
rect 16762 2136 16818 2145
rect 16762 2071 16818 2080
rect 19798 2136 19854 2145
rect 19798 2071 19854 2080
rect 19904 480 19932 3567
rect 20272 2650 20300 3567
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20074 2544 20130 2553
rect 20548 2514 20576 3402
rect 20824 3398 20852 3429
rect 20628 3392 20680 3398
rect 20812 3392 20864 3398
rect 20628 3334 20680 3340
rect 20810 3360 20812 3369
rect 20864 3360 20866 3369
rect 20640 2904 20668 3334
rect 20810 3295 20866 3304
rect 20824 3194 20852 3295
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 21652 2990 21680 4082
rect 21928 3738 21956 4558
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22020 4060 22048 4422
rect 22100 4072 22152 4078
rect 22020 4032 22100 4060
rect 22152 4032 22232 4060
rect 22100 4014 22152 4020
rect 22112 3949 22140 4014
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21928 2990 21956 3674
rect 22204 3097 22232 4032
rect 22296 3466 22324 5170
rect 22742 4992 22798 5001
rect 22742 4927 22798 4936
rect 22466 4856 22522 4865
rect 22466 4791 22522 4800
rect 22376 4684 22428 4690
rect 22376 4626 22428 4632
rect 22388 4486 22416 4626
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22388 4146 22416 4422
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22388 3738 22416 4082
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 22190 3088 22246 3097
rect 22388 3058 22416 3334
rect 22190 3023 22246 3032
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22480 2990 22508 4791
rect 22756 4690 22784 4927
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22756 4282 22784 4626
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22650 4040 22706 4049
rect 22650 3975 22706 3984
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 21640 2984 21692 2990
rect 21560 2944 21640 2972
rect 20720 2916 20772 2922
rect 20640 2876 20720 2904
rect 20640 2650 20668 2876
rect 20720 2858 20772 2864
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 21560 2514 21588 2944
rect 21640 2926 21692 2932
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22112 2514 22140 2926
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22388 2514 22416 2858
rect 22480 2553 22508 2926
rect 22572 2922 22600 3878
rect 22664 3126 22692 3975
rect 22756 3602 22784 4218
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 22836 4004 22888 4010
rect 22836 3946 22888 3952
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22756 3194 22784 3538
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 22652 3120 22704 3126
rect 22848 3097 22876 3946
rect 22652 3062 22704 3068
rect 22834 3088 22890 3097
rect 22834 3023 22890 3032
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 22466 2544 22522 2553
rect 20074 2479 20076 2488
rect 20128 2479 20130 2488
rect 20536 2508 20588 2514
rect 20076 2450 20128 2456
rect 20536 2450 20588 2456
rect 21548 2508 21600 2514
rect 21548 2450 21600 2456
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 22376 2508 22428 2514
rect 22940 2514 22968 4082
rect 22466 2479 22522 2488
rect 22928 2508 22980 2514
rect 22376 2450 22428 2456
rect 22928 2450 22980 2456
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 23032 1601 23060 7210
rect 23308 7177 23336 9007
rect 23294 7168 23350 7177
rect 23294 7103 23350 7112
rect 23308 6458 23336 7103
rect 23400 7002 23428 10639
rect 29734 10432 29790 10441
rect 27622 10364 27918 10384
rect 29734 10367 29790 10376
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 28814 9616 28870 9625
rect 28814 9551 28870 9560
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 24766 8528 24822 8537
rect 24766 8463 24822 8472
rect 24674 8392 24730 8401
rect 24674 8327 24730 8336
rect 24688 7313 24716 8327
rect 24780 7449 24808 8463
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 24766 7440 24822 7449
rect 24766 7375 24822 7384
rect 24214 7304 24270 7313
rect 24214 7239 24270 7248
rect 24674 7304 24730 7313
rect 24674 7239 24730 7248
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23492 6186 23520 6802
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 24044 5710 24072 6054
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 23388 5568 23440 5574
rect 23388 5510 23440 5516
rect 23400 5234 23428 5510
rect 24228 5370 24256 7239
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24504 6458 24532 6802
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24596 5846 24624 6598
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 24492 5704 24544 5710
rect 24492 5646 24544 5652
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 24228 5166 24256 5306
rect 24216 5160 24268 5166
rect 24216 5102 24268 5108
rect 23296 5024 23348 5030
rect 23296 4966 23348 4972
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23308 4690 23336 4966
rect 23492 4826 23520 4966
rect 24504 4826 24532 5646
rect 24596 5370 24624 5782
rect 24584 5364 24636 5370
rect 24584 5306 24636 5312
rect 24688 5030 24716 6394
rect 24872 6322 24900 6598
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24872 6202 24900 6258
rect 24780 6174 24900 6202
rect 25240 6186 25268 6326
rect 25412 6316 25464 6322
rect 25412 6258 25464 6264
rect 25228 6180 25280 6186
rect 24780 5302 24808 6174
rect 25228 6122 25280 6128
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25056 5642 25084 6054
rect 25240 5778 25268 6122
rect 25318 6080 25374 6089
rect 25318 6015 25374 6024
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25044 5636 25096 5642
rect 25044 5578 25096 5584
rect 24952 5568 25004 5574
rect 24952 5510 25004 5516
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24768 5092 24820 5098
rect 24964 5080 24992 5510
rect 25056 5234 25084 5578
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 24820 5052 24992 5080
rect 24768 5034 24820 5040
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 24492 4820 24544 4826
rect 24492 4762 24544 4768
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23308 3942 23336 4626
rect 23492 4146 23520 4762
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 23584 4214 23612 4626
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 23572 4208 23624 4214
rect 23572 4150 23624 4156
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23296 3936 23348 3942
rect 23480 3936 23532 3942
rect 23296 3878 23348 3884
rect 23478 3904 23480 3913
rect 23532 3904 23534 3913
rect 23308 3602 23336 3878
rect 23478 3839 23534 3848
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 23756 3596 23808 3602
rect 23756 3538 23808 3544
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23492 2922 23520 3334
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23480 2916 23532 2922
rect 23480 2858 23532 2864
rect 23110 2680 23166 2689
rect 23110 2615 23166 2624
rect 23124 2582 23152 2615
rect 23112 2576 23164 2582
rect 23112 2518 23164 2524
rect 23492 2514 23520 2858
rect 23480 2508 23532 2514
rect 23480 2450 23532 2456
rect 23018 1592 23074 1601
rect 23018 1527 23074 1536
rect 23584 480 23612 3130
rect 23768 3058 23796 3538
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 24136 2990 24164 4558
rect 24688 4078 24716 4966
rect 24860 4752 24912 4758
rect 24860 4694 24912 4700
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24780 4010 24808 4558
rect 24768 4004 24820 4010
rect 24768 3946 24820 3952
rect 24780 3670 24808 3946
rect 24872 3942 24900 4694
rect 24860 3936 24912 3942
rect 24860 3878 24912 3884
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24596 2990 24624 3334
rect 24872 3126 24900 3878
rect 24964 3534 24992 5052
rect 25240 4826 25268 5714
rect 25228 4820 25280 4826
rect 25228 4762 25280 4768
rect 25332 4078 25360 6015
rect 25424 5574 25452 6258
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 27252 5772 27304 5778
rect 27252 5714 27304 5720
rect 26148 5704 26200 5710
rect 26148 5646 26200 5652
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25320 4072 25372 4078
rect 25320 4014 25372 4020
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25412 3664 25464 3670
rect 25412 3606 25464 3612
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 25424 3194 25452 3606
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 24584 2984 24636 2990
rect 24584 2926 24636 2932
rect 24136 2514 24164 2926
rect 25042 2544 25098 2553
rect 24124 2508 24176 2514
rect 25042 2479 25044 2488
rect 24124 2450 24176 2456
rect 25096 2479 25098 2488
rect 25044 2450 25096 2456
rect 25516 1329 25544 4014
rect 25872 3936 25924 3942
rect 25872 3878 25924 3884
rect 25884 3738 25912 3878
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 26160 3670 26188 5646
rect 26882 5536 26938 5545
rect 26882 5471 26938 5480
rect 26330 5264 26386 5273
rect 26330 5199 26386 5208
rect 26344 5166 26372 5199
rect 26896 5166 26924 5471
rect 27264 5370 27292 5714
rect 27988 5704 28040 5710
rect 27988 5646 28040 5652
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27632 5250 27660 5510
rect 27540 5234 27660 5250
rect 27528 5228 27660 5234
rect 27580 5222 27660 5228
rect 27528 5170 27580 5176
rect 26332 5160 26384 5166
rect 26332 5102 26384 5108
rect 26884 5160 26936 5166
rect 26884 5102 26936 5108
rect 26792 5024 26844 5030
rect 26792 4966 26844 4972
rect 26804 4758 26832 4966
rect 27540 4826 27568 5170
rect 28000 5098 28028 5646
rect 28828 5250 28856 9551
rect 28906 5264 28962 5273
rect 28828 5222 28906 5250
rect 28906 5199 28962 5208
rect 29000 5160 29052 5166
rect 29000 5102 29052 5108
rect 27988 5092 28040 5098
rect 27988 5034 28040 5040
rect 28264 5092 28316 5098
rect 28264 5034 28316 5040
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 26792 4752 26844 4758
rect 26606 4720 26662 4729
rect 26792 4694 26844 4700
rect 27620 4752 27672 4758
rect 27620 4694 27672 4700
rect 27712 4752 27764 4758
rect 27712 4694 27764 4700
rect 26606 4655 26608 4664
rect 26660 4655 26662 4664
rect 26608 4626 26660 4632
rect 26516 4548 26568 4554
rect 26516 4490 26568 4496
rect 26528 4078 26556 4490
rect 26620 4282 26648 4626
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26608 4276 26660 4282
rect 26608 4218 26660 4224
rect 26516 4072 26568 4078
rect 26514 4040 26516 4049
rect 26568 4040 26570 4049
rect 26804 4010 26832 4422
rect 27632 4282 27660 4694
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27724 4010 27752 4694
rect 26514 3975 26570 3984
rect 26792 4004 26844 4010
rect 26792 3946 26844 3952
rect 27712 4004 27764 4010
rect 27712 3946 27764 3952
rect 26804 3670 26832 3946
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 26148 3664 26200 3670
rect 26148 3606 26200 3612
rect 26332 3664 26384 3670
rect 26332 3606 26384 3612
rect 26792 3664 26844 3670
rect 26792 3606 26844 3612
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26252 3058 26280 3334
rect 26344 3126 26372 3606
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26332 3120 26384 3126
rect 26332 3062 26384 3068
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 26252 2689 26280 2994
rect 26344 2922 26372 3062
rect 26436 2990 26464 3470
rect 27436 3392 27488 3398
rect 27434 3360 27436 3369
rect 28000 3369 28028 5034
rect 28276 4758 28304 5034
rect 28264 4752 28316 4758
rect 29012 4729 29040 5102
rect 28264 4694 28316 4700
rect 28998 4720 29054 4729
rect 28276 3738 28304 4694
rect 28998 4655 29054 4664
rect 29184 4684 29236 4690
rect 29184 4626 29236 4632
rect 29196 4282 29224 4626
rect 29552 4480 29604 4486
rect 29552 4422 29604 4428
rect 29184 4276 29236 4282
rect 29184 4218 29236 4224
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 29104 3777 29132 4014
rect 29090 3768 29146 3777
rect 28264 3732 28316 3738
rect 29090 3703 29146 3712
rect 28264 3674 28316 3680
rect 29196 3670 29224 4218
rect 29276 3936 29328 3942
rect 29276 3878 29328 3884
rect 28540 3664 28592 3670
rect 28540 3606 28592 3612
rect 29184 3664 29236 3670
rect 29184 3606 29236 3612
rect 27488 3360 27490 3369
rect 27434 3295 27490 3304
rect 27986 3360 28042 3369
rect 27986 3295 28042 3304
rect 28552 3194 28580 3606
rect 28908 3460 28960 3466
rect 28908 3402 28960 3408
rect 28540 3188 28592 3194
rect 28540 3130 28592 3136
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26332 2916 26384 2922
rect 26332 2858 26384 2864
rect 26238 2680 26294 2689
rect 26238 2615 26294 2624
rect 26344 2582 26372 2858
rect 27436 2848 27488 2854
rect 27436 2790 27488 2796
rect 26332 2576 26384 2582
rect 26332 2518 26384 2524
rect 27160 2576 27212 2582
rect 27160 2518 27212 2524
rect 25502 1320 25558 1329
rect 25502 1255 25558 1264
rect 27172 480 27200 2518
rect 27448 2514 27476 2790
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 27620 2576 27672 2582
rect 27618 2544 27620 2553
rect 27672 2544 27674 2553
rect 27436 2508 27488 2514
rect 27618 2479 27674 2488
rect 27802 2544 27858 2553
rect 28920 2514 28948 3402
rect 29090 3360 29146 3369
rect 29090 3295 29146 3304
rect 29104 2990 29132 3295
rect 29288 3058 29316 3878
rect 29276 3052 29328 3058
rect 29276 2994 29328 3000
rect 29000 2984 29052 2990
rect 29000 2926 29052 2932
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29012 2650 29040 2926
rect 29564 2650 29592 4422
rect 29748 4078 29776 10367
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34978 7848 35034 7857
rect 34978 7783 35034 7792
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 34992 7342 35020 7783
rect 34980 7336 35032 7342
rect 34980 7278 35032 7284
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 33782 5536 33838 5545
rect 33782 5471 33838 5480
rect 30654 5264 30710 5273
rect 30654 5199 30710 5208
rect 30668 4690 30696 5199
rect 33796 4865 33824 5471
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 35084 5370 35112 12815
rect 35268 6730 35296 13767
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 35452 10470 35480 11154
rect 35440 10464 35492 10470
rect 35438 10432 35440 10441
rect 35492 10432 35494 10441
rect 35438 10367 35494 10376
rect 35440 10124 35492 10130
rect 35440 10066 35492 10072
rect 35452 9518 35480 10066
rect 35440 9512 35492 9518
rect 35438 9480 35440 9489
rect 35492 9480 35494 9489
rect 35438 9415 35494 9424
rect 35438 9072 35494 9081
rect 35438 9007 35440 9016
rect 35492 9007 35494 9016
rect 35440 8978 35492 8984
rect 35452 8634 35480 8978
rect 35440 8628 35492 8634
rect 35440 8570 35492 8576
rect 35438 8528 35494 8537
rect 35438 8463 35494 8472
rect 35452 8430 35480 8463
rect 35440 8424 35492 8430
rect 35440 8366 35492 8372
rect 35544 8090 35572 15535
rect 35806 14648 35862 14657
rect 35806 14583 35862 14592
rect 35622 12064 35678 12073
rect 35622 11999 35678 12008
rect 35636 11354 35664 11999
rect 35624 11348 35676 11354
rect 35624 11290 35676 11296
rect 35622 11112 35678 11121
rect 35622 11047 35678 11056
rect 35636 10266 35664 11047
rect 35714 10296 35770 10305
rect 35624 10260 35676 10266
rect 35714 10231 35770 10240
rect 35624 10202 35676 10208
rect 35622 9344 35678 9353
rect 35622 9279 35678 9288
rect 35636 8634 35664 9279
rect 35728 9178 35756 10231
rect 35716 9172 35768 9178
rect 35716 9114 35768 9120
rect 35624 8628 35676 8634
rect 35624 8570 35676 8576
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35438 7984 35494 7993
rect 35438 7919 35440 7928
rect 35492 7919 35494 7928
rect 35440 7890 35492 7896
rect 35452 7546 35480 7890
rect 35820 7546 35848 14583
rect 36726 8528 36782 8537
rect 36726 8463 36782 8472
rect 36542 8256 36598 8265
rect 36542 8191 36598 8200
rect 35440 7540 35492 7546
rect 35440 7482 35492 7488
rect 35808 7540 35860 7546
rect 35808 7482 35860 7488
rect 36556 7342 36584 8191
rect 36740 7546 36768 8463
rect 36728 7540 36780 7546
rect 36728 7482 36780 7488
rect 36544 7336 36596 7342
rect 36544 7278 36596 7284
rect 35440 6860 35492 6866
rect 35440 6802 35492 6808
rect 35256 6724 35308 6730
rect 35256 6666 35308 6672
rect 35452 6390 35480 6802
rect 35440 6384 35492 6390
rect 35438 6352 35440 6361
rect 35492 6352 35494 6361
rect 35438 6287 35494 6296
rect 35072 5364 35124 5370
rect 35072 5306 35124 5312
rect 33782 4856 33838 4865
rect 33782 4791 33838 4800
rect 30656 4684 30708 4690
rect 30656 4626 30708 4632
rect 30564 4480 30616 4486
rect 30564 4422 30616 4428
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 30484 4010 30512 4082
rect 30380 4004 30432 4010
rect 30380 3946 30432 3952
rect 30472 4004 30524 4010
rect 30472 3946 30524 3952
rect 30392 3738 30420 3946
rect 30484 3738 30512 3946
rect 30380 3732 30432 3738
rect 30380 3674 30432 3680
rect 30472 3732 30524 3738
rect 30472 3674 30524 3680
rect 30576 3670 30604 4422
rect 30668 4282 30696 4626
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 30656 4276 30708 4282
rect 30656 4218 30708 4224
rect 31300 4276 31352 4282
rect 31300 4218 31352 4224
rect 31312 4185 31340 4218
rect 31298 4176 31354 4185
rect 31298 4111 31354 4120
rect 31024 4004 31076 4010
rect 31024 3946 31076 3952
rect 30564 3664 30616 3670
rect 30564 3606 30616 3612
rect 30656 3664 30708 3670
rect 30656 3606 30708 3612
rect 30838 3632 30894 3641
rect 30668 3194 30696 3606
rect 30838 3567 30894 3576
rect 30656 3188 30708 3194
rect 30656 3130 30708 3136
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 27802 2479 27804 2488
rect 27436 2450 27488 2456
rect 27856 2479 27858 2488
rect 28908 2508 28960 2514
rect 27804 2450 27856 2456
rect 28908 2450 28960 2456
rect 28906 2408 28962 2417
rect 28906 2343 28908 2352
rect 28960 2343 28962 2352
rect 28908 2314 28960 2320
rect 30852 480 30880 3567
rect 31036 3534 31064 3946
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31036 3210 31064 3470
rect 31036 3182 31248 3210
rect 32232 3194 32260 3538
rect 32496 3392 32548 3398
rect 32496 3334 32548 3340
rect 31220 2922 31248 3182
rect 32220 3188 32272 3194
rect 32220 3130 32272 3136
rect 32508 3058 32536 3334
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 32036 3052 32088 3058
rect 32036 2994 32088 3000
rect 32496 3052 32548 3058
rect 32496 2994 32548 3000
rect 30932 2916 30984 2922
rect 30932 2858 30984 2864
rect 31208 2916 31260 2922
rect 31208 2858 31260 2864
rect 30944 2650 30972 2858
rect 31312 2650 31340 2994
rect 31666 2816 31722 2825
rect 31666 2751 31722 2760
rect 31680 2650 31708 2751
rect 32048 2650 32076 2994
rect 32588 2916 32640 2922
rect 32588 2858 32640 2864
rect 30932 2644 30984 2650
rect 30932 2586 30984 2592
rect 31300 2644 31352 2650
rect 31300 2586 31352 2592
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 32036 2644 32088 2650
rect 32036 2586 32088 2592
rect 30944 2446 30972 2586
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 31312 2378 31340 2586
rect 32600 2582 32628 2858
rect 34150 2816 34206 2825
rect 34150 2751 34206 2760
rect 32588 2576 32640 2582
rect 32586 2544 32588 2553
rect 32640 2544 32642 2553
rect 32586 2479 32642 2488
rect 31300 2372 31352 2378
rect 31300 2314 31352 2320
rect 34164 1442 34192 2751
rect 38106 2408 38162 2417
rect 38106 2343 38162 2352
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 34164 1414 34468 1442
rect 34440 480 34468 1414
rect 38120 480 38148 2343
rect 4250 232 4306 241
rect 4250 167 4306 176
rect 5354 0 5410 480
rect 9034 0 9090 480
rect 12622 0 12678 480
rect 16302 0 16358 480
rect 19338 96 19394 105
rect 19338 31 19340 40
rect 19392 31 19394 40
rect 19340 2 19392 8
rect 19890 0 19946 480
rect 23570 0 23626 480
rect 27158 0 27214 480
rect 28906 96 28962 105
rect 28906 31 28908 40
rect 28960 31 28962 40
rect 28908 2 28960 8
rect 30838 0 30894 480
rect 34426 0 34482 480
rect 38106 0 38162 480
<< via2 >>
rect 1766 15544 1822 15600
rect 1490 12824 1546 12880
rect 1582 12008 1638 12064
rect 1582 11056 1638 11112
rect 1490 10240 1546 10296
rect 1582 9288 1638 9344
rect 1674 8880 1730 8936
rect 35530 15544 35586 15600
rect 1858 14592 1914 14648
rect 1950 13776 2006 13832
rect 2042 9036 2098 9072
rect 3422 9560 3478 9616
rect 2042 9016 2044 9036
rect 2044 9016 2096 9036
rect 2096 9016 2098 9036
rect 2502 8472 2558 8528
rect 2042 7792 2098 7848
rect 5078 8492 5134 8528
rect 5078 8472 5080 8492
rect 5080 8472 5132 8492
rect 5132 8472 5134 8492
rect 2686 8064 2742 8120
rect 2594 7520 2650 7576
rect 2042 5888 2098 5944
rect 2042 5228 2098 5264
rect 2042 5208 2044 5228
rect 2044 5208 2096 5228
rect 2096 5208 2098 5228
rect 2778 3984 2834 4040
rect 2778 3712 2834 3768
rect 1766 2352 1822 2408
rect 3054 8200 3110 8256
rect 5078 8084 5134 8120
rect 5078 8064 5080 8084
rect 5080 8064 5132 8084
rect 5132 8064 5134 8084
rect 3974 7656 4030 7712
rect 3422 3848 3478 3904
rect 2962 3440 3018 3496
rect 4342 7520 4398 7576
rect 3606 4528 3662 4584
rect 5630 8064 5686 8120
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 16670 11600 16726 11656
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 12990 9016 13046 9072
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 12990 8336 13046 8392
rect 5630 7656 5686 7712
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 6826 7384 6882 7440
rect 3974 4120 4030 4176
rect 6826 6568 6882 6624
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 10690 7656 10746 7712
rect 3974 3032 4030 3088
rect 2870 448 2926 504
rect 5906 6160 5962 6216
rect 7194 6160 7250 6216
rect 5262 3848 5318 3904
rect 6458 3884 6460 3904
rect 6460 3884 6512 3904
rect 6512 3884 6514 3904
rect 6458 3848 6514 3884
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 7010 2932 7012 2952
rect 7012 2932 7064 2952
rect 7064 2932 7066 2952
rect 7010 2896 7066 2932
rect 5538 2796 5540 2816
rect 5540 2796 5592 2816
rect 5592 2796 5594 2816
rect 5538 2760 5594 2796
rect 9862 6160 9918 6216
rect 9862 5888 9918 5944
rect 10598 4936 10654 4992
rect 10138 4528 10194 4584
rect 9126 3884 9128 3904
rect 9128 3884 9180 3904
rect 9180 3884 9182 3904
rect 9126 3848 9182 3884
rect 9126 3576 9182 3632
rect 8758 3440 8814 3496
rect 8850 3304 8906 3360
rect 8666 2760 8722 2816
rect 9310 3168 9366 3224
rect 10230 3712 10286 3768
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14186 7520 14242 7576
rect 14370 7540 14426 7576
rect 14370 7520 14372 7540
rect 14372 7520 14424 7540
rect 14424 7520 14426 7540
rect 11334 6604 11336 6624
rect 11336 6604 11388 6624
rect 11388 6604 11390 6624
rect 11334 6568 11390 6604
rect 11150 5752 11206 5808
rect 12254 3576 12310 3632
rect 11058 3460 11114 3496
rect 11058 3440 11060 3460
rect 11060 3440 11112 3460
rect 11112 3440 11114 3460
rect 11518 3052 11574 3088
rect 11518 3032 11520 3052
rect 11520 3032 11572 3052
rect 11572 3032 11574 3052
rect 11886 3168 11942 3224
rect 12530 4936 12586 4992
rect 13726 7268 13782 7304
rect 13726 7248 13728 7268
rect 13728 7248 13780 7268
rect 13780 7248 13782 7268
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 35254 13776 35310 13832
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 35070 12824 35126 12880
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 33322 11600 33378 11656
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 19982 10648 20038 10704
rect 23386 10648 23442 10704
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 18878 9424 18934 9480
rect 17222 7656 17278 7712
rect 15382 7248 15438 7304
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14002 6568 14058 6624
rect 12806 4392 12862 4448
rect 12530 4256 12586 4312
rect 12530 3732 12586 3768
rect 12530 3712 12532 3732
rect 12532 3712 12584 3732
rect 12584 3712 12586 3732
rect 10690 2624 10746 2680
rect 12254 2760 12310 2816
rect 11426 2524 11428 2544
rect 11428 2524 11480 2544
rect 11480 2524 11482 2544
rect 11426 2488 11482 2524
rect 10506 2372 10562 2408
rect 10506 2352 10508 2372
rect 10508 2352 10560 2372
rect 10560 2352 10562 2372
rect 12070 2388 12072 2408
rect 12072 2388 12124 2408
rect 12124 2388 12126 2408
rect 12070 2352 12126 2388
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 15198 6024 15254 6080
rect 16394 6160 16450 6216
rect 15750 5652 15752 5672
rect 15752 5652 15804 5672
rect 15804 5652 15806 5672
rect 15750 5616 15806 5652
rect 15106 5092 15162 5128
rect 15106 5072 15108 5092
rect 15108 5072 15160 5092
rect 15160 5072 15162 5092
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 13174 3576 13230 3632
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14278 3596 14334 3632
rect 14278 3576 14280 3596
rect 14280 3576 14332 3596
rect 14332 3576 14334 3596
rect 14186 3304 14242 3360
rect 15566 4528 15622 4584
rect 15474 4276 15530 4312
rect 15474 4256 15476 4276
rect 15476 4256 15528 4276
rect 15528 4256 15530 4276
rect 13818 2896 13874 2952
rect 13726 2508 13782 2544
rect 13726 2488 13728 2508
rect 13728 2488 13780 2508
rect 13780 2488 13782 2508
rect 13634 2352 13690 2408
rect 14002 2488 14058 2544
rect 15382 3460 15438 3496
rect 16026 4428 16028 4448
rect 16028 4428 16080 4448
rect 16080 4428 16082 4448
rect 16026 4392 16082 4428
rect 16394 4120 16450 4176
rect 17222 7112 17278 7168
rect 18234 6860 18290 6896
rect 18234 6840 18236 6860
rect 18236 6840 18288 6860
rect 18288 6840 18290 6860
rect 17498 6316 17554 6352
rect 17498 6296 17500 6316
rect 17500 6296 17552 6316
rect 17552 6296 17554 6316
rect 18418 6196 18420 6216
rect 18420 6196 18472 6216
rect 18472 6196 18474 6216
rect 18418 6160 18474 6196
rect 15382 3440 15384 3460
rect 15384 3440 15436 3460
rect 15436 3440 15438 3460
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 16670 3304 16726 3360
rect 15658 2372 15714 2408
rect 15658 2352 15660 2372
rect 15660 2352 15712 2372
rect 15712 2352 15714 2372
rect 13174 1264 13230 1320
rect 17038 4800 17094 4856
rect 17774 5092 17830 5128
rect 17774 5072 17776 5092
rect 17776 5072 17828 5092
rect 17828 5072 17830 5092
rect 17682 4936 17738 4992
rect 17130 3188 17186 3224
rect 17130 3168 17132 3188
rect 17132 3168 17184 3188
rect 17184 3168 17186 3188
rect 18326 3304 18382 3360
rect 23294 9016 23350 9072
rect 20074 8880 20130 8936
rect 19982 8200 20038 8256
rect 19890 7792 19946 7848
rect 19062 6976 19118 7032
rect 19246 6160 19302 6216
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 21086 6180 21142 6216
rect 21086 6160 21088 6180
rect 21088 6160 21140 6180
rect 21140 6160 21142 6180
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 21362 4972 21364 4992
rect 21364 4972 21416 4992
rect 21416 4972 21418 4992
rect 21362 4936 21418 4972
rect 21638 4936 21694 4992
rect 21362 4800 21418 4856
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20810 3848 20866 3904
rect 21638 4528 21694 4584
rect 19890 3576 19946 3632
rect 20258 3576 20314 3632
rect 19338 3304 19394 3360
rect 17406 2508 17462 2544
rect 17406 2488 17408 2508
rect 17408 2488 17460 2508
rect 17460 2488 17462 2508
rect 16762 2080 16818 2136
rect 19798 2080 19854 2136
rect 20074 2508 20130 2544
rect 20810 3340 20812 3360
rect 20812 3340 20864 3360
rect 20864 3340 20866 3360
rect 20810 3304 20866 3340
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 22742 4936 22798 4992
rect 22466 4800 22522 4856
rect 22190 3032 22246 3088
rect 22650 3984 22706 4040
rect 22834 3032 22890 3088
rect 20074 2488 20076 2508
rect 20076 2488 20128 2508
rect 20128 2488 20130 2508
rect 22466 2488 22522 2544
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 23294 7112 23350 7168
rect 29734 10376 29790 10432
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 28814 9560 28870 9616
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 24766 8472 24822 8528
rect 24674 8336 24730 8392
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 24766 7384 24822 7440
rect 24214 7248 24270 7304
rect 24674 7248 24730 7304
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 25318 6024 25374 6080
rect 23478 3884 23480 3904
rect 23480 3884 23532 3904
rect 23532 3884 23534 3904
rect 23478 3848 23534 3884
rect 23110 2624 23166 2680
rect 23018 1536 23074 1592
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 25042 2508 25098 2544
rect 25042 2488 25044 2508
rect 25044 2488 25096 2508
rect 25096 2488 25098 2508
rect 26882 5480 26938 5536
rect 26330 5208 26386 5264
rect 28906 5208 28962 5264
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 26606 4684 26662 4720
rect 26606 4664 26608 4684
rect 26608 4664 26660 4684
rect 26660 4664 26662 4684
rect 26514 4020 26516 4040
rect 26516 4020 26568 4040
rect 26568 4020 26570 4040
rect 26514 3984 26570 4020
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 28998 4664 29054 4720
rect 29090 3712 29146 3768
rect 27434 3340 27436 3360
rect 27436 3340 27488 3360
rect 27488 3340 27490 3360
rect 27434 3304 27490 3340
rect 27986 3304 28042 3360
rect 26238 2624 26294 2680
rect 25502 1264 25558 1320
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 27618 2524 27620 2544
rect 27620 2524 27672 2544
rect 27672 2524 27674 2544
rect 27618 2488 27674 2524
rect 27802 2508 27858 2544
rect 29090 3304 29146 3360
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 34978 7792 35034 7848
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 33782 5480 33838 5536
rect 30654 5208 30710 5264
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 35438 10412 35440 10432
rect 35440 10412 35492 10432
rect 35492 10412 35494 10432
rect 35438 10376 35494 10412
rect 35438 9460 35440 9480
rect 35440 9460 35492 9480
rect 35492 9460 35494 9480
rect 35438 9424 35494 9460
rect 35438 9036 35494 9072
rect 35438 9016 35440 9036
rect 35440 9016 35492 9036
rect 35492 9016 35494 9036
rect 35438 8472 35494 8528
rect 35806 14592 35862 14648
rect 35622 12008 35678 12064
rect 35622 11056 35678 11112
rect 35714 10240 35770 10296
rect 35622 9288 35678 9344
rect 35438 7948 35494 7984
rect 35438 7928 35440 7948
rect 35440 7928 35492 7948
rect 35492 7928 35494 7948
rect 36726 8472 36782 8528
rect 36542 8200 36598 8256
rect 35438 6332 35440 6352
rect 35440 6332 35492 6352
rect 35492 6332 35494 6352
rect 35438 6296 35494 6332
rect 33782 4800 33838 4856
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 31298 4120 31354 4176
rect 30838 3576 30894 3632
rect 27802 2488 27804 2508
rect 27804 2488 27856 2508
rect 27856 2488 27858 2508
rect 28906 2372 28962 2408
rect 28906 2352 28908 2372
rect 28908 2352 28960 2372
rect 28960 2352 28962 2372
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 31666 2760 31722 2816
rect 34150 2760 34206 2816
rect 32586 2524 32588 2544
rect 32588 2524 32640 2544
rect 32640 2524 32642 2544
rect 32586 2488 32642 2524
rect 38106 2352 38162 2408
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 4250 176 4306 232
rect 19338 60 19394 96
rect 19338 40 19340 60
rect 19340 40 19392 60
rect 19392 40 19394 60
rect 28906 60 28962 96
rect 28906 40 28908 60
rect 28908 40 28960 60
rect 28960 40 28962 60
<< metal3 >>
rect 0 15602 480 15632
rect 1761 15602 1827 15605
rect 0 15600 1827 15602
rect 0 15544 1766 15600
rect 1822 15544 1827 15600
rect 0 15542 1827 15544
rect 0 15512 480 15542
rect 1761 15539 1827 15542
rect 35525 15602 35591 15605
rect 39520 15602 40000 15632
rect 35525 15600 40000 15602
rect 35525 15544 35530 15600
rect 35586 15544 40000 15600
rect 35525 15542 40000 15544
rect 35525 15539 35591 15542
rect 39520 15512 40000 15542
rect 0 14650 480 14680
rect 1853 14650 1919 14653
rect 0 14648 1919 14650
rect 0 14592 1858 14648
rect 1914 14592 1919 14648
rect 0 14590 1919 14592
rect 0 14560 480 14590
rect 1853 14587 1919 14590
rect 35801 14650 35867 14653
rect 39520 14650 40000 14680
rect 35801 14648 40000 14650
rect 35801 14592 35806 14648
rect 35862 14592 40000 14648
rect 35801 14590 40000 14592
rect 35801 14587 35867 14590
rect 39520 14560 40000 14590
rect 0 13834 480 13864
rect 1945 13834 2011 13837
rect 0 13832 2011 13834
rect 0 13776 1950 13832
rect 2006 13776 2011 13832
rect 0 13774 2011 13776
rect 0 13744 480 13774
rect 1945 13771 2011 13774
rect 35249 13834 35315 13837
rect 39520 13834 40000 13864
rect 35249 13832 40000 13834
rect 35249 13776 35254 13832
rect 35310 13776 40000 13832
rect 35249 13774 40000 13776
rect 35249 13771 35315 13774
rect 39520 13744 40000 13774
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 0 12882 480 12912
rect 1485 12882 1551 12885
rect 0 12880 1551 12882
rect 0 12824 1490 12880
rect 1546 12824 1551 12880
rect 0 12822 1551 12824
rect 0 12792 480 12822
rect 1485 12819 1551 12822
rect 35065 12882 35131 12885
rect 39520 12882 40000 12912
rect 35065 12880 40000 12882
rect 35065 12824 35070 12880
rect 35126 12824 40000 12880
rect 35065 12822 40000 12824
rect 35065 12819 35131 12822
rect 39520 12792 40000 12822
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 0 12066 480 12096
rect 1577 12066 1643 12069
rect 0 12064 1643 12066
rect 0 12008 1582 12064
rect 1638 12008 1643 12064
rect 0 12006 1643 12008
rect 0 11976 480 12006
rect 1577 12003 1643 12006
rect 35617 12066 35683 12069
rect 39520 12066 40000 12096
rect 35617 12064 40000 12066
rect 35617 12008 35622 12064
rect 35678 12008 40000 12064
rect 35617 12006 40000 12008
rect 35617 12003 35683 12006
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 39520 11976 40000 12006
rect 34277 11935 34597 11936
rect 16665 11658 16731 11661
rect 33317 11658 33383 11661
rect 16665 11656 33383 11658
rect 16665 11600 16670 11656
rect 16726 11600 33322 11656
rect 33378 11600 33383 11656
rect 16665 11598 33383 11600
rect 16665 11595 16731 11598
rect 33317 11595 33383 11598
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 0 11114 480 11144
rect 1577 11114 1643 11117
rect 0 11112 1643 11114
rect 0 11056 1582 11112
rect 1638 11056 1643 11112
rect 0 11054 1643 11056
rect 0 11024 480 11054
rect 1577 11051 1643 11054
rect 35617 11114 35683 11117
rect 39520 11114 40000 11144
rect 35617 11112 40000 11114
rect 35617 11056 35622 11112
rect 35678 11056 40000 11112
rect 35617 11054 40000 11056
rect 35617 11051 35683 11054
rect 39520 11024 40000 11054
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 19977 10706 20043 10709
rect 23381 10706 23447 10709
rect 19977 10704 23447 10706
rect 19977 10648 19982 10704
rect 20038 10648 23386 10704
rect 23442 10648 23447 10704
rect 19977 10646 23447 10648
rect 19977 10643 20043 10646
rect 23381 10643 23447 10646
rect 29729 10434 29795 10437
rect 35433 10434 35499 10437
rect 29729 10432 35499 10434
rect 29729 10376 29734 10432
rect 29790 10376 35438 10432
rect 35494 10376 35499 10432
rect 29729 10374 35499 10376
rect 29729 10371 29795 10374
rect 35433 10371 35499 10374
rect 14277 10368 14597 10369
rect 0 10298 480 10328
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 480 10238
rect 1485 10235 1551 10238
rect 35709 10298 35775 10301
rect 39520 10298 40000 10328
rect 35709 10296 40000 10298
rect 35709 10240 35714 10296
rect 35770 10240 40000 10296
rect 35709 10238 40000 10240
rect 35709 10235 35775 10238
rect 39520 10208 40000 10238
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 3417 9618 3483 9621
rect 28809 9618 28875 9621
rect 3417 9616 28875 9618
rect 3417 9560 3422 9616
rect 3478 9560 28814 9616
rect 28870 9560 28875 9616
rect 3417 9558 28875 9560
rect 3417 9555 3483 9558
rect 28809 9555 28875 9558
rect 18873 9482 18939 9485
rect 35433 9482 35499 9485
rect 18873 9480 35499 9482
rect 18873 9424 18878 9480
rect 18934 9424 35438 9480
rect 35494 9424 35499 9480
rect 18873 9422 35499 9424
rect 18873 9419 18939 9422
rect 35433 9419 35499 9422
rect 0 9346 480 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 480 9286
rect 1577 9283 1643 9286
rect 35617 9346 35683 9349
rect 39520 9346 40000 9376
rect 35617 9344 40000 9346
rect 35617 9288 35622 9344
rect 35678 9288 40000 9344
rect 35617 9286 40000 9288
rect 35617 9283 35683 9286
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 39520 9256 40000 9286
rect 27610 9215 27930 9216
rect 2037 9074 2103 9077
rect 12985 9074 13051 9077
rect 2037 9072 13051 9074
rect 2037 9016 2042 9072
rect 2098 9016 12990 9072
rect 13046 9016 13051 9072
rect 2037 9014 13051 9016
rect 2037 9011 2103 9014
rect 12985 9011 13051 9014
rect 23289 9074 23355 9077
rect 35433 9074 35499 9077
rect 23289 9072 35499 9074
rect 23289 9016 23294 9072
rect 23350 9016 35438 9072
rect 35494 9016 35499 9072
rect 23289 9014 35499 9016
rect 23289 9011 23355 9014
rect 35433 9011 35499 9014
rect 1669 8938 1735 8941
rect 20069 8938 20135 8941
rect 1669 8936 20135 8938
rect 1669 8880 1674 8936
rect 1730 8880 20074 8936
rect 20130 8880 20135 8936
rect 1669 8878 20135 8880
rect 1669 8875 1735 8878
rect 20069 8875 20135 8878
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 0 8530 480 8560
rect 2497 8530 2563 8533
rect 0 8528 2563 8530
rect 0 8472 2502 8528
rect 2558 8472 2563 8528
rect 0 8470 2563 8472
rect 0 8440 480 8470
rect 2497 8467 2563 8470
rect 5073 8530 5139 8533
rect 24761 8530 24827 8533
rect 35433 8530 35499 8533
rect 5073 8528 24827 8530
rect 5073 8472 5078 8528
rect 5134 8472 24766 8528
rect 24822 8472 24827 8528
rect 5073 8470 24827 8472
rect 5073 8467 5139 8470
rect 24761 8467 24827 8470
rect 24902 8528 35499 8530
rect 24902 8472 35438 8528
rect 35494 8472 35499 8528
rect 24902 8470 35499 8472
rect 12985 8394 13051 8397
rect 24669 8394 24735 8397
rect 24902 8394 24962 8470
rect 35433 8467 35499 8470
rect 36721 8530 36787 8533
rect 39520 8530 40000 8560
rect 36721 8528 40000 8530
rect 36721 8472 36726 8528
rect 36782 8472 40000 8528
rect 36721 8470 40000 8472
rect 36721 8467 36787 8470
rect 39520 8440 40000 8470
rect 12985 8392 14842 8394
rect 12985 8336 12990 8392
rect 13046 8336 14842 8392
rect 12985 8334 14842 8336
rect 12985 8331 13051 8334
rect 3049 8258 3115 8261
rect 14782 8258 14842 8334
rect 24669 8392 24962 8394
rect 24669 8336 24674 8392
rect 24730 8336 24962 8392
rect 24669 8334 24962 8336
rect 27478 8334 28090 8394
rect 24669 8331 24735 8334
rect 19977 8258 20043 8261
rect 27478 8258 27538 8334
rect 3049 8256 14106 8258
rect 3049 8200 3054 8256
rect 3110 8200 14106 8256
rect 3049 8198 14106 8200
rect 14782 8256 20043 8258
rect 14782 8200 19982 8256
rect 20038 8200 20043 8256
rect 14782 8198 20043 8200
rect 3049 8195 3115 8198
rect 2681 8122 2747 8125
rect 5073 8122 5139 8125
rect 2681 8120 5139 8122
rect 2681 8064 2686 8120
rect 2742 8064 5078 8120
rect 5134 8064 5139 8120
rect 2681 8062 5139 8064
rect 2681 8059 2747 8062
rect 5073 8059 5139 8062
rect 5625 8122 5691 8125
rect 5625 8120 8402 8122
rect 5625 8064 5630 8120
rect 5686 8064 8402 8120
rect 5625 8062 8402 8064
rect 5625 8059 5691 8062
rect 2037 7850 2103 7853
rect 8342 7850 8402 8062
rect 14046 7986 14106 8198
rect 19977 8195 20043 8198
rect 20118 8198 27538 8258
rect 28030 8258 28090 8334
rect 36537 8258 36603 8261
rect 28030 8256 36603 8258
rect 28030 8200 36542 8256
rect 36598 8200 36603 8256
rect 28030 8198 36603 8200
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 20118 8122 20178 8198
rect 36537 8195 36603 8198
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 14782 8062 20178 8122
rect 14782 7986 14842 8062
rect 35433 7986 35499 7989
rect 14046 7926 14842 7986
rect 17174 7984 35499 7986
rect 17174 7928 35438 7984
rect 35494 7928 35499 7984
rect 17174 7926 35499 7928
rect 17174 7850 17234 7926
rect 35433 7923 35499 7926
rect 2037 7848 8218 7850
rect 2037 7792 2042 7848
rect 2098 7792 8218 7848
rect 2037 7790 8218 7792
rect 8342 7790 17234 7850
rect 19885 7850 19951 7853
rect 34973 7850 35039 7853
rect 19885 7848 35039 7850
rect 19885 7792 19890 7848
rect 19946 7792 34978 7848
rect 35034 7792 35039 7848
rect 19885 7790 35039 7792
rect 2037 7787 2103 7790
rect 3969 7714 4035 7717
rect 5625 7714 5691 7717
rect 1350 7712 5691 7714
rect 1350 7656 3974 7712
rect 4030 7656 5630 7712
rect 5686 7656 5691 7712
rect 1350 7654 5691 7656
rect 0 7578 480 7608
rect 1350 7578 1410 7654
rect 3969 7651 4035 7654
rect 5625 7651 5691 7654
rect 7610 7648 7930 7649
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 0 7518 1410 7578
rect 2589 7578 2655 7581
rect 4337 7578 4403 7581
rect 2589 7576 4403 7578
rect 2589 7520 2594 7576
rect 2650 7520 4342 7576
rect 4398 7520 4403 7576
rect 2589 7518 4403 7520
rect 8158 7578 8218 7790
rect 19885 7787 19951 7790
rect 34973 7787 35039 7790
rect 10685 7714 10751 7717
rect 17217 7714 17283 7717
rect 10685 7712 17283 7714
rect 10685 7656 10690 7712
rect 10746 7656 17222 7712
rect 17278 7656 17283 7712
rect 10685 7654 17283 7656
rect 10685 7651 10751 7654
rect 17217 7651 17283 7654
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 14181 7578 14247 7581
rect 8158 7576 14247 7578
rect 8158 7520 14186 7576
rect 14242 7520 14247 7576
rect 8158 7518 14247 7520
rect 0 7488 480 7518
rect 2589 7515 2655 7518
rect 4337 7515 4403 7518
rect 14181 7515 14247 7518
rect 14365 7578 14431 7581
rect 39520 7578 40000 7608
rect 14365 7576 17418 7578
rect 14365 7520 14370 7576
rect 14426 7520 17418 7576
rect 14365 7518 17418 7520
rect 14365 7515 14431 7518
rect 6821 7442 6887 7445
rect 6821 7440 17050 7442
rect 6821 7384 6826 7440
rect 6882 7384 17050 7440
rect 6821 7382 17050 7384
rect 6821 7379 6887 7382
rect 13721 7306 13787 7309
rect 15377 7306 15443 7309
rect 13721 7304 15443 7306
rect 13721 7248 13726 7304
rect 13782 7248 15382 7304
rect 15438 7248 15443 7304
rect 13721 7246 15443 7248
rect 13721 7243 13787 7246
rect 15377 7243 15443 7246
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 16990 7034 17050 7382
rect 17358 7306 17418 7518
rect 34838 7518 40000 7578
rect 24761 7442 24827 7445
rect 34838 7442 34898 7518
rect 39520 7488 40000 7518
rect 24761 7440 34898 7442
rect 24761 7384 24766 7440
rect 24822 7384 34898 7440
rect 24761 7382 34898 7384
rect 24761 7379 24827 7382
rect 24209 7306 24275 7309
rect 24669 7306 24735 7309
rect 17358 7304 24735 7306
rect 17358 7248 24214 7304
rect 24270 7248 24674 7304
rect 24730 7248 24735 7304
rect 17358 7246 24735 7248
rect 24209 7243 24275 7246
rect 24669 7243 24735 7246
rect 17217 7170 17283 7173
rect 23289 7170 23355 7173
rect 17217 7168 23355 7170
rect 17217 7112 17222 7168
rect 17278 7112 23294 7168
rect 23350 7112 23355 7168
rect 17217 7110 23355 7112
rect 17217 7107 17283 7110
rect 23289 7107 23355 7110
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 19057 7034 19123 7037
rect 16990 7032 19123 7034
rect 16990 6976 19062 7032
rect 19118 6976 19123 7032
rect 16990 6974 19123 6976
rect 19057 6971 19123 6974
rect 18229 6898 18295 6901
rect 18229 6896 35634 6898
rect 18229 6840 18234 6896
rect 18290 6840 35634 6896
rect 18229 6838 35634 6840
rect 18229 6835 18295 6838
rect 0 6626 480 6656
rect 6821 6626 6887 6629
rect 0 6624 6887 6626
rect 0 6568 6826 6624
rect 6882 6568 6887 6624
rect 0 6566 6887 6568
rect 0 6536 480 6566
rect 6821 6563 6887 6566
rect 11329 6626 11395 6629
rect 13997 6626 14063 6629
rect 11329 6624 14063 6626
rect 11329 6568 11334 6624
rect 11390 6568 14002 6624
rect 14058 6568 14063 6624
rect 11329 6566 14063 6568
rect 35574 6626 35634 6838
rect 39520 6626 40000 6656
rect 35574 6566 40000 6626
rect 11329 6563 11395 6566
rect 13997 6563 14063 6566
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 39520 6536 40000 6566
rect 34277 6495 34597 6496
rect 17493 6354 17559 6357
rect 35433 6354 35499 6357
rect 1166 6352 35499 6354
rect 1166 6296 17498 6352
rect 17554 6296 35438 6352
rect 35494 6296 35499 6352
rect 1166 6294 35499 6296
rect 0 5810 480 5840
rect 1166 5810 1226 6294
rect 17493 6291 17559 6294
rect 35433 6291 35499 6294
rect 5901 6218 5967 6221
rect 7189 6218 7255 6221
rect 5901 6216 7255 6218
rect 5901 6160 5906 6216
rect 5962 6160 7194 6216
rect 7250 6160 7255 6216
rect 5901 6158 7255 6160
rect 5901 6155 5967 6158
rect 7189 6155 7255 6158
rect 9857 6218 9923 6221
rect 16389 6218 16455 6221
rect 18413 6218 18479 6221
rect 9857 6216 14106 6218
rect 9857 6160 9862 6216
rect 9918 6160 14106 6216
rect 9857 6158 14106 6160
rect 9857 6155 9923 6158
rect 2037 5946 2103 5949
rect 9857 5946 9923 5949
rect 2037 5944 9923 5946
rect 2037 5888 2042 5944
rect 2098 5888 9862 5944
rect 9918 5888 9923 5944
rect 2037 5886 9923 5888
rect 2037 5883 2103 5886
rect 9857 5883 9923 5886
rect 0 5750 1226 5810
rect 11145 5810 11211 5813
rect 14046 5810 14106 6158
rect 16389 6216 18479 6218
rect 16389 6160 16394 6216
rect 16450 6160 18418 6216
rect 18474 6160 18479 6216
rect 16389 6158 18479 6160
rect 16389 6155 16455 6158
rect 18413 6155 18479 6158
rect 19241 6218 19307 6221
rect 21081 6218 21147 6221
rect 19241 6216 21147 6218
rect 19241 6160 19246 6216
rect 19302 6160 21086 6216
rect 21142 6160 21147 6216
rect 19241 6158 21147 6160
rect 19241 6155 19307 6158
rect 21081 6155 21147 6158
rect 15193 6082 15259 6085
rect 25313 6082 25379 6085
rect 15193 6080 25379 6082
rect 15193 6024 15198 6080
rect 15254 6024 25318 6080
rect 25374 6024 25379 6080
rect 15193 6022 25379 6024
rect 15193 6019 15259 6022
rect 25313 6019 25379 6022
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 39520 5810 40000 5840
rect 11145 5808 13922 5810
rect 11145 5752 11150 5808
rect 11206 5752 13922 5808
rect 11145 5750 13922 5752
rect 14046 5750 40000 5810
rect 0 5720 480 5750
rect 11145 5747 11211 5750
rect 13862 5674 13922 5750
rect 39520 5720 40000 5750
rect 15745 5674 15811 5677
rect 13862 5672 15811 5674
rect 13862 5616 15750 5672
rect 15806 5616 15811 5672
rect 13862 5614 15811 5616
rect 15745 5611 15811 5614
rect 26877 5538 26943 5541
rect 33777 5538 33843 5541
rect 26877 5536 33843 5538
rect 26877 5480 26882 5536
rect 26938 5480 33782 5536
rect 33838 5480 33843 5536
rect 26877 5478 33843 5480
rect 26877 5475 26943 5478
rect 33777 5475 33843 5478
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 2037 5266 2103 5269
rect 26325 5266 26391 5269
rect 2037 5264 26391 5266
rect 2037 5208 2042 5264
rect 2098 5208 26330 5264
rect 26386 5208 26391 5264
rect 2037 5206 26391 5208
rect 2037 5203 2103 5206
rect 26325 5203 26391 5206
rect 28901 5266 28967 5269
rect 30649 5266 30715 5269
rect 28901 5264 30715 5266
rect 28901 5208 28906 5264
rect 28962 5208 30654 5264
rect 30710 5208 30715 5264
rect 28901 5206 30715 5208
rect 28901 5203 28967 5206
rect 30649 5203 30715 5206
rect 15101 5130 15167 5133
rect 17769 5130 17835 5133
rect 15101 5128 17835 5130
rect 15101 5072 15106 5128
rect 15162 5072 17774 5128
rect 17830 5072 17835 5128
rect 15101 5070 17835 5072
rect 15101 5067 15167 5070
rect 17769 5067 17835 5070
rect 10593 4994 10659 4997
rect 12525 4994 12591 4997
rect 10593 4992 12591 4994
rect 10593 4936 10598 4992
rect 10654 4936 12530 4992
rect 12586 4936 12591 4992
rect 10593 4934 12591 4936
rect 10593 4931 10659 4934
rect 12525 4931 12591 4934
rect 17677 4994 17743 4997
rect 21357 4994 21423 4997
rect 17677 4992 21423 4994
rect 17677 4936 17682 4992
rect 17738 4936 21362 4992
rect 21418 4936 21423 4992
rect 17677 4934 21423 4936
rect 17677 4931 17743 4934
rect 21357 4931 21423 4934
rect 21633 4994 21699 4997
rect 22737 4994 22803 4997
rect 21633 4992 22803 4994
rect 21633 4936 21638 4992
rect 21694 4936 22742 4992
rect 22798 4936 22803 4992
rect 21633 4934 22803 4936
rect 21633 4931 21699 4934
rect 22737 4931 22803 4934
rect 14277 4928 14597 4929
rect 0 4858 480 4888
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 17033 4858 17099 4861
rect 21357 4858 21423 4861
rect 22461 4858 22527 4861
rect 0 4824 12312 4858
rect 12390 4824 14106 4858
rect 0 4798 14106 4824
rect 0 4768 480 4798
rect 12252 4764 12450 4798
rect 14046 4722 14106 4798
rect 17033 4856 22527 4858
rect 17033 4800 17038 4856
rect 17094 4800 21362 4856
rect 21418 4800 22466 4856
rect 22522 4800 22527 4856
rect 17033 4798 22527 4800
rect 17033 4795 17099 4798
rect 21357 4795 21423 4798
rect 22461 4795 22527 4798
rect 33777 4858 33843 4861
rect 39520 4858 40000 4888
rect 33777 4856 40000 4858
rect 33777 4800 33782 4856
rect 33838 4800 40000 4856
rect 33777 4798 40000 4800
rect 33777 4795 33843 4798
rect 39520 4768 40000 4798
rect 26601 4722 26667 4725
rect 28993 4722 29059 4725
rect 14046 4720 29059 4722
rect 14046 4664 26606 4720
rect 26662 4664 28998 4720
rect 29054 4664 29059 4720
rect 14046 4662 29059 4664
rect 26601 4659 26667 4662
rect 28993 4659 29059 4662
rect 3601 4586 3667 4589
rect 10133 4586 10199 4589
rect 3601 4584 10199 4586
rect 3601 4528 3606 4584
rect 3662 4528 10138 4584
rect 10194 4528 10199 4584
rect 3601 4526 10199 4528
rect 3601 4523 3667 4526
rect 10133 4523 10199 4526
rect 15561 4586 15627 4589
rect 21633 4586 21699 4589
rect 15561 4584 21699 4586
rect 15561 4528 15566 4584
rect 15622 4528 21638 4584
rect 21694 4528 21699 4584
rect 15561 4526 21699 4528
rect 15561 4523 15627 4526
rect 21633 4523 21699 4526
rect 12801 4450 12867 4453
rect 16021 4450 16087 4453
rect 12801 4448 16087 4450
rect 12801 4392 12806 4448
rect 12862 4392 16026 4448
rect 16082 4392 16087 4448
rect 12801 4390 16087 4392
rect 12801 4387 12867 4390
rect 16021 4387 16087 4390
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 12525 4314 12591 4317
rect 15469 4314 15535 4317
rect 12525 4312 15535 4314
rect 12525 4256 12530 4312
rect 12586 4256 15474 4312
rect 15530 4256 15535 4312
rect 12525 4254 15535 4256
rect 12525 4251 12591 4254
rect 15469 4251 15535 4254
rect 3969 4178 4035 4181
rect 16389 4178 16455 4181
rect 3969 4176 16455 4178
rect 3969 4120 3974 4176
rect 4030 4120 16394 4176
rect 16450 4120 16455 4176
rect 3969 4118 16455 4120
rect 3969 4115 4035 4118
rect 16389 4115 16455 4118
rect 31293 4178 31359 4181
rect 31293 4176 35634 4178
rect 31293 4120 31298 4176
rect 31354 4120 35634 4176
rect 31293 4118 35634 4120
rect 31293 4115 31359 4118
rect 0 4042 480 4072
rect 2773 4042 2839 4045
rect 0 4040 2839 4042
rect 0 3984 2778 4040
rect 2834 3984 2839 4040
rect 0 3982 2839 3984
rect 0 3952 480 3982
rect 2773 3979 2839 3982
rect 22645 4042 22711 4045
rect 26509 4042 26575 4045
rect 22645 4040 26575 4042
rect 22645 3984 22650 4040
rect 22706 3984 26514 4040
rect 26570 3984 26575 4040
rect 22645 3982 26575 3984
rect 35574 4042 35634 4118
rect 39520 4042 40000 4072
rect 35574 3982 40000 4042
rect 22645 3979 22711 3982
rect 26509 3979 26575 3982
rect 39520 3952 40000 3982
rect 3417 3906 3483 3909
rect 5257 3906 5323 3909
rect 6453 3906 6519 3909
rect 9121 3906 9187 3909
rect 3417 3904 9187 3906
rect 3417 3848 3422 3904
rect 3478 3848 5262 3904
rect 5318 3848 6458 3904
rect 6514 3848 9126 3904
rect 9182 3848 9187 3904
rect 3417 3846 9187 3848
rect 3417 3843 3483 3846
rect 5257 3843 5323 3846
rect 6453 3843 6519 3846
rect 9121 3843 9187 3846
rect 20805 3906 20871 3909
rect 23473 3906 23539 3909
rect 20805 3904 23539 3906
rect 20805 3848 20810 3904
rect 20866 3848 23478 3904
rect 23534 3848 23539 3904
rect 20805 3846 23539 3848
rect 20805 3843 20871 3846
rect 23473 3843 23539 3846
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 2773 3772 2839 3773
rect 2773 3770 2820 3772
rect 2728 3768 2820 3770
rect 2728 3712 2778 3768
rect 2728 3710 2820 3712
rect 2773 3708 2820 3710
rect 2884 3708 2890 3772
rect 10225 3770 10291 3773
rect 12525 3770 12591 3773
rect 10225 3768 12591 3770
rect 10225 3712 10230 3768
rect 10286 3712 12530 3768
rect 12586 3712 12591 3768
rect 10225 3710 12591 3712
rect 2773 3707 2839 3708
rect 10225 3707 10291 3710
rect 12525 3707 12591 3710
rect 28942 3708 28948 3772
rect 29012 3770 29018 3772
rect 29085 3770 29151 3773
rect 29012 3768 29151 3770
rect 29012 3712 29090 3768
rect 29146 3712 29151 3768
rect 29012 3710 29151 3712
rect 29012 3708 29018 3710
rect 29085 3707 29151 3710
rect 9121 3634 9187 3637
rect 12249 3634 12315 3637
rect 13169 3634 13235 3637
rect 9121 3632 13235 3634
rect 9121 3576 9126 3632
rect 9182 3576 12254 3632
rect 12310 3576 13174 3632
rect 13230 3576 13235 3632
rect 9121 3574 13235 3576
rect 9121 3571 9187 3574
rect 12249 3571 12315 3574
rect 13169 3571 13235 3574
rect 14273 3634 14339 3637
rect 19885 3634 19951 3637
rect 14273 3632 19951 3634
rect 14273 3576 14278 3632
rect 14334 3576 19890 3632
rect 19946 3576 19951 3632
rect 14273 3574 19951 3576
rect 14273 3571 14339 3574
rect 19885 3571 19951 3574
rect 20253 3634 20319 3637
rect 30833 3634 30899 3637
rect 20253 3632 30899 3634
rect 20253 3576 20258 3632
rect 20314 3576 30838 3632
rect 30894 3576 30899 3632
rect 20253 3574 30899 3576
rect 20253 3571 20319 3574
rect 30833 3571 30899 3574
rect 2957 3498 3023 3501
rect 8753 3498 8819 3501
rect 2957 3496 8819 3498
rect 2957 3440 2962 3496
rect 3018 3440 8758 3496
rect 8814 3440 8819 3496
rect 2957 3438 8819 3440
rect 2957 3435 3023 3438
rect 8753 3435 8819 3438
rect 11053 3498 11119 3501
rect 15377 3498 15443 3501
rect 11053 3496 15443 3498
rect 11053 3440 11058 3496
rect 11114 3440 15382 3496
rect 15438 3440 15443 3496
rect 11053 3438 15443 3440
rect 11053 3435 11119 3438
rect 15377 3435 15443 3438
rect 8845 3362 8911 3365
rect 14181 3362 14247 3365
rect 16665 3362 16731 3365
rect 18321 3362 18387 3365
rect 19333 3362 19399 3365
rect 20805 3362 20871 3365
rect 8845 3360 20871 3362
rect 8845 3304 8850 3360
rect 8906 3304 14186 3360
rect 14242 3304 16670 3360
rect 16726 3304 18326 3360
rect 18382 3304 19338 3360
rect 19394 3304 20810 3360
rect 20866 3304 20871 3360
rect 8845 3302 20871 3304
rect 8845 3299 8911 3302
rect 14181 3299 14247 3302
rect 16665 3299 16731 3302
rect 18321 3299 18387 3302
rect 19333 3299 19399 3302
rect 20805 3299 20871 3302
rect 27429 3362 27495 3365
rect 27981 3362 28047 3365
rect 29085 3362 29151 3365
rect 27429 3360 29151 3362
rect 27429 3304 27434 3360
rect 27490 3304 27986 3360
rect 28042 3304 29090 3360
rect 29146 3304 29151 3360
rect 27429 3302 29151 3304
rect 27429 3299 27495 3302
rect 27981 3299 28047 3302
rect 29085 3299 29151 3302
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 9305 3226 9371 3229
rect 11881 3226 11947 3229
rect 17125 3226 17191 3229
rect 9305 3224 17191 3226
rect 9305 3168 9310 3224
rect 9366 3168 11886 3224
rect 11942 3168 17130 3224
rect 17186 3168 17191 3224
rect 9305 3166 17191 3168
rect 9305 3163 9371 3166
rect 11881 3163 11947 3166
rect 17125 3163 17191 3166
rect 0 3090 480 3120
rect 3969 3090 4035 3093
rect 0 3088 4035 3090
rect 0 3032 3974 3088
rect 4030 3032 4035 3088
rect 0 3030 4035 3032
rect 0 3000 480 3030
rect 3969 3027 4035 3030
rect 11513 3090 11579 3093
rect 22185 3090 22251 3093
rect 11513 3088 22251 3090
rect 11513 3032 11518 3088
rect 11574 3032 22190 3088
rect 22246 3032 22251 3088
rect 11513 3030 22251 3032
rect 11513 3027 11579 3030
rect 22185 3027 22251 3030
rect 22829 3090 22895 3093
rect 39520 3090 40000 3120
rect 22829 3088 40000 3090
rect 22829 3032 22834 3088
rect 22890 3032 40000 3088
rect 22829 3030 40000 3032
rect 22829 3027 22895 3030
rect 39520 3000 40000 3030
rect 7005 2954 7071 2957
rect 13813 2954 13879 2957
rect 7005 2952 13879 2954
rect 7005 2896 7010 2952
rect 7066 2896 13818 2952
rect 13874 2896 13879 2952
rect 7005 2894 13879 2896
rect 7005 2891 7071 2894
rect 13813 2891 13879 2894
rect 5533 2818 5599 2821
rect 8661 2818 8727 2821
rect 12249 2818 12315 2821
rect 5533 2816 12315 2818
rect 5533 2760 5538 2816
rect 5594 2760 8666 2816
rect 8722 2760 12254 2816
rect 12310 2760 12315 2816
rect 5533 2758 12315 2760
rect 5533 2755 5599 2758
rect 8661 2755 8727 2758
rect 12249 2755 12315 2758
rect 31661 2818 31727 2821
rect 34145 2818 34211 2821
rect 31661 2816 34211 2818
rect 31661 2760 31666 2816
rect 31722 2760 34150 2816
rect 34206 2760 34211 2816
rect 31661 2758 34211 2760
rect 31661 2755 31727 2758
rect 34145 2755 34211 2758
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 10685 2682 10751 2685
rect 1350 2680 10751 2682
rect 1350 2624 10690 2680
rect 10746 2624 10751 2680
rect 1350 2622 10751 2624
rect 0 2274 480 2304
rect 1350 2274 1410 2622
rect 10685 2619 10751 2622
rect 23105 2682 23171 2685
rect 26233 2682 26299 2685
rect 23105 2680 26299 2682
rect 23105 2624 23110 2680
rect 23166 2624 26238 2680
rect 26294 2624 26299 2680
rect 23105 2622 26299 2624
rect 23105 2619 23171 2622
rect 26233 2619 26299 2622
rect 11421 2546 11487 2549
rect 13721 2546 13787 2549
rect 13997 2546 14063 2549
rect 11421 2544 14063 2546
rect 11421 2488 11426 2544
rect 11482 2488 13726 2544
rect 13782 2488 14002 2544
rect 14058 2488 14063 2544
rect 11421 2486 14063 2488
rect 11421 2483 11487 2486
rect 13721 2483 13787 2486
rect 13997 2483 14063 2486
rect 17401 2546 17467 2549
rect 20069 2546 20135 2549
rect 17401 2544 20135 2546
rect 17401 2488 17406 2544
rect 17462 2488 20074 2544
rect 20130 2488 20135 2544
rect 17401 2486 20135 2488
rect 17401 2483 17467 2486
rect 20069 2483 20135 2486
rect 22461 2546 22527 2549
rect 25037 2546 25103 2549
rect 27613 2546 27679 2549
rect 22461 2544 27679 2546
rect 22461 2488 22466 2544
rect 22522 2488 25042 2544
rect 25098 2488 27618 2544
rect 27674 2488 27679 2544
rect 22461 2486 27679 2488
rect 22461 2483 22527 2486
rect 25037 2483 25103 2486
rect 27613 2483 27679 2486
rect 27797 2546 27863 2549
rect 32581 2546 32647 2549
rect 27797 2544 32647 2546
rect 27797 2488 27802 2544
rect 27858 2488 32586 2544
rect 32642 2488 32647 2544
rect 27797 2486 32647 2488
rect 27797 2483 27863 2486
rect 32581 2483 32647 2486
rect 1761 2410 1827 2413
rect 10501 2410 10567 2413
rect 1761 2408 10567 2410
rect 1761 2352 1766 2408
rect 1822 2352 10506 2408
rect 10562 2352 10567 2408
rect 1761 2350 10567 2352
rect 1761 2347 1827 2350
rect 10501 2347 10567 2350
rect 12065 2410 12131 2413
rect 13629 2410 13695 2413
rect 15653 2410 15719 2413
rect 12065 2408 13554 2410
rect 12065 2352 12070 2408
rect 12126 2352 13554 2408
rect 12065 2350 13554 2352
rect 12065 2347 12131 2350
rect 0 2214 1410 2274
rect 0 2184 480 2214
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 13494 2138 13554 2350
rect 13629 2408 15719 2410
rect 13629 2352 13634 2408
rect 13690 2352 15658 2408
rect 15714 2352 15719 2408
rect 13629 2350 15719 2352
rect 13629 2347 13695 2350
rect 15653 2347 15719 2350
rect 28901 2410 28967 2413
rect 38101 2410 38167 2413
rect 28901 2408 38167 2410
rect 28901 2352 28906 2408
rect 28962 2352 38106 2408
rect 38162 2352 38167 2408
rect 28901 2350 38167 2352
rect 28901 2347 28967 2350
rect 38101 2347 38167 2350
rect 39520 2274 40000 2304
rect 34838 2214 40000 2274
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 16757 2138 16823 2141
rect 19793 2138 19859 2141
rect 13494 2136 19859 2138
rect 13494 2080 16762 2136
rect 16818 2080 19798 2136
rect 19854 2080 19859 2136
rect 13494 2078 19859 2080
rect 16757 2075 16823 2078
rect 19793 2075 19859 2078
rect 28942 1940 28948 2004
rect 29012 2002 29018 2004
rect 34838 2002 34898 2214
rect 39520 2184 40000 2214
rect 29012 1942 34898 2002
rect 29012 1940 29018 1942
rect 23013 1594 23079 1597
rect 28942 1594 28948 1596
rect 23013 1592 28948 1594
rect 23013 1536 23018 1592
rect 23074 1536 28948 1592
rect 23013 1534 28948 1536
rect 23013 1531 23079 1534
rect 28942 1532 28948 1534
rect 29012 1532 29018 1596
rect 0 1322 480 1352
rect 13169 1322 13235 1325
rect 0 1320 13235 1322
rect 0 1264 13174 1320
rect 13230 1264 13235 1320
rect 0 1262 13235 1264
rect 0 1232 480 1262
rect 13169 1259 13235 1262
rect 25497 1322 25563 1325
rect 39520 1322 40000 1352
rect 25497 1320 40000 1322
rect 25497 1264 25502 1320
rect 25558 1264 40000 1320
rect 25497 1262 40000 1264
rect 25497 1259 25563 1262
rect 39520 1232 40000 1262
rect 0 506 480 536
rect 2865 506 2931 509
rect 0 504 2931 506
rect 0 448 2870 504
rect 2926 448 2931 504
rect 0 446 2931 448
rect 0 416 480 446
rect 2865 443 2931 446
rect 28942 444 28948 508
rect 29012 506 29018 508
rect 39520 506 40000 536
rect 29012 446 40000 506
rect 29012 444 29018 446
rect 39520 416 40000 446
rect 4245 234 4311 237
rect 4245 232 9690 234
rect 4245 176 4250 232
rect 4306 176 9690 232
rect 4245 174 9690 176
rect 4245 171 4311 174
rect 9630 98 9690 174
rect 19333 98 19399 101
rect 9630 96 19399 98
rect 9630 40 19338 96
rect 19394 40 19399 96
rect 9630 38 19399 40
rect 19333 35 19399 38
rect 28901 100 28967 101
rect 28901 96 28948 100
rect 29012 98 29018 100
rect 28901 40 28906 96
rect 28901 36 28948 40
rect 29012 38 29094 98
rect 29012 36 29018 38
rect 28901 35 28967 36
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 2820 3768 2884 3772
rect 2820 3712 2834 3768
rect 2834 3712 2884 3768
rect 2820 3708 2884 3712
rect 28948 3708 29012 3772
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
rect 28948 1940 29012 2004
rect 28948 1532 29012 1596
rect 28948 444 29012 508
rect 28948 96 29012 100
rect 28948 40 28962 96
rect 28962 40 29012 96
rect 28948 36 29012 40
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
rect 28947 2004 29013 2005
rect 28947 1940 28948 2004
rect 29012 1940 29013 2004
rect 28947 1939 29013 1940
rect 28950 1597 29010 1939
rect 28947 1596 29013 1597
rect 28947 1532 28948 1596
rect 29012 1532 29013 1596
rect 28947 1531 29013 1532
rect 28947 508 29013 509
rect 28947 444 28948 508
rect 29012 444 29013 508
rect 28947 443 29013 444
rect 28950 101 29010 443
rect 28947 100 29013 101
rect 28947 36 28948 100
rect 29012 36 29013 100
rect 28947 35 29013 36
<< via4 >>
rect 2734 3772 2970 3858
rect 2734 3708 2820 3772
rect 2820 3708 2884 3772
rect 2884 3708 2970 3772
rect 2734 3622 2970 3708
rect 28862 3772 29098 3858
rect 28862 3708 28948 3772
rect 28948 3708 29012 3772
rect 29012 3708 29098 3772
rect 28862 3622 29098 3708
<< metal5 >>
rect 2692 3858 29140 3900
rect 2692 3622 2734 3858
rect 2970 3622 28862 3858
rect 29098 3622 29140 3858
rect 2692 3580 29140 3622
use scs8hd_decap_3  FILLER_1_8 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_8 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__050__B tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_13 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_16 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__D
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__C
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _049_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_19
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__044__D
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__B
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _045_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_53 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_49
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_45
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__C
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_59
timestamp 1586364061
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_67
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _043_
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__D
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _037_
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__037__A
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_nor4_4  _056_
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 1602 592
use scs8hd_decap_8  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_104
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use scs8hd_or2_4  _076_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 682 592
use scs8hd_inv_8  _041_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__038__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__039__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _039_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _064_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__C
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_or4_4  _042_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__B
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__D
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _055_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_or4_4  _054_
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_167
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__D
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_176
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 866 592
use scs8hd_nor4_4  _068_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_201
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_198
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_205
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_202
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__C
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_209
timestamp 1586364061
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__D
timestamp 1586364061
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_213
timestamp 1586364061
transform 1 0 20700 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__D
timestamp 1586364061
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _083_
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 1602 592
use scs8hd_nor4_4  _084_
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__D
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__D
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__D
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__D
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_nor4_4  _085_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1602 592
use scs8hd_nor4_4  _082_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25392 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_266
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_262
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_270
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_270
timestamp 1586364061
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 25760 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_284
timestamp 1586364061
transform 1 0 27232 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_278
timestamp 1586364061
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_288
timestamp 1586364061
transform 1 0 27600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_292
timestamp 1586364061
transform 1 0 27968 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_291
timestamp 1586364061
transform 1 0 27876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27784 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 28060 0 -1 2720
box -38 -48 222 592
use scs8hd_conb_1  _097_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_296
timestamp 1586364061
transform 1 0 28336 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_295
timestamp 1586364061
transform 1 0 28244 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_300
timestamp 1586364061
transform 1 0 28704 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28520 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 28428 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28612 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_306
timestamp 1586364061
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_321
timestamp 1586364061
transform 1 0 30636 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_315
timestamp 1586364061
transform 1 0 30084 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_320
timestamp 1586364061
transform 1 0 30544 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _091_
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_0_329
timestamp 1586364061
transform 1 0 31372 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_325
timestamp 1586364061
transform 1 0 31004 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31188 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_336
timestamp 1586364061
transform 1 0 32016 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_332
timestamp 1586364061
transform 1 0 31648 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_337
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_333
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 32108 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31464 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30820 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33396 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_351
timestamp 1586364061
transform 1 0 33396 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_339
timestamp 1586364061
transform 1 0 32292 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_349
timestamp 1586364061
transform 1 0 33212 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_353
timestamp 1586364061
transform 1 0 33580 0 1 2720
box -38 -48 1142 592
use scs8hd_conb_1  _096_
timestamp 1586364061
transform 1 0 34132 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_362
timestamp 1586364061
transform 1 0 34408 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_370
timestamp 1586364061
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_365
timestamp 1586364061
transform 1 0 34684 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__050__D
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__C
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_8
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__052__C
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_22
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_26
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 590 592
use scs8hd_nor4_4  _044_
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_38
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_62
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_70
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__C
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_1  _060_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_100
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _038_
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__C
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _053_
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__D
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__D
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_133
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 314 592
use scs8hd_or4_4  _066_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__054__D
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _070_
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_195
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_conb_1  _095_
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__D
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__C
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__D
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _079_
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_2_249
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_253
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_257
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_271
timestamp 1586364061
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28244 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_287
timestamp 1586364061
transform 1 0 27508 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30268 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29900 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29256 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_304
timestamp 1586364061
transform 1 0 29072 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_308
timestamp 1586364061
transform 1 0 29440 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_315
timestamp 1586364061
transform 1 0 30084 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_328
timestamp 1586364061
transform 1 0 31280 0 -1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_346
timestamp 1586364061
transform 1 0 32936 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_350
timestamp 1586364061
transform 1 0 33304 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_362
timestamp 1586364061
transform 1 0 34408 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_374
timestamp 1586364061
transform 1 0 35512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_386
timestamp 1586364061
transform 1 0 36616 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_394
timestamp 1586364061
transform 1 0 37352 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_nor4_4  _052_
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 1602 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__D
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__B
timestamp 1586364061
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_48
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__D
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_60
timestamp 1586364061
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__046__C
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_67
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _057_
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__C
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__D
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_96
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_100
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_104
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _061_
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_nor4_4  _063_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _072_
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__C
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_150
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_154
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _073_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_224
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__D
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_256
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_260
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_267
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_271
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27692 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_287
timestamp 1586364061
transform 1 0 27508 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_291
timestamp 1586364061
transform 1 0 27876 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_295
timestamp 1586364061
transform 1 0 28244 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30268 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_309
timestamp 1586364061
transform 1 0 29532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_313
timestamp 1586364061
transform 1 0 29900 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31280 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_326
timestamp 1586364061
transform 1 0 31096 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _050_
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 1602 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__051__D
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_35
timestamp 1586364061
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _046_
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_39
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_69
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__057__D
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use scs8hd_nor4_4  _059_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _062_
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__058__D
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_115
timestamp 1586364061
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__D
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__C
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_160
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _071_
timestamp 1586364061
transform 1 0 16192 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__071__C
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _074_
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_181
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_185
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _078_
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 1602 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 21344 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_222
timestamp 1586364061
transform 1 0 21528 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_266
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 26956 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_279
timestamp 1586364061
transform 1 0 26772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_283
timestamp 1586364061
transform 1 0 27140 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27508 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_296
timestamp 1586364061
transform 1 0 28336 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 29072 0 -1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30636 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_313
timestamp 1586364061
transform 1 0 29900 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _051_
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1602 592
use scs8hd_buf_2  _101_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _092_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_65
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_69
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_103
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_107
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _048_
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use scs8hd_nor4_4  _058_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_140
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_144
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_or2_4  _081_
timestamp 1586364061
transform 1 0 16468 0 1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__D
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_163
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__C
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_218
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__C
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_235
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_239
timestamp 1586364061
transform 1 0 23092 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_248
timestamp 1586364061
transform 1 0 23920 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_252
timestamp 1586364061
transform 1 0 24288 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_265
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 27232 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_5_278
timestamp 1586364061
transform 1 0 26680 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_282
timestamp 1586364061
transform 1 0 27048 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27416 0 1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_5_295
timestamp 1586364061
transform 1 0 28244 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_303
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 35420 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_377
timestamp 1586364061
transform 1 0 35788 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_381
timestamp 1586364061
transform 1 0 36156 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_393
timestamp 1586364061
transform 1 0 37260 0 1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_5_405
timestamp 1586364061
transform 1 0 38364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_8
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__051__C
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_43
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_63
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_101
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__058__C
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__040__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  _040_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_130
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_126
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_164
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_171
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_189
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_193
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__D
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_212
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_226
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_230
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_229
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_243
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_conb_1  _093_
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_262
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_266
timestamp 1586364061
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_252
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_256
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _087_
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_285
timestamp 1586364061
transform 1 0 27324 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27508 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27876 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_289
timestamp 1586364061
transform 1 0 27692 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_293
timestamp 1586364061
transform 1 0 28060 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_305
timestamp 1586364061
transform 1 0 29164 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_317
timestamp 1586364061
transform 1 0 30268 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_329
timestamp 1586364061
transform 1 0 31372 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_335
timestamp 1586364061
transform 1 0 31924 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 35420 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_375
timestamp 1586364061
transform 1 0 35604 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_387
timestamp 1586364061
transform 1 0 36708 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_399
timestamp 1586364061
transform 1 0 37812 0 1 5984
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _094_
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_76
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_112
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_124
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_128
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _067_
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_240
timestamp 1586364061
transform 1 0 23184 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_244
timestamp 1586364061
transform 1 0 23552 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_8  _086_
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_261
timestamp 1586364061
transform 1 0 25116 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_265
timestamp 1586364061
transform 1 0 25484 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_377
timestamp 1586364061
transform 1 0 35788 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_389
timestamp 1586364061
transform 1 0 36892 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_30
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_47
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_55
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_106
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_165
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_192
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_198
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_202
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_209
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_213
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_342
timestamp 1586364061
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_354
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 35420 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 35236 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 36524 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_377
timestamp 1586364061
transform 1 0 35788 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_381
timestamp 1586364061
transform 1 0 36156 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_389
timestamp 1586364061
transform 1 0 36892 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_393
timestamp 1586364061
transform 1 0 37260 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_405
timestamp 1586364061
transform 1 0 38364 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_52
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_98
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_122
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_199
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_300
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_312
timestamp 1586364061
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_349
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_377
timestamp 1586364061
transform 1 0 35788 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_389
timestamp 1586364061
transform 1 0 36892 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_18
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_22
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_44
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_318
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_330
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_354
timestamp 1586364061
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 35420 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 35236 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 35972 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_377
timestamp 1586364061
transform 1 0 35788 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_381
timestamp 1586364061
transform 1 0 36156 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_393
timestamp 1586364061
transform 1 0 37260 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_11_405
timestamp 1586364061
transform 1 0 38364 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_349
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_361
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_377
timestamp 1586364061
transform 1 0 35788 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_389
timestamp 1586364061
transform 1 0 36892 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_293
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_300
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_312
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_324
timestamp 1586364061
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_342
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 35420 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_375
timestamp 1586364061
transform 1 0 35604 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_387
timestamp 1586364061
transform 1 0 36708 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_377
timestamp 1586364061
transform 1 0 35788 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_389
timestamp 1586364061
transform 1 0 36892 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_399
timestamp 1586364061
transform 1 0 37812 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_43
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_354
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 35420 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_375
timestamp 1586364061
transform 1 0 35604 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_387
timestamp 1586364061
transform 1 0 36708 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_399
timestamp 1586364061
transform 1 0 37812 0 1 10336
box -38 -48 774 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_288
timestamp 1586364061
transform 1 0 27600 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_300
timestamp 1586364061
transform 1 0 28704 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_312
timestamp 1586364061
transform 1 0 29808 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_324
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_361
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_293
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_379
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_391
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_403
timestamp 1586364061
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5354 0 5410 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 9034 0 9090 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 12622 0 12678 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 16302 0 16358 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 19890 0 19946 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 23570 0 23626 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 30838 0 30894 480 6 bottom_grid_pin_0_
port 6 nsew default tristate
rlabel metal2 s 34426 0 34482 480 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal2 s 38106 0 38162 480 6 bottom_grid_pin_8_
port 8 nsew default tristate
rlabel metal3 s 0 416 480 536 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 0 1232 480 1352 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal3 s 0 2184 480 2304 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 0 10208 480 10328 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 39520 416 40000 536 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 39520 2184 40000 2304 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 39520 3000 40000 3120 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 39520 3952 40000 4072 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 39520 4768 40000 4888 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 39520 5720 40000 5840 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal3 s 39520 6536 40000 6656 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 39520 7488 40000 7608 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 39520 8440 40000 8560 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 39520 9256 40000 9376 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 39520 10208 40000 10328 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 39520 11024 40000 11144 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 39520 11976 40000 12096 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 39520 12792 40000 12912 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 39520 13744 40000 13864 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 39520 15512 40000 15632 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 27158 0 27214 480 6 data_in
port 45 nsew default input
rlabel metal2 s 1766 0 1822 480 6 enable
port 46 nsew default input
rlabel metal2 s 33322 15520 33378 16000 6 top_grid_pin_14_
port 47 nsew default tristate
rlabel metal2 s 6642 15520 6698 16000 6 top_grid_pin_2_
port 48 nsew default tristate
rlabel metal2 s 19982 15520 20038 16000 6 top_grid_pin_6_
port 49 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 50 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 51 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 16000
<< end >>
