magic
tech sky130A
magscale 1 2
timestamp 1606223695
<< locali >>
rect 9505 12155 9539 12257
rect 7665 11067 7699 11237
rect 14105 10591 14139 10761
<< viali >>
rect 1685 12393 1719 12427
rect 4537 12393 4571 12427
rect 7941 12393 7975 12427
rect 2053 12257 2087 12291
rect 4445 12257 4479 12291
rect 6653 12257 6687 12291
rect 7849 12257 7883 12291
rect 8677 12257 8711 12291
rect 9505 12257 9539 12291
rect 15853 12257 15887 12291
rect 2145 12189 2179 12223
rect 2329 12189 2363 12223
rect 4629 12189 4663 12223
rect 6745 12189 6779 12223
rect 6929 12189 6963 12223
rect 8033 12189 8067 12223
rect 9505 12121 9539 12155
rect 4077 12053 4111 12087
rect 6285 12053 6319 12087
rect 7481 12053 7515 12087
rect 16037 12053 16071 12087
rect 1961 11849 1995 11883
rect 3985 11849 4019 11883
rect 8585 11849 8619 11883
rect 2513 11713 2547 11747
rect 4537 11713 4571 11747
rect 8033 11713 8067 11747
rect 9137 11713 9171 11747
rect 13001 11713 13035 11747
rect 15577 11713 15611 11747
rect 2329 11645 2363 11679
rect 3157 11645 3191 11679
rect 7757 11645 7791 11679
rect 8953 11645 8987 11679
rect 9045 11577 9079 11611
rect 15301 11577 15335 11611
rect 2421 11509 2455 11543
rect 3341 11509 3375 11543
rect 4353 11509 4387 11543
rect 4445 11509 4479 11543
rect 5181 11509 5215 11543
rect 7389 11509 7423 11543
rect 7849 11509 7883 11543
rect 12449 11509 12483 11543
rect 12817 11509 12851 11543
rect 12909 11509 12943 11543
rect 14933 11509 14967 11543
rect 15393 11509 15427 11543
rect 3341 11305 3375 11339
rect 4537 11305 4571 11339
rect 4905 11305 4939 11339
rect 9137 11305 9171 11339
rect 14289 11305 14323 11339
rect 15393 11305 15427 11339
rect 15761 11305 15795 11339
rect 4997 11237 5031 11271
rect 7665 11237 7699 11271
rect 8002 11237 8036 11271
rect 2228 11169 2262 11203
rect 5825 11169 5859 11203
rect 6092 11169 6126 11203
rect 1961 11101 1995 11135
rect 5181 11101 5215 11135
rect 7757 11169 7791 11203
rect 12909 11169 12943 11203
rect 13176 11169 13210 11203
rect 15853 11169 15887 11203
rect 15945 11101 15979 11135
rect 7205 11033 7239 11067
rect 7665 11033 7699 11067
rect 1685 10761 1719 10795
rect 4261 10761 4295 10795
rect 4721 10761 4755 10795
rect 12909 10761 12943 10795
rect 14105 10761 14139 10795
rect 15577 10761 15611 10795
rect 2329 10625 2363 10659
rect 5273 10625 5307 10659
rect 7849 10625 7883 10659
rect 13369 10625 13403 10659
rect 13553 10625 13587 10659
rect 2881 10557 2915 10591
rect 5089 10557 5123 10591
rect 7665 10557 7699 10591
rect 8677 10557 8711 10591
rect 8933 10557 8967 10591
rect 10517 10557 10551 10591
rect 14105 10557 14139 10591
rect 14197 10557 14231 10591
rect 3148 10489 3182 10523
rect 10784 10489 10818 10523
rect 14464 10489 14498 10523
rect 2053 10421 2087 10455
rect 2145 10421 2179 10455
rect 5181 10421 5215 10455
rect 7297 10421 7331 10455
rect 7757 10421 7791 10455
rect 10057 10421 10091 10455
rect 11897 10421 11931 10455
rect 13277 10421 13311 10455
rect 2329 10217 2363 10251
rect 2697 10217 2731 10251
rect 2789 10217 2823 10251
rect 12173 10217 12207 10251
rect 14381 10217 14415 10251
rect 15393 10217 15427 10251
rect 4874 10149 4908 10183
rect 10048 10149 10082 10183
rect 15853 10149 15887 10183
rect 1593 10081 1627 10115
rect 7573 10081 7607 10115
rect 8769 10081 8803 10115
rect 12265 10081 12299 10115
rect 14473 10081 14507 10115
rect 15761 10081 15795 10115
rect 2881 10013 2915 10047
rect 4629 10013 4663 10047
rect 7665 10013 7699 10047
rect 7849 10013 7883 10047
rect 8861 10013 8895 10047
rect 9045 10013 9079 10047
rect 9781 10013 9815 10047
rect 12357 10013 12391 10047
rect 13369 10013 13403 10047
rect 14657 10013 14691 10047
rect 15945 10013 15979 10047
rect 1777 9945 1811 9979
rect 6009 9945 6043 9979
rect 8401 9945 8435 9979
rect 7205 9877 7239 9911
rect 11161 9877 11195 9911
rect 11805 9877 11839 9911
rect 14013 9877 14047 9911
rect 2053 9673 2087 9707
rect 4721 9673 4755 9707
rect 5181 9673 5215 9707
rect 8217 9673 8251 9707
rect 5549 9605 5583 9639
rect 8677 9605 8711 9639
rect 15393 9605 15427 9639
rect 2697 9537 2731 9571
rect 6193 9537 6227 9571
rect 9229 9537 9263 9571
rect 10793 9537 10827 9571
rect 15945 9537 15979 9571
rect 3341 9469 3375 9503
rect 5365 9469 5399 9503
rect 6844 9469 6878 9503
rect 7104 9469 7138 9503
rect 11621 9469 11655 9503
rect 12449 9469 12483 9503
rect 14657 9469 14691 9503
rect 3586 9401 3620 9435
rect 6009 9401 6043 9435
rect 10701 9401 10735 9435
rect 12705 9401 12739 9435
rect 15853 9401 15887 9435
rect 2421 9333 2455 9367
rect 2513 9333 2547 9367
rect 5917 9333 5951 9367
rect 9045 9333 9079 9367
rect 9137 9333 9171 9367
rect 10241 9333 10275 9367
rect 10609 9333 10643 9367
rect 11437 9333 11471 9367
rect 13829 9333 13863 9367
rect 14841 9333 14875 9367
rect 15761 9333 15795 9367
rect 2053 9129 2087 9163
rect 6929 9129 6963 9163
rect 7297 9129 7331 9163
rect 8125 9129 8159 9163
rect 12541 9129 12575 9163
rect 13001 9129 13035 9163
rect 13369 9129 13403 9163
rect 15669 9129 15703 9163
rect 15761 9129 15795 9163
rect 10333 9061 10367 9095
rect 2421 8993 2455 9027
rect 3249 8993 3283 9027
rect 4077 8993 4111 9027
rect 5089 8993 5123 9027
rect 5345 8993 5379 9027
rect 8493 8993 8527 9027
rect 11161 8993 11195 9027
rect 11417 8993 11451 9027
rect 14473 8993 14507 9027
rect 1409 8925 1443 8959
rect 2513 8925 2547 8959
rect 2697 8925 2731 8959
rect 7389 8925 7423 8959
rect 7481 8925 7515 8959
rect 8585 8925 8619 8959
rect 8769 8925 8803 8959
rect 10425 8925 10459 8959
rect 10517 8925 10551 8959
rect 13461 8925 13495 8959
rect 13553 8925 13587 8959
rect 15853 8925 15887 8959
rect 6469 8857 6503 8891
rect 15301 8857 15335 8891
rect 3433 8789 3467 8823
rect 4261 8789 4295 8823
rect 9965 8789 9999 8823
rect 14657 8789 14691 8823
rect 3525 8585 3559 8619
rect 5365 8585 5399 8619
rect 6837 8585 6871 8619
rect 9873 8517 9907 8551
rect 11069 8517 11103 8551
rect 16037 8517 16071 8551
rect 3985 8449 4019 8483
rect 7389 8449 7423 8483
rect 10517 8449 10551 8483
rect 11621 8449 11655 8483
rect 13277 8449 13311 8483
rect 13461 8449 13495 8483
rect 14013 8449 14047 8483
rect 1409 8381 1443 8415
rect 2145 8381 2179 8415
rect 4252 8381 4286 8415
rect 5825 8381 5859 8415
rect 8033 8381 8067 8415
rect 10241 8381 10275 8415
rect 11437 8381 11471 8415
rect 15853 8381 15887 8415
rect 2412 8313 2446 8347
rect 7297 8313 7331 8347
rect 8300 8313 8334 8347
rect 11529 8313 11563 8347
rect 13185 8313 13219 8347
rect 14258 8313 14292 8347
rect 1593 8245 1627 8279
rect 6009 8245 6043 8279
rect 7205 8245 7239 8279
rect 9413 8245 9447 8279
rect 10333 8245 10367 8279
rect 12817 8245 12851 8279
rect 15393 8245 15427 8279
rect 1961 8041 1995 8075
rect 2789 8041 2823 8075
rect 3157 8041 3191 8075
rect 6745 8041 6779 8075
rect 8861 8041 8895 8075
rect 10149 8041 10183 8075
rect 10241 8041 10275 8075
rect 12541 8041 12575 8075
rect 13737 8041 13771 8075
rect 15669 8041 15703 8075
rect 15761 8041 15795 8075
rect 3249 7973 3283 8007
rect 11345 7973 11379 8007
rect 4905 7905 4939 7939
rect 5733 7905 5767 7939
rect 6653 7905 6687 7939
rect 7113 7905 7147 7939
rect 8769 7905 8803 7939
rect 11437 7905 11471 7939
rect 2053 7837 2087 7871
rect 2237 7837 2271 7871
rect 3341 7837 3375 7871
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 7205 7837 7239 7871
rect 7389 7837 7423 7871
rect 9045 7837 9079 7871
rect 10425 7837 10459 7871
rect 11529 7837 11563 7871
rect 12633 7837 12667 7871
rect 12817 7837 12851 7871
rect 13829 7837 13863 7871
rect 13921 7837 13955 7871
rect 14565 7837 14599 7871
rect 15853 7837 15887 7871
rect 5917 7769 5951 7803
rect 13369 7769 13403 7803
rect 1593 7701 1627 7735
rect 4537 7701 4571 7735
rect 6469 7701 6503 7735
rect 8401 7701 8435 7735
rect 9781 7701 9815 7735
rect 10977 7701 11011 7735
rect 12173 7701 12207 7735
rect 15301 7701 15335 7735
rect 2513 7497 2547 7531
rect 4905 7497 4939 7531
rect 9413 7497 9447 7531
rect 13829 7497 13863 7531
rect 11437 7429 11471 7463
rect 2973 7361 3007 7395
rect 3157 7361 3191 7395
rect 4169 7361 4203 7395
rect 4261 7361 4295 7395
rect 5457 7361 5491 7395
rect 6101 7361 6135 7395
rect 7389 7361 7423 7395
rect 11897 7361 11931 7395
rect 12081 7361 12115 7395
rect 14841 7361 14875 7395
rect 1581 7293 1615 7327
rect 2881 7293 2915 7327
rect 4077 7293 4111 7327
rect 7297 7293 7331 7327
rect 8125 7293 8159 7327
rect 9965 7293 9999 7327
rect 12449 7293 12483 7327
rect 12716 7293 12750 7327
rect 15853 7293 15887 7327
rect 5365 7225 5399 7259
rect 10210 7225 10244 7259
rect 11805 7225 11839 7259
rect 14749 7225 14783 7259
rect 1777 7157 1811 7191
rect 3709 7157 3743 7191
rect 5273 7157 5307 7191
rect 6837 7157 6871 7191
rect 7205 7157 7239 7191
rect 11345 7157 11379 7191
rect 14289 7157 14323 7191
rect 14657 7157 14691 7191
rect 16037 7157 16071 7191
rect 5089 6953 5123 6987
rect 7665 6953 7699 6987
rect 13185 6953 13219 6987
rect 15669 6953 15703 6987
rect 5457 6885 5491 6919
rect 13553 6885 13587 6919
rect 15761 6885 15795 6919
rect 1409 6817 1443 6851
rect 2412 6817 2446 6851
rect 4077 6817 4111 6851
rect 4997 6817 5031 6851
rect 6541 6817 6575 6851
rect 8493 6817 8527 6851
rect 8953 6817 8987 6851
rect 10149 6817 10183 6851
rect 11060 6817 11094 6851
rect 13645 6817 13679 6851
rect 14473 6817 14507 6851
rect 2145 6749 2179 6783
rect 5549 6749 5583 6783
rect 5641 6749 5675 6783
rect 6285 6749 6319 6783
rect 8585 6749 8619 6783
rect 8769 6749 8803 6783
rect 9229 6749 9263 6783
rect 10793 6749 10827 6783
rect 13829 6749 13863 6783
rect 15853 6749 15887 6783
rect 3525 6681 3559 6715
rect 8125 6681 8159 6715
rect 14657 6681 14691 6715
rect 1593 6613 1627 6647
rect 4261 6613 4295 6647
rect 4813 6613 4847 6647
rect 12173 6613 12207 6647
rect 15301 6613 15335 6647
rect 6837 6409 6871 6443
rect 11345 6409 11379 6443
rect 11805 6409 11839 6443
rect 16037 6409 16071 6443
rect 5825 6341 5859 6375
rect 8769 6341 8803 6375
rect 7389 6273 7423 6307
rect 9413 6273 9447 6307
rect 12909 6273 12943 6307
rect 13093 6273 13127 6307
rect 1685 6205 1719 6239
rect 2605 6205 2639 6239
rect 4445 6205 4479 6239
rect 9229 6205 9263 6239
rect 9965 6205 9999 6239
rect 11989 6205 12023 6239
rect 13645 6205 13679 6239
rect 13912 6205 13946 6239
rect 15853 6205 15887 6239
rect 1961 6137 1995 6171
rect 2850 6137 2884 6171
rect 4690 6137 4724 6171
rect 10232 6137 10266 6171
rect 3985 6069 4019 6103
rect 7205 6069 7239 6103
rect 7297 6069 7331 6103
rect 9137 6069 9171 6103
rect 12449 6069 12483 6103
rect 12817 6069 12851 6103
rect 15025 6069 15059 6103
rect 1961 5865 1995 5899
rect 2789 5865 2823 5899
rect 3157 5865 3191 5899
rect 3249 5865 3283 5899
rect 4445 5865 4479 5899
rect 4905 5865 4939 5899
rect 6745 5865 6779 5899
rect 8769 5865 8803 5899
rect 8861 5865 8895 5899
rect 14013 5865 14047 5899
rect 14381 5865 14415 5899
rect 6837 5797 6871 5831
rect 12072 5797 12106 5831
rect 14473 5797 14507 5831
rect 2053 5729 2087 5763
rect 4813 5729 4847 5763
rect 10517 5729 10551 5763
rect 15853 5729 15887 5763
rect 2237 5661 2271 5695
rect 3341 5661 3375 5695
rect 5089 5661 5123 5695
rect 7021 5661 7055 5695
rect 7573 5661 7607 5695
rect 9045 5661 9079 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 11805 5661 11839 5695
rect 14565 5661 14599 5695
rect 8401 5593 8435 5627
rect 1593 5525 1627 5559
rect 6377 5525 6411 5559
rect 10149 5525 10183 5559
rect 13185 5525 13219 5559
rect 16037 5525 16071 5559
rect 1961 5321 1995 5355
rect 3157 5321 3191 5355
rect 8217 5321 8251 5355
rect 10057 5253 10091 5287
rect 10517 5253 10551 5287
rect 11713 5253 11747 5287
rect 2421 5185 2455 5219
rect 2605 5185 2639 5219
rect 3709 5185 3743 5219
rect 4813 5185 4847 5219
rect 4997 5185 5031 5219
rect 6009 5185 6043 5219
rect 6193 5185 6227 5219
rect 11069 5185 11103 5219
rect 13093 5185 13127 5219
rect 14289 5185 14323 5219
rect 2329 5117 2363 5151
rect 4721 5117 4755 5151
rect 6837 5117 6871 5151
rect 8677 5117 8711 5151
rect 11897 5117 11931 5151
rect 13001 5117 13035 5151
rect 15853 5117 15887 5151
rect 7082 5049 7116 5083
rect 8944 5049 8978 5083
rect 14197 5049 14231 5083
rect 3525 4981 3559 5015
rect 3617 4981 3651 5015
rect 4353 4981 4387 5015
rect 5549 4981 5583 5015
rect 5917 4981 5951 5015
rect 10885 4981 10919 5015
rect 10977 4981 11011 5015
rect 12541 4981 12575 5015
rect 12909 4981 12943 5015
rect 13737 4981 13771 5015
rect 14105 4981 14139 5015
rect 16037 4981 16071 5015
rect 3525 4777 3559 4811
rect 5549 4777 5583 4811
rect 6377 4777 6411 4811
rect 6745 4777 6779 4811
rect 8125 4777 8159 4811
rect 9965 4777 9999 4811
rect 11621 4777 11655 4811
rect 12541 4777 12575 4811
rect 12909 4709 12943 4743
rect 13001 4709 13035 4743
rect 1409 4641 1443 4675
rect 2145 4641 2179 4675
rect 2412 4641 2446 4675
rect 4077 4641 4111 4675
rect 5641 4641 5675 4675
rect 10333 4641 10367 4675
rect 11529 4641 11563 4675
rect 15853 4641 15887 4675
rect 5825 4573 5859 4607
rect 6837 4573 6871 4607
rect 7021 4573 7055 4607
rect 8217 4573 8251 4607
rect 8309 4573 8343 4607
rect 10425 4573 10459 4607
rect 10609 4573 10643 4607
rect 11805 4573 11839 4607
rect 13093 4573 13127 4607
rect 1593 4437 1627 4471
rect 4261 4437 4295 4471
rect 5181 4437 5215 4471
rect 7757 4437 7791 4471
rect 11161 4437 11195 4471
rect 16037 4437 16071 4471
rect 2973 4233 3007 4267
rect 5549 4233 5583 4267
rect 7481 4233 7515 4267
rect 3433 4097 3467 4131
rect 3617 4097 3651 4131
rect 8125 4097 8159 4131
rect 10517 4097 10551 4131
rect 11713 4097 11747 4131
rect 13001 4097 13035 4131
rect 1593 4029 1627 4063
rect 3341 4029 3375 4063
rect 4169 4029 4203 4063
rect 7941 4029 7975 4063
rect 8677 4029 8711 4063
rect 8933 4029 8967 4063
rect 11529 4029 11563 4063
rect 14381 4029 14415 4063
rect 15117 4029 15151 4063
rect 15853 4029 15887 4063
rect 4436 3961 4470 3995
rect 12817 3961 12851 3995
rect 1777 3893 1811 3927
rect 7849 3893 7883 3927
rect 10057 3893 10091 3927
rect 11161 3893 11195 3927
rect 11621 3893 11655 3927
rect 12449 3893 12483 3927
rect 12909 3893 12943 3927
rect 14565 3893 14599 3927
rect 15301 3893 15335 3927
rect 16037 3893 16071 3927
rect 6837 3689 6871 3723
rect 8769 3689 8803 3723
rect 10149 3689 10183 3723
rect 10885 3689 10919 3723
rect 11345 3689 11379 3723
rect 5724 3621 5758 3655
rect 11253 3621 11287 3655
rect 1501 3553 1535 3587
rect 2421 3553 2455 3587
rect 3157 3553 3191 3587
rect 4077 3553 4111 3587
rect 5457 3553 5491 3587
rect 8677 3553 8711 3587
rect 10057 3553 10091 3587
rect 14473 3553 14507 3587
rect 15853 3553 15887 3587
rect 1685 3485 1719 3519
rect 8953 3485 8987 3519
rect 10241 3485 10275 3519
rect 11529 3485 11563 3519
rect 2605 3349 2639 3383
rect 3341 3349 3375 3383
rect 4261 3349 4295 3383
rect 8309 3349 8343 3383
rect 9689 3349 9723 3383
rect 14657 3349 14691 3383
rect 16037 3349 16071 3383
rect 1961 3145 1995 3179
rect 7021 3145 7055 3179
rect 9597 3145 9631 3179
rect 10977 3145 11011 3179
rect 7573 3009 7607 3043
rect 8217 3009 8251 3043
rect 11437 3009 11471 3043
rect 11529 3009 11563 3043
rect 1777 2941 1811 2975
rect 2513 2941 2547 2975
rect 3801 2941 3835 2975
rect 4721 2941 4755 2975
rect 5825 2941 5859 2975
rect 7389 2941 7423 2975
rect 10057 2941 10091 2975
rect 11345 2941 11379 2975
rect 12817 2941 12851 2975
rect 14197 2941 14231 2975
rect 14933 2941 14967 2975
rect 15853 2941 15887 2975
rect 4077 2873 4111 2907
rect 4997 2873 5031 2907
rect 6101 2873 6135 2907
rect 8484 2873 8518 2907
rect 10333 2873 10367 2907
rect 13093 2873 13127 2907
rect 2697 2805 2731 2839
rect 7481 2805 7515 2839
rect 14381 2805 14415 2839
rect 15117 2805 15151 2839
rect 16037 2805 16071 2839
rect 7665 2601 7699 2635
rect 8125 2601 8159 2635
rect 8033 2533 8067 2567
rect 1961 2465 1995 2499
rect 2697 2465 2731 2499
rect 11345 2465 11379 2499
rect 14657 2465 14691 2499
rect 15853 2465 15887 2499
rect 8217 2397 8251 2431
rect 11529 2397 11563 2431
rect 2145 2261 2179 2295
rect 2881 2261 2915 2295
rect 14841 2261 14875 2295
rect 16037 2261 16071 2295
<< metal1 >>
rect 3878 15240 3884 15292
rect 3936 15280 3942 15292
rect 6546 15280 6552 15292
rect 3936 15252 6552 15280
rect 3936 15240 3942 15252
rect 6546 15240 6552 15252
rect 6604 15240 6610 15292
rect 11882 15172 11888 15224
rect 11940 15212 11946 15224
rect 14918 15212 14924 15224
rect 11940 15184 14924 15212
rect 11940 15172 11946 15184
rect 14918 15172 14924 15184
rect 14976 15172 14982 15224
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 10318 14804 10324 14816
rect 3568 14776 10324 14804
rect 3568 14764 3574 14776
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 1104 14714 16836 14736
rect 1104 14662 6246 14714
rect 6298 14662 6310 14714
rect 6362 14662 6374 14714
rect 6426 14662 6438 14714
rect 6490 14662 11510 14714
rect 11562 14662 11574 14714
rect 11626 14662 11638 14714
rect 11690 14662 11702 14714
rect 11754 14662 16836 14714
rect 1104 14640 16836 14662
rect 1104 14170 16836 14192
rect 1104 14118 3614 14170
rect 3666 14118 3678 14170
rect 3730 14118 3742 14170
rect 3794 14118 3806 14170
rect 3858 14118 8878 14170
rect 8930 14118 8942 14170
rect 8994 14118 9006 14170
rect 9058 14118 9070 14170
rect 9122 14118 14142 14170
rect 14194 14118 14206 14170
rect 14258 14118 14270 14170
rect 14322 14118 14334 14170
rect 14386 14118 16836 14170
rect 1104 14096 16836 14118
rect 1104 13626 16836 13648
rect 1104 13574 6246 13626
rect 6298 13574 6310 13626
rect 6362 13574 6374 13626
rect 6426 13574 6438 13626
rect 6490 13574 11510 13626
rect 11562 13574 11574 13626
rect 11626 13574 11638 13626
rect 11690 13574 11702 13626
rect 11754 13574 16836 13626
rect 1104 13552 16836 13574
rect 1104 13082 16836 13104
rect 1104 13030 3614 13082
rect 3666 13030 3678 13082
rect 3730 13030 3742 13082
rect 3794 13030 3806 13082
rect 3858 13030 8878 13082
rect 8930 13030 8942 13082
rect 8994 13030 9006 13082
rect 9058 13030 9070 13082
rect 9122 13030 14142 13082
rect 14194 13030 14206 13082
rect 14258 13030 14270 13082
rect 14322 13030 14334 13082
rect 14386 13030 16836 13082
rect 1104 13008 16836 13030
rect 3510 12656 3516 12708
rect 3568 12696 3574 12708
rect 7650 12696 7656 12708
rect 3568 12668 7656 12696
rect 3568 12656 3574 12668
rect 7650 12656 7656 12668
rect 7708 12656 7714 12708
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 10778 12628 10784 12640
rect 4120 12600 10784 12628
rect 4120 12588 4126 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 1104 12538 16836 12560
rect 1104 12486 6246 12538
rect 6298 12486 6310 12538
rect 6362 12486 6374 12538
rect 6426 12486 6438 12538
rect 6490 12486 11510 12538
rect 11562 12486 11574 12538
rect 11626 12486 11638 12538
rect 11690 12486 11702 12538
rect 11754 12486 16836 12538
rect 1104 12464 16836 12486
rect 1673 12427 1731 12433
rect 1673 12393 1685 12427
rect 1719 12424 1731 12427
rect 4525 12427 4583 12433
rect 4525 12424 4537 12427
rect 1719 12396 4537 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 4525 12393 4537 12396
rect 4571 12393 4583 12427
rect 7926 12424 7932 12436
rect 7887 12396 7932 12424
rect 4525 12387 4583 12393
rect 7926 12384 7932 12396
rect 7984 12424 7990 12436
rect 13814 12424 13820 12436
rect 7984 12396 13820 12424
rect 7984 12384 7990 12396
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 9214 12356 9220 12368
rect 2924 12328 9220 12356
rect 2924 12316 2930 12328
rect 9214 12316 9220 12328
rect 9272 12316 9278 12368
rect 1946 12248 1952 12300
rect 2004 12288 2010 12300
rect 2041 12291 2099 12297
rect 2041 12288 2053 12291
rect 2004 12260 2053 12288
rect 2004 12248 2010 12260
rect 2041 12257 2053 12260
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 4028 12260 4445 12288
rect 4028 12248 4034 12260
rect 4433 12257 4445 12260
rect 4479 12257 4491 12291
rect 6638 12288 6644 12300
rect 6599 12260 6644 12288
rect 4433 12251 4491 12257
rect 6638 12248 6644 12260
rect 6696 12248 6702 12300
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 7650 12288 7656 12300
rect 7432 12260 7656 12288
rect 7432 12248 7438 12260
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 7883 12260 8677 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 8665 12257 8677 12260
rect 8711 12257 8723 12291
rect 8665 12251 8723 12257
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12288 9551 12291
rect 15841 12291 15899 12297
rect 15841 12288 15853 12291
rect 9539 12260 15853 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 15841 12257 15853 12260
rect 15887 12257 15899 12291
rect 15841 12251 15899 12257
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 3326 12220 3332 12232
rect 2363 12192 3332 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 4304 12192 4629 12220
rect 4304 12180 4310 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 5592 12192 6745 12220
rect 5592 12180 5598 12192
rect 6733 12189 6745 12192
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 6932 12152 6960 12183
rect 8018 12180 8024 12232
rect 8076 12220 8082 12232
rect 8076 12192 8121 12220
rect 8076 12180 8082 12192
rect 8202 12180 8208 12232
rect 8260 12220 8266 12232
rect 15654 12220 15660 12232
rect 8260 12192 15660 12220
rect 8260 12180 8266 12192
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 7834 12152 7840 12164
rect 6932 12124 7840 12152
rect 7834 12112 7840 12124
rect 7892 12112 7898 12164
rect 9493 12155 9551 12161
rect 9493 12152 9505 12155
rect 9232 12124 9505 12152
rect 3234 12044 3240 12096
rect 3292 12084 3298 12096
rect 4065 12087 4123 12093
rect 4065 12084 4077 12087
rect 3292 12056 4077 12084
rect 3292 12044 3298 12056
rect 4065 12053 4077 12056
rect 4111 12053 4123 12087
rect 4065 12047 4123 12053
rect 6086 12044 6092 12096
rect 6144 12084 6150 12096
rect 6273 12087 6331 12093
rect 6273 12084 6285 12087
rect 6144 12056 6285 12084
rect 6144 12044 6150 12056
rect 6273 12053 6285 12056
rect 6319 12053 6331 12087
rect 7466 12084 7472 12096
rect 7427 12056 7472 12084
rect 6273 12047 6331 12053
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 7650 12044 7656 12096
rect 7708 12084 7714 12096
rect 9232 12084 9260 12124
rect 9493 12121 9505 12124
rect 9539 12121 9551 12155
rect 9493 12115 9551 12121
rect 7708 12056 9260 12084
rect 7708 12044 7714 12056
rect 9306 12044 9312 12096
rect 9364 12084 9370 12096
rect 14826 12084 14832 12096
rect 9364 12056 14832 12084
rect 9364 12044 9370 12056
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 16025 12087 16083 12093
rect 16025 12053 16037 12087
rect 16071 12084 16083 12087
rect 16206 12084 16212 12096
rect 16071 12056 16212 12084
rect 16071 12053 16083 12056
rect 16025 12047 16083 12053
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 1104 11994 16836 12016
rect 1104 11942 3614 11994
rect 3666 11942 3678 11994
rect 3730 11942 3742 11994
rect 3794 11942 3806 11994
rect 3858 11942 8878 11994
rect 8930 11942 8942 11994
rect 8994 11942 9006 11994
rect 9058 11942 9070 11994
rect 9122 11942 14142 11994
rect 14194 11942 14206 11994
rect 14258 11942 14270 11994
rect 14322 11942 14334 11994
rect 14386 11942 16836 11994
rect 1104 11920 16836 11942
rect 1946 11880 1952 11892
rect 1907 11852 1952 11880
rect 1946 11840 1952 11852
rect 2004 11840 2010 11892
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3510 11880 3516 11892
rect 3016 11852 3516 11880
rect 3016 11840 3022 11852
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 3970 11880 3976 11892
rect 3931 11852 3976 11880
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 6638 11840 6644 11892
rect 6696 11880 6702 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 6696 11852 8585 11880
rect 6696 11840 6702 11852
rect 8573 11849 8585 11852
rect 8619 11849 8631 11883
rect 8573 11843 8631 11849
rect 3418 11772 3424 11824
rect 3476 11812 3482 11824
rect 5994 11812 6000 11824
rect 3476 11784 6000 11812
rect 3476 11772 3482 11784
rect 5994 11772 6000 11784
rect 6052 11772 6058 11824
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 9030 11812 9036 11824
rect 7892 11784 9036 11812
rect 7892 11772 7898 11784
rect 9030 11772 9036 11784
rect 9088 11772 9094 11824
rect 12158 11772 12164 11824
rect 12216 11812 12222 11824
rect 14550 11812 14556 11824
rect 12216 11784 14556 11812
rect 12216 11772 12222 11784
rect 14550 11772 14556 11784
rect 14608 11772 14614 11824
rect 2222 11704 2228 11756
rect 2280 11744 2286 11756
rect 2501 11747 2559 11753
rect 2501 11744 2513 11747
rect 2280 11716 2513 11744
rect 2280 11704 2286 11716
rect 2501 11713 2513 11716
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 4525 11747 4583 11753
rect 4525 11744 4537 11747
rect 3384 11716 4537 11744
rect 3384 11704 3390 11716
rect 4525 11713 4537 11716
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 7650 11704 7656 11756
rect 7708 11704 7714 11756
rect 8018 11744 8024 11756
rect 7979 11716 8024 11744
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9125 11747 9183 11753
rect 9125 11744 9137 11747
rect 8904 11716 9137 11744
rect 8904 11704 8910 11716
rect 9125 11713 9137 11716
rect 9171 11713 9183 11747
rect 9125 11707 9183 11713
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 11388 11716 13001 11744
rect 11388 11704 11394 11716
rect 12989 11713 13001 11716
rect 13035 11744 13047 11747
rect 13446 11744 13452 11756
rect 13035 11716 13452 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 13446 11704 13452 11716
rect 13504 11744 13510 11756
rect 14274 11744 14280 11756
rect 13504 11716 14280 11744
rect 13504 11704 13510 11716
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 15562 11744 15568 11756
rect 15523 11716 15568 11744
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 2314 11676 2320 11688
rect 2275 11648 2320 11676
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 3145 11679 3203 11685
rect 3145 11645 3157 11679
rect 3191 11676 3203 11679
rect 4982 11676 4988 11688
rect 3191 11648 4988 11676
rect 3191 11645 3203 11648
rect 3145 11639 3203 11645
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 5810 11636 5816 11688
rect 5868 11676 5874 11688
rect 7668 11676 7696 11704
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 5868 11648 7757 11676
rect 5868 11636 5874 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 7834 11636 7840 11688
rect 7892 11676 7898 11688
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 7892 11648 8953 11676
rect 7892 11636 7898 11648
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 15838 11676 15844 11688
rect 9456 11648 15844 11676
rect 9456 11636 9462 11648
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 9033 11611 9091 11617
rect 9033 11608 9045 11611
rect 7392 11580 9045 11608
rect 2406 11500 2412 11552
rect 2464 11540 2470 11552
rect 2464 11512 2509 11540
rect 2464 11500 2470 11512
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3329 11543 3387 11549
rect 3329 11540 3341 11543
rect 2832 11512 3341 11540
rect 2832 11500 2838 11512
rect 3329 11509 3341 11512
rect 3375 11509 3387 11543
rect 4338 11540 4344 11552
rect 4299 11512 4344 11540
rect 3329 11503 3387 11509
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 4430 11500 4436 11552
rect 4488 11540 4494 11552
rect 4488 11512 4533 11540
rect 4488 11500 4494 11512
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 7392 11549 7420 11580
rect 9033 11577 9045 11580
rect 9079 11577 9091 11611
rect 9033 11571 9091 11577
rect 15289 11611 15347 11617
rect 15289 11577 15301 11611
rect 15335 11608 15347 11611
rect 15654 11608 15660 11620
rect 15335 11580 15660 11608
rect 15335 11577 15347 11580
rect 15289 11571 15347 11577
rect 15654 11568 15660 11580
rect 15712 11568 15718 11620
rect 5169 11543 5227 11549
rect 5169 11540 5181 11543
rect 4948 11512 5181 11540
rect 4948 11500 4954 11512
rect 5169 11509 5181 11512
rect 5215 11509 5227 11543
rect 5169 11503 5227 11509
rect 7377 11543 7435 11549
rect 7377 11509 7389 11543
rect 7423 11509 7435 11543
rect 7377 11503 7435 11509
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 7837 11543 7895 11549
rect 7837 11540 7849 11543
rect 7616 11512 7849 11540
rect 7616 11500 7622 11512
rect 7837 11509 7849 11512
rect 7883 11540 7895 11543
rect 9306 11540 9312 11552
rect 7883 11512 9312 11540
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12802 11540 12808 11552
rect 12492 11512 12537 11540
rect 12763 11512 12808 11540
rect 12492 11500 12498 11512
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 14918 11540 14924 11552
rect 12952 11512 12997 11540
rect 14879 11512 14924 11540
rect 12952 11500 12958 11512
rect 14918 11500 14924 11512
rect 14976 11500 14982 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15436 11512 15481 11540
rect 15436 11500 15442 11512
rect 1104 11450 16836 11472
rect 1104 11398 6246 11450
rect 6298 11398 6310 11450
rect 6362 11398 6374 11450
rect 6426 11398 6438 11450
rect 6490 11398 11510 11450
rect 11562 11398 11574 11450
rect 11626 11398 11638 11450
rect 11690 11398 11702 11450
rect 11754 11398 16836 11450
rect 1104 11376 16836 11398
rect 3326 11336 3332 11348
rect 3287 11308 3332 11336
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4396 11308 4537 11336
rect 4396 11296 4402 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 4890 11336 4896 11348
rect 4851 11308 4896 11336
rect 4525 11299 4583 11305
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 8754 11296 8760 11348
rect 8812 11336 8818 11348
rect 9030 11336 9036 11348
rect 8812 11308 9036 11336
rect 8812 11296 8818 11308
rect 9030 11296 9036 11308
rect 9088 11336 9094 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 9088 11308 9137 11336
rect 9088 11296 9094 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 14274 11336 14280 11348
rect 14235 11308 14280 11336
rect 9125 11299 9183 11305
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 15378 11336 15384 11348
rect 15339 11308 15384 11336
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15746 11336 15752 11348
rect 15707 11308 15752 11336
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 4982 11268 4988 11280
rect 4943 11240 4988 11268
rect 4982 11228 4988 11240
rect 5040 11228 5046 11280
rect 6730 11268 6736 11280
rect 5828 11240 6736 11268
rect 2222 11209 2228 11212
rect 2216 11200 2228 11209
rect 2183 11172 2228 11200
rect 2216 11163 2228 11172
rect 2222 11160 2228 11163
rect 2280 11160 2286 11212
rect 5828 11209 5856 11240
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 7653 11271 7711 11277
rect 7653 11237 7665 11271
rect 7699 11268 7711 11271
rect 7990 11271 8048 11277
rect 7990 11268 8002 11271
rect 7699 11240 8002 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 7990 11237 8002 11240
rect 8036 11268 8048 11271
rect 8846 11268 8852 11280
rect 8036 11240 8852 11268
rect 8036 11237 8048 11240
rect 7990 11231 8048 11237
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 9214 11228 9220 11280
rect 9272 11268 9278 11280
rect 9272 11240 13676 11268
rect 9272 11228 9278 11240
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 6080 11203 6138 11209
rect 6080 11169 6092 11203
rect 6126 11200 6138 11203
rect 6638 11200 6644 11212
rect 6126 11172 6644 11200
rect 6126 11169 6138 11172
rect 6080 11163 6138 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 6748 11200 6776 11228
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 6748 11172 7757 11200
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 11882 11200 11888 11212
rect 8352 11172 11888 11200
rect 8352 11160 8358 11172
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 12897 11203 12955 11209
rect 12897 11169 12909 11203
rect 12943 11200 12955 11203
rect 12986 11200 12992 11212
rect 12943 11172 12992 11200
rect 12943 11169 12955 11172
rect 12897 11163 12955 11169
rect 12986 11160 12992 11172
rect 13044 11160 13050 11212
rect 13164 11203 13222 11209
rect 13164 11169 13176 11203
rect 13210 11200 13222 11203
rect 13538 11200 13544 11212
rect 13210 11172 13544 11200
rect 13210 11169 13222 11172
rect 13164 11163 13222 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 13648 11200 13676 11240
rect 13998 11228 14004 11280
rect 14056 11268 14062 11280
rect 15764 11268 15792 11296
rect 14056 11240 15792 11268
rect 14056 11228 14062 11240
rect 15841 11203 15899 11209
rect 15841 11200 15853 11203
rect 13648 11172 15853 11200
rect 15841 11169 15853 11172
rect 15887 11200 15899 11203
rect 16298 11200 16304 11212
rect 15887 11172 16304 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 16298 11160 16304 11172
rect 16356 11160 16362 11212
rect 1946 11132 1952 11144
rect 1907 11104 1952 11132
rect 1946 11092 1952 11104
rect 2004 11092 2010 11144
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5258 11132 5264 11144
rect 5215 11104 5264 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 15930 11092 15936 11144
rect 15988 11132 15994 11144
rect 15988 11104 16033 11132
rect 15988 11092 15994 11104
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 5810 11064 5816 11076
rect 4120 11036 5816 11064
rect 4120 11024 4126 11036
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 6822 11024 6828 11076
rect 6880 11064 6886 11076
rect 7193 11067 7251 11073
rect 7193 11064 7205 11067
rect 6880 11036 7205 11064
rect 6880 11024 6886 11036
rect 7193 11033 7205 11036
rect 7239 11064 7251 11067
rect 7653 11067 7711 11073
rect 7653 11064 7665 11067
rect 7239 11036 7665 11064
rect 7239 11033 7251 11036
rect 7193 11027 7251 11033
rect 7653 11033 7665 11036
rect 7699 11033 7711 11067
rect 7653 11027 7711 11033
rect 2590 10956 2596 11008
rect 2648 10996 2654 11008
rect 3142 10996 3148 11008
rect 2648 10968 3148 10996
rect 2648 10956 2654 10968
rect 3142 10956 3148 10968
rect 3200 10996 3206 11008
rect 13262 10996 13268 11008
rect 3200 10968 13268 10996
rect 3200 10956 3206 10968
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 1104 10906 16836 10928
rect 1104 10854 3614 10906
rect 3666 10854 3678 10906
rect 3730 10854 3742 10906
rect 3794 10854 3806 10906
rect 3858 10854 8878 10906
rect 8930 10854 8942 10906
rect 8994 10854 9006 10906
rect 9058 10854 9070 10906
rect 9122 10854 14142 10906
rect 14194 10854 14206 10906
rect 14258 10854 14270 10906
rect 14322 10854 14334 10906
rect 14386 10854 16836 10906
rect 1104 10832 16836 10854
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 2130 10792 2136 10804
rect 1719 10764 2136 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 4246 10792 4252 10804
rect 4207 10764 4252 10792
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4709 10795 4767 10801
rect 4709 10792 4721 10795
rect 4488 10764 4721 10792
rect 4488 10752 4494 10764
rect 4709 10761 4721 10764
rect 4755 10761 4767 10795
rect 4709 10755 4767 10761
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 11882 10792 11888 10804
rect 4856 10764 11888 10792
rect 4856 10752 4862 10764
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12894 10792 12900 10804
rect 12855 10764 12900 10792
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 12986 10752 12992 10804
rect 13044 10792 13050 10804
rect 14093 10795 14151 10801
rect 14093 10792 14105 10795
rect 13044 10764 14105 10792
rect 13044 10752 13050 10764
rect 14093 10761 14105 10764
rect 14139 10761 14151 10795
rect 15562 10792 15568 10804
rect 14093 10755 14151 10761
rect 14200 10764 15568 10792
rect 4062 10684 4068 10736
rect 4120 10724 4126 10736
rect 8202 10724 8208 10736
rect 4120 10696 8208 10724
rect 4120 10684 4126 10696
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 13998 10724 14004 10736
rect 11532 10696 14004 10724
rect 2222 10616 2228 10668
rect 2280 10656 2286 10668
rect 2317 10659 2375 10665
rect 2317 10656 2329 10659
rect 2280 10628 2329 10656
rect 2280 10616 2286 10628
rect 2317 10625 2329 10628
rect 2363 10656 2375 10659
rect 2363 10628 3004 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 1946 10548 1952 10600
rect 2004 10588 2010 10600
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2004 10560 2881 10588
rect 2004 10548 2010 10560
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 2976 10588 3004 10628
rect 4798 10616 4804 10668
rect 4856 10656 4862 10668
rect 4856 10628 5120 10656
rect 4856 10616 4862 10628
rect 5092 10597 5120 10628
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5316 10628 5409 10656
rect 5316 10616 5322 10628
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 7834 10656 7840 10668
rect 6696 10628 7840 10656
rect 6696 10616 6702 10628
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 9692 10628 10640 10656
rect 5077 10591 5135 10597
rect 2976 10560 4752 10588
rect 2869 10551 2927 10557
rect 2884 10520 2912 10551
rect 4724 10532 4752 10560
rect 5077 10557 5089 10591
rect 5123 10557 5135 10591
rect 5077 10551 5135 10557
rect 2958 10520 2964 10532
rect 2884 10492 2964 10520
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 3136 10523 3194 10529
rect 3136 10489 3148 10523
rect 3182 10520 3194 10523
rect 3326 10520 3332 10532
rect 3182 10492 3332 10520
rect 3182 10489 3194 10492
rect 3136 10483 3194 10489
rect 3326 10480 3332 10492
rect 3384 10480 3390 10532
rect 4706 10480 4712 10532
rect 4764 10520 4770 10532
rect 5276 10520 5304 10616
rect 5994 10548 6000 10600
rect 6052 10588 6058 10600
rect 7374 10588 7380 10600
rect 6052 10560 7380 10588
rect 6052 10548 6058 10560
rect 7374 10548 7380 10560
rect 7432 10588 7438 10600
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 7432 10560 7665 10588
rect 7432 10548 7438 10560
rect 7653 10557 7665 10560
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10557 8723 10591
rect 8665 10551 8723 10557
rect 4764 10492 5304 10520
rect 4764 10480 4770 10492
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 8680 10520 8708 10551
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 8921 10591 8979 10597
rect 8921 10588 8933 10591
rect 8812 10560 8933 10588
rect 8812 10548 8818 10560
rect 8921 10557 8933 10560
rect 8967 10557 8979 10591
rect 8921 10551 8979 10557
rect 9214 10548 9220 10600
rect 9272 10588 9278 10600
rect 9692 10588 9720 10628
rect 9272 10560 9720 10588
rect 9272 10548 9278 10560
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 10505 10591 10563 10597
rect 10505 10588 10517 10591
rect 9824 10560 10517 10588
rect 9824 10548 9830 10560
rect 10505 10557 10517 10560
rect 10551 10557 10563 10591
rect 10612 10588 10640 10628
rect 11532 10588 11560 10696
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 13354 10656 13360 10668
rect 13315 10628 13360 10656
rect 13354 10616 13360 10628
rect 13412 10616 13418 10668
rect 13538 10656 13544 10668
rect 13451 10628 13544 10656
rect 13538 10616 13544 10628
rect 13596 10656 13602 10668
rect 14200 10656 14228 10764
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 13596 10628 14228 10656
rect 13596 10616 13602 10628
rect 10612 10560 11560 10588
rect 10505 10551 10563 10557
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 14093 10591 14151 10597
rect 11940 10560 13124 10588
rect 11940 10548 11946 10560
rect 7064 10492 8616 10520
rect 8680 10492 8892 10520
rect 7064 10480 7070 10492
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 5169 10455 5227 10461
rect 2188 10424 2233 10452
rect 2188 10412 2194 10424
rect 5169 10421 5181 10455
rect 5215 10452 5227 10455
rect 5258 10452 5264 10464
rect 5215 10424 5264 10452
rect 5215 10421 5227 10424
rect 5169 10415 5227 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 7282 10452 7288 10464
rect 7243 10424 7288 10452
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7745 10455 7803 10461
rect 7745 10421 7757 10455
rect 7791 10452 7803 10455
rect 8110 10452 8116 10464
rect 7791 10424 8116 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 8588 10452 8616 10492
rect 8754 10452 8760 10464
rect 8588 10424 8760 10452
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 8864 10452 8892 10492
rect 9306 10480 9312 10532
rect 9364 10520 9370 10532
rect 10594 10520 10600 10532
rect 9364 10492 10600 10520
rect 9364 10480 9370 10492
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 10772 10523 10830 10529
rect 10772 10489 10784 10523
rect 10818 10520 10830 10523
rect 11330 10520 11336 10532
rect 10818 10492 11336 10520
rect 10818 10489 10830 10492
rect 10772 10483 10830 10489
rect 11330 10480 11336 10492
rect 11388 10480 11394 10532
rect 13096 10520 13124 10560
rect 14093 10557 14105 10591
rect 14139 10588 14151 10591
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 14139 10560 14197 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 13814 10520 13820 10532
rect 13096 10492 13820 10520
rect 13814 10480 13820 10492
rect 13872 10480 13878 10532
rect 14452 10523 14510 10529
rect 14452 10489 14464 10523
rect 14498 10520 14510 10523
rect 15194 10520 15200 10532
rect 14498 10492 15200 10520
rect 14498 10489 14510 10492
rect 14452 10483 14510 10489
rect 15194 10480 15200 10492
rect 15252 10480 15258 10532
rect 9766 10452 9772 10464
rect 8864 10424 9772 10452
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 11885 10455 11943 10461
rect 11885 10421 11897 10455
rect 11931 10452 11943 10455
rect 12710 10452 12716 10464
rect 11931 10424 12716 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 13262 10452 13268 10464
rect 13175 10424 13268 10452
rect 13262 10412 13268 10424
rect 13320 10452 13326 10464
rect 14550 10452 14556 10464
rect 13320 10424 14556 10452
rect 13320 10412 13326 10424
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 1104 10362 16836 10384
rect 1104 10310 6246 10362
rect 6298 10310 6310 10362
rect 6362 10310 6374 10362
rect 6426 10310 6438 10362
rect 6490 10310 11510 10362
rect 11562 10310 11574 10362
rect 11626 10310 11638 10362
rect 11690 10310 11702 10362
rect 11754 10310 16836 10362
rect 1104 10288 16836 10310
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2406 10248 2412 10260
rect 2363 10220 2412 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 2682 10248 2688 10260
rect 2643 10220 2688 10248
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 2866 10248 2872 10260
rect 2823 10220 2872 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 4614 10248 4620 10260
rect 3200 10220 4620 10248
rect 3200 10208 3206 10220
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5258 10248 5264 10260
rect 5132 10220 5264 10248
rect 5132 10208 5138 10220
rect 5258 10208 5264 10220
rect 5316 10248 5322 10260
rect 12161 10251 12219 10257
rect 5316 10220 10180 10248
rect 5316 10208 5322 10220
rect 1596 10152 4200 10180
rect 1596 10121 1624 10152
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 2958 10112 2964 10124
rect 2740 10084 2964 10112
rect 2740 10072 2746 10084
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 4172 10112 4200 10152
rect 4246 10140 4252 10192
rect 4304 10180 4310 10192
rect 4862 10183 4920 10189
rect 4862 10180 4874 10183
rect 4304 10152 4874 10180
rect 4304 10140 4310 10152
rect 4862 10149 4874 10152
rect 4908 10149 4920 10183
rect 4862 10143 4920 10149
rect 7374 10140 7380 10192
rect 7432 10180 7438 10192
rect 10042 10189 10048 10192
rect 10036 10180 10048 10189
rect 7432 10152 9904 10180
rect 10003 10152 10048 10180
rect 7432 10140 7438 10152
rect 7561 10115 7619 10121
rect 4172 10084 7512 10112
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10013 4675 10047
rect 4617 10007 4675 10013
rect 1765 9979 1823 9985
rect 1765 9945 1777 9979
rect 1811 9976 1823 9979
rect 1811 9948 2452 9976
rect 1811 9945 1823 9948
rect 1765 9939 1823 9945
rect 2424 9908 2452 9948
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 2884 9976 2912 10007
rect 2740 9948 2912 9976
rect 2740 9936 2746 9948
rect 4062 9908 4068 9920
rect 2424 9880 4068 9908
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4632 9908 4660 10007
rect 5997 9979 6055 9985
rect 5997 9945 6009 9979
rect 6043 9976 6055 9979
rect 7098 9976 7104 9988
rect 6043 9948 7104 9976
rect 6043 9945 6055 9948
rect 5997 9939 6055 9945
rect 7098 9936 7104 9948
rect 7156 9936 7162 9988
rect 4798 9908 4804 9920
rect 4632 9880 4804 9908
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7193 9911 7251 9917
rect 7193 9908 7205 9911
rect 6972 9880 7205 9908
rect 6972 9868 6978 9880
rect 7193 9877 7205 9880
rect 7239 9877 7251 9911
rect 7484 9908 7512 10084
rect 7561 10081 7573 10115
rect 7607 10112 7619 10115
rect 8662 10112 8668 10124
rect 7607 10084 8668 10112
rect 7607 10081 7619 10084
rect 7561 10075 7619 10081
rect 8662 10072 8668 10084
rect 8720 10072 8726 10124
rect 8754 10072 8760 10124
rect 8812 10112 8818 10124
rect 9876 10112 9904 10152
rect 10036 10143 10048 10152
rect 10042 10140 10048 10143
rect 10100 10140 10106 10192
rect 10152 10180 10180 10220
rect 12161 10217 12173 10251
rect 12207 10248 12219 10251
rect 12434 10248 12440 10260
rect 12207 10220 12440 10248
rect 12207 10217 12219 10220
rect 12161 10211 12219 10217
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 12618 10208 12624 10260
rect 12676 10248 12682 10260
rect 13078 10248 13084 10260
rect 12676 10220 13084 10248
rect 12676 10208 12682 10220
rect 13078 10208 13084 10220
rect 13136 10248 13142 10260
rect 13354 10248 13360 10260
rect 13136 10220 13360 10248
rect 13136 10208 13142 10220
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 14369 10251 14427 10257
rect 14369 10217 14381 10251
rect 14415 10248 14427 10251
rect 15381 10251 15439 10257
rect 15381 10248 15393 10251
rect 14415 10220 15393 10248
rect 14415 10217 14427 10220
rect 14369 10211 14427 10217
rect 15381 10217 15393 10220
rect 15427 10217 15439 10251
rect 15381 10211 15439 10217
rect 13722 10180 13728 10192
rect 10152 10152 13728 10180
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 15102 10180 15108 10192
rect 14384 10152 15108 10180
rect 12253 10115 12311 10121
rect 8812 10084 9444 10112
rect 9876 10084 12204 10112
rect 8812 10072 8818 10084
rect 7650 10044 7656 10056
rect 7611 10016 7656 10044
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7834 10044 7840 10056
rect 7795 10016 7840 10044
rect 7834 10004 7840 10016
rect 7892 10004 7898 10056
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 8168 10016 8432 10044
rect 8168 10004 8174 10016
rect 8404 9985 8432 10016
rect 8478 10004 8484 10056
rect 8536 10044 8542 10056
rect 8849 10047 8907 10053
rect 8849 10044 8861 10047
rect 8536 10016 8861 10044
rect 8536 10004 8542 10016
rect 8849 10013 8861 10016
rect 8895 10013 8907 10047
rect 8849 10007 8907 10013
rect 9033 10047 9091 10053
rect 9033 10013 9045 10047
rect 9079 10044 9091 10047
rect 9214 10044 9220 10056
rect 9079 10016 9220 10044
rect 9079 10013 9091 10016
rect 9033 10007 9091 10013
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 8389 9979 8447 9985
rect 8389 9945 8401 9979
rect 8435 9945 8447 9979
rect 8389 9939 8447 9945
rect 8754 9908 8760 9920
rect 7484 9880 8760 9908
rect 7193 9871 7251 9877
rect 8754 9868 8760 9880
rect 8812 9908 8818 9920
rect 9306 9908 9312 9920
rect 8812 9880 9312 9908
rect 8812 9868 8818 9880
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9416 9908 9444 10084
rect 9766 10044 9772 10056
rect 9727 10016 9772 10044
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 12176 9976 12204 10084
rect 12253 10081 12265 10115
rect 12299 10112 12311 10115
rect 13998 10112 14004 10124
rect 12299 10084 14004 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10044 12403 10047
rect 12710 10044 12716 10056
rect 12391 10016 12716 10044
rect 12391 10013 12403 10016
rect 12345 10007 12403 10013
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 13354 10044 13360 10056
rect 13315 10016 13360 10044
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 14384 10044 14412 10152
rect 15102 10140 15108 10152
rect 15160 10140 15166 10192
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 15841 10183 15899 10189
rect 15841 10180 15853 10183
rect 15344 10152 15853 10180
rect 15344 10140 15350 10152
rect 15841 10149 15853 10152
rect 15887 10149 15899 10183
rect 15841 10143 15899 10149
rect 14461 10115 14519 10121
rect 14461 10081 14473 10115
rect 14507 10112 14519 10115
rect 15378 10112 15384 10124
rect 14507 10084 15384 10112
rect 14507 10081 14519 10084
rect 14461 10075 14519 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15749 10115 15807 10121
rect 15749 10081 15761 10115
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 13556 10016 14412 10044
rect 14645 10047 14703 10053
rect 13556 9976 13584 10016
rect 14645 10013 14657 10047
rect 14691 10044 14703 10047
rect 15562 10044 15568 10056
rect 14691 10016 15568 10044
rect 14691 10013 14703 10016
rect 14645 10007 14703 10013
rect 15562 10004 15568 10016
rect 15620 10004 15626 10056
rect 11072 9948 12112 9976
rect 12176 9948 13584 9976
rect 11072 9908 11100 9948
rect 9416 9880 11100 9908
rect 11149 9911 11207 9917
rect 11149 9877 11161 9911
rect 11195 9908 11207 9911
rect 11238 9908 11244 9920
rect 11195 9880 11244 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 11793 9911 11851 9917
rect 11793 9877 11805 9911
rect 11839 9908 11851 9911
rect 11974 9908 11980 9920
rect 11839 9880 11980 9908
rect 11839 9877 11851 9880
rect 11793 9871 11851 9877
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 12084 9908 12112 9948
rect 13630 9936 13636 9988
rect 13688 9976 13694 9988
rect 15764 9976 15792 10075
rect 15930 10004 15936 10056
rect 15988 10044 15994 10056
rect 15988 10016 16033 10044
rect 15988 10004 15994 10016
rect 16022 9976 16028 9988
rect 13688 9948 16028 9976
rect 13688 9936 13694 9948
rect 16022 9936 16028 9948
rect 16080 9936 16086 9988
rect 13906 9908 13912 9920
rect 12084 9880 13912 9908
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14001 9911 14059 9917
rect 14001 9877 14013 9911
rect 14047 9908 14059 9911
rect 15746 9908 15752 9920
rect 14047 9880 15752 9908
rect 14047 9877 14059 9880
rect 14001 9871 14059 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 1104 9818 16836 9840
rect 1104 9766 3614 9818
rect 3666 9766 3678 9818
rect 3730 9766 3742 9818
rect 3794 9766 3806 9818
rect 3858 9766 8878 9818
rect 8930 9766 8942 9818
rect 8994 9766 9006 9818
rect 9058 9766 9070 9818
rect 9122 9766 14142 9818
rect 14194 9766 14206 9818
rect 14258 9766 14270 9818
rect 14322 9766 14334 9818
rect 14386 9766 16836 9818
rect 1104 9744 16836 9766
rect 2038 9704 2044 9716
rect 1999 9676 2044 9704
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 4062 9704 4068 9716
rect 3016 9676 4068 9704
rect 3016 9664 3022 9676
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 4706 9704 4712 9716
rect 4667 9676 4712 9704
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 5169 9707 5227 9713
rect 5169 9704 5181 9707
rect 4856 9676 5181 9704
rect 4856 9664 4862 9676
rect 5169 9673 5181 9676
rect 5215 9704 5227 9707
rect 6730 9704 6736 9716
rect 5215 9676 6736 9704
rect 5215 9673 5227 9676
rect 5169 9667 5227 9673
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7156 9676 7788 9704
rect 7156 9664 7162 9676
rect 2314 9596 2320 9648
rect 2372 9636 2378 9648
rect 5534 9636 5540 9648
rect 2372 9608 3372 9636
rect 5495 9608 5540 9636
rect 2372 9596 2378 9608
rect 2682 9568 2688 9580
rect 2595 9540 2688 9568
rect 2682 9528 2688 9540
rect 2740 9568 2746 9580
rect 3344 9568 3372 9608
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 6822 9636 6828 9648
rect 6196 9608 6828 9636
rect 6196 9577 6224 9608
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 7760 9636 7788 9676
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 7892 9676 8217 9704
rect 7892 9664 7898 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 8205 9667 8263 9673
rect 12452 9676 13400 9704
rect 8662 9636 8668 9648
rect 7760 9608 8524 9636
rect 8623 9608 8668 9636
rect 6181 9571 6239 9577
rect 2740 9540 3096 9568
rect 3344 9540 3464 9568
rect 2740 9528 2746 9540
rect 3068 9432 3096 9540
rect 3326 9500 3332 9512
rect 3287 9472 3332 9500
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 3436 9500 3464 9540
rect 5184 9540 6132 9568
rect 5184 9500 5212 9540
rect 5350 9500 5356 9512
rect 3436 9472 5212 9500
rect 5311 9472 5356 9500
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 6104 9500 6132 9540
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 8496 9568 8524 9608
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 10318 9596 10324 9648
rect 10376 9636 10382 9648
rect 12452 9636 12480 9676
rect 10376 9608 12480 9636
rect 13372 9636 13400 9676
rect 14642 9664 14648 9716
rect 14700 9704 14706 9716
rect 16390 9704 16396 9716
rect 14700 9676 16396 9704
rect 14700 9664 14706 9676
rect 16390 9664 16396 9676
rect 16448 9664 16454 9716
rect 15010 9636 15016 9648
rect 13372 9608 15016 9636
rect 10376 9596 10382 9608
rect 15010 9596 15016 9608
rect 15068 9596 15074 9648
rect 15378 9636 15384 9648
rect 15339 9608 15384 9636
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 9214 9568 9220 9580
rect 6181 9531 6239 9537
rect 6656 9540 6960 9568
rect 8496 9540 9220 9568
rect 6656 9500 6684 9540
rect 6104 9472 6684 9500
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 6832 9503 6890 9509
rect 6832 9500 6844 9503
rect 6788 9472 6844 9500
rect 6788 9460 6794 9472
rect 6832 9469 6844 9472
rect 6878 9469 6890 9503
rect 6932 9500 6960 9540
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 10502 9568 10508 9580
rect 10100 9540 10508 9568
rect 10100 9528 10106 9540
rect 10502 9528 10508 9540
rect 10560 9568 10566 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10560 9540 10793 9568
rect 10560 9528 10566 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10870 9528 10876 9580
rect 10928 9568 10934 9580
rect 14458 9568 14464 9580
rect 10928 9540 12572 9568
rect 10928 9528 10934 9540
rect 7098 9509 7104 9512
rect 6932 9472 7052 9500
rect 6832 9463 6890 9469
rect 3510 9432 3516 9444
rect 3068 9404 3516 9432
rect 3510 9392 3516 9404
rect 3568 9441 3574 9444
rect 3568 9435 3632 9441
rect 3568 9401 3586 9435
rect 3620 9401 3632 9435
rect 3568 9395 3632 9401
rect 3568 9392 3574 9395
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 5626 9432 5632 9444
rect 4212 9404 5632 9432
rect 4212 9392 4218 9404
rect 5626 9392 5632 9404
rect 5684 9392 5690 9444
rect 5997 9435 6055 9441
rect 5997 9401 6009 9435
rect 6043 9432 6055 9435
rect 6914 9432 6920 9444
rect 6043 9404 6920 9432
rect 6043 9401 6055 9404
rect 5997 9395 6055 9401
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 7024 9432 7052 9472
rect 7092 9463 7104 9509
rect 7156 9500 7162 9512
rect 7156 9472 7192 9500
rect 7098 9460 7104 9463
rect 7156 9460 7162 9472
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 11609 9503 11667 9509
rect 7432 9472 10732 9500
rect 7432 9460 7438 9472
rect 10704 9444 10732 9472
rect 11609 9469 11621 9503
rect 11655 9500 11667 9503
rect 11790 9500 11796 9512
rect 11655 9472 11796 9500
rect 11655 9469 11667 9472
rect 11609 9463 11667 9469
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12544 9500 12572 9540
rect 13464 9540 14464 9568
rect 13464 9500 13492 9540
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 14826 9528 14832 9580
rect 14884 9528 14890 9580
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 15930 9568 15936 9580
rect 15252 9540 15936 9568
rect 15252 9528 15258 9540
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 12544 9472 13492 9500
rect 12437 9463 12495 9469
rect 10686 9432 10692 9444
rect 7024 9404 10548 9432
rect 10647 9404 10692 9432
rect 2406 9364 2412 9376
rect 2367 9336 2412 9364
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 2501 9367 2559 9373
rect 2501 9333 2513 9367
rect 2547 9364 2559 9367
rect 2866 9364 2872 9376
rect 2547 9336 2872 9364
rect 2547 9333 2559 9336
rect 2501 9327 2559 9333
rect 2866 9324 2872 9336
rect 2924 9364 2930 9376
rect 5718 9364 5724 9376
rect 2924 9336 5724 9364
rect 2924 9324 2930 9336
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 5905 9367 5963 9373
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 7282 9364 7288 9376
rect 5951 9336 7288 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 10226 9364 10232 9376
rect 9180 9336 9225 9364
rect 10187 9336 10232 9364
rect 9180 9324 9186 9336
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 10520 9364 10548 9404
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 12452 9432 12480 9463
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14645 9503 14703 9509
rect 14645 9500 14657 9503
rect 13872 9472 14657 9500
rect 13872 9460 13878 9472
rect 14645 9469 14657 9472
rect 14691 9469 14703 9503
rect 14645 9463 14703 9469
rect 12701 9441 12707 9444
rect 11440 9404 12480 9432
rect 10594 9364 10600 9376
rect 10520 9336 10600 9364
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11440 9373 11468 9404
rect 11425 9367 11483 9373
rect 11425 9364 11437 9367
rect 11020 9336 11437 9364
rect 11020 9324 11026 9336
rect 11425 9333 11437 9336
rect 11471 9333 11483 9367
rect 12452 9364 12480 9404
rect 12693 9435 12707 9441
rect 12693 9401 12705 9435
rect 12759 9432 12765 9444
rect 12759 9404 12793 9432
rect 12693 9395 12707 9401
rect 12701 9392 12707 9395
rect 12759 9392 12765 9404
rect 13630 9392 13636 9444
rect 13688 9432 13694 9444
rect 14844 9432 14872 9528
rect 13688 9404 14872 9432
rect 13688 9392 13694 9404
rect 15378 9392 15384 9444
rect 15436 9432 15442 9444
rect 15841 9435 15899 9441
rect 15841 9432 15853 9435
rect 15436 9404 15853 9432
rect 15436 9392 15442 9404
rect 15841 9401 15853 9404
rect 15887 9401 15899 9435
rect 15841 9395 15899 9401
rect 12894 9364 12900 9376
rect 12452 9336 12900 9364
rect 11425 9327 11483 9333
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13780 9336 13829 9364
rect 13780 9324 13786 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 14826 9364 14832 9376
rect 14787 9336 14832 9364
rect 13817 9327 13875 9333
rect 14826 9324 14832 9336
rect 14884 9324 14890 9376
rect 15749 9367 15807 9373
rect 15749 9333 15761 9367
rect 15795 9364 15807 9367
rect 15930 9364 15936 9376
rect 15795 9336 15936 9364
rect 15795 9333 15807 9336
rect 15749 9327 15807 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 1104 9274 16836 9296
rect 1104 9222 6246 9274
rect 6298 9222 6310 9274
rect 6362 9222 6374 9274
rect 6426 9222 6438 9274
rect 6490 9222 11510 9274
rect 11562 9222 11574 9274
rect 11626 9222 11638 9274
rect 11690 9222 11702 9274
rect 11754 9222 16836 9274
rect 1104 9200 16836 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2130 9160 2136 9172
rect 2087 9132 2136 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 4246 9160 4252 9172
rect 3068 9132 4252 9160
rect 2314 8984 2320 9036
rect 2372 9024 2378 9036
rect 2409 9027 2467 9033
rect 2409 9024 2421 9027
rect 2372 8996 2421 9024
rect 2372 8984 2378 8996
rect 2409 8993 2421 8996
rect 2455 8993 2467 9027
rect 3068 9024 3096 9132
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 6917 9163 6975 9169
rect 6917 9160 6929 9163
rect 4396 9132 6929 9160
rect 4396 9120 4402 9132
rect 6917 9129 6929 9132
rect 6963 9129 6975 9163
rect 7282 9160 7288 9172
rect 7243 9132 7288 9160
rect 6917 9123 6975 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 7708 9132 8125 9160
rect 7708 9120 7714 9132
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 8113 9123 8171 9129
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 12434 9160 12440 9172
rect 8260 9132 12440 9160
rect 8260 9120 8266 9132
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9129 12587 9163
rect 12529 9123 12587 9129
rect 3142 9052 3148 9104
rect 3200 9092 3206 9104
rect 7098 9092 7104 9104
rect 3200 9064 7104 9092
rect 3200 9052 3206 9064
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 7208 9064 7604 9092
rect 3237 9027 3295 9033
rect 3237 9024 3249 9027
rect 3068 8996 3249 9024
rect 2409 8987 2467 8993
rect 3237 8993 3249 8996
rect 3283 8993 3295 9027
rect 3237 8987 3295 8993
rect 3326 8984 3332 9036
rect 3384 9024 3390 9036
rect 4065 9027 4123 9033
rect 3384 8996 4016 9024
rect 3384 8984 3390 8996
rect 3988 8968 4016 8996
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4154 9024 4160 9036
rect 4111 8996 4160 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 4246 8984 4252 9036
rect 4304 9024 4310 9036
rect 4890 9024 4896 9036
rect 4304 8996 4896 9024
rect 4304 8984 4310 8996
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8925 1455 8959
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 1397 8919 1455 8925
rect 1412 8888 1440 8919
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 3510 8956 3516 8968
rect 2731 8928 3516 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4798 8956 4804 8968
rect 4028 8928 4804 8956
rect 4028 8916 4034 8928
rect 4798 8916 4804 8928
rect 4856 8956 4862 8968
rect 5092 8956 5120 8987
rect 5166 8984 5172 9036
rect 5224 9024 5230 9036
rect 5333 9027 5391 9033
rect 5333 9024 5345 9027
rect 5224 8996 5345 9024
rect 5224 8984 5230 8996
rect 5333 8993 5345 8996
rect 5379 8993 5391 9027
rect 5333 8987 5391 8993
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 7208 9024 7236 9064
rect 5776 8996 7236 9024
rect 5776 8984 5782 8996
rect 4856 8928 5120 8956
rect 6472 8928 6684 8956
rect 4856 8916 4862 8928
rect 3142 8888 3148 8900
rect 1412 8860 3148 8888
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 3326 8848 3332 8900
rect 3384 8888 3390 8900
rect 5074 8888 5080 8900
rect 3384 8860 5080 8888
rect 3384 8848 3390 8860
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 6472 8897 6500 8928
rect 6457 8891 6515 8897
rect 6457 8857 6469 8891
rect 6503 8857 6515 8891
rect 6656 8888 6684 8928
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 6880 8928 7389 8956
rect 6880 8916 6886 8928
rect 7377 8925 7389 8928
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 7484 8888 7512 8919
rect 6656 8860 7512 8888
rect 7576 8888 7604 9064
rect 7742 9052 7748 9104
rect 7800 9092 7806 9104
rect 10321 9095 10379 9101
rect 10321 9092 10333 9095
rect 7800 9064 10333 9092
rect 7800 9052 7806 9064
rect 10321 9061 10333 9064
rect 10367 9092 10379 9095
rect 10410 9092 10416 9104
rect 10367 9064 10416 9092
rect 10367 9061 10379 9064
rect 10321 9055 10379 9061
rect 10410 9052 10416 9064
rect 10468 9052 10474 9104
rect 12544 9092 12572 9123
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12860 9132 13001 9160
rect 12860 9120 12866 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 13354 9160 13360 9172
rect 13315 9132 13360 9160
rect 12989 9123 13047 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 14918 9120 14924 9172
rect 14976 9160 14982 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 14976 9132 15669 9160
rect 14976 9120 14982 9132
rect 15657 9129 15669 9132
rect 15703 9129 15715 9163
rect 15657 9123 15715 9129
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 15804 9132 15849 9160
rect 15804 9120 15810 9132
rect 15194 9092 15200 9104
rect 12544 9064 15200 9092
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 8478 9024 8484 9036
rect 8439 8996 8484 9024
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 10962 9024 10968 9036
rect 9824 8996 10968 9024
rect 9824 8984 9830 8996
rect 10962 8984 10968 8996
rect 11020 9024 11026 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 11020 8996 11161 9024
rect 11020 8984 11026 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 11405 9027 11463 9033
rect 11405 9024 11417 9027
rect 11296 8996 11417 9024
rect 11296 8984 11302 8996
rect 11405 8993 11417 8996
rect 11451 8993 11463 9027
rect 11405 8987 11463 8993
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 14458 9024 14464 9036
rect 13412 8996 14464 9024
rect 13412 8984 13418 8996
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8573 8959 8631 8965
rect 8573 8956 8585 8959
rect 8352 8928 8585 8956
rect 8352 8916 8358 8928
rect 8573 8925 8585 8928
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9214 8956 9220 8968
rect 8803 8928 9220 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10428 8888 10456 8919
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 10560 8928 10605 8956
rect 10560 8916 10566 8928
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 13170 8956 13176 8968
rect 12492 8928 13176 8956
rect 12492 8916 12498 8928
rect 13170 8916 13176 8928
rect 13228 8956 13234 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 13228 8928 13461 8956
rect 13228 8916 13234 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 13596 8928 13641 8956
rect 13924 8928 15853 8956
rect 13596 8916 13602 8928
rect 7576 8860 10456 8888
rect 6457 8851 6515 8857
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2498 8820 2504 8832
rect 2372 8792 2504 8820
rect 2372 8780 2378 8792
rect 2498 8780 2504 8792
rect 2556 8780 2562 8832
rect 3418 8820 3424 8832
rect 3379 8792 3424 8820
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 4246 8820 4252 8832
rect 4207 8792 4252 8820
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 5258 8780 5264 8832
rect 5316 8820 5322 8832
rect 6472 8820 6500 8851
rect 9950 8820 9956 8832
rect 5316 8792 6500 8820
rect 9911 8792 9956 8820
rect 5316 8780 5322 8792
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 10428 8820 10456 8860
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 13814 8888 13820 8900
rect 12584 8860 13820 8888
rect 12584 8848 12590 8860
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 13262 8820 13268 8832
rect 10428 8792 13268 8820
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 13924 8820 13952 8928
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 13998 8848 14004 8900
rect 14056 8888 14062 8900
rect 15289 8891 15347 8897
rect 15289 8888 15301 8891
rect 14056 8860 15301 8888
rect 14056 8848 14062 8860
rect 15289 8857 15301 8860
rect 15335 8857 15347 8891
rect 15289 8851 15347 8857
rect 14642 8820 14648 8832
rect 13504 8792 13952 8820
rect 14603 8792 14648 8820
rect 13504 8780 13510 8792
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 1104 8730 16836 8752
rect 1104 8678 3614 8730
rect 3666 8678 3678 8730
rect 3730 8678 3742 8730
rect 3794 8678 3806 8730
rect 3858 8678 8878 8730
rect 8930 8678 8942 8730
rect 8994 8678 9006 8730
rect 9058 8678 9070 8730
rect 9122 8678 14142 8730
rect 14194 8678 14206 8730
rect 14258 8678 14270 8730
rect 14322 8678 14334 8730
rect 14386 8678 16836 8730
rect 1104 8656 16836 8678
rect 3326 8616 3332 8628
rect 1412 8588 3332 8616
rect 1412 8421 1440 8588
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3510 8616 3516 8628
rect 3471 8588 3516 8616
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 5353 8619 5411 8625
rect 5353 8616 5365 8619
rect 3896 8588 5365 8616
rect 3896 8560 3924 8588
rect 5353 8585 5365 8588
rect 5399 8585 5411 8619
rect 6822 8616 6828 8628
rect 6783 8588 6828 8616
rect 5353 8579 5411 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 13354 8616 13360 8628
rect 7156 8588 13360 8616
rect 7156 8576 7162 8588
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 3878 8508 3884 8560
rect 3936 8508 3942 8560
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 7926 8548 7932 8560
rect 5040 8520 7932 8548
rect 5040 8508 5046 8520
rect 7926 8508 7932 8520
rect 7984 8508 7990 8560
rect 9858 8548 9864 8560
rect 9819 8520 9864 8548
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 11057 8551 11115 8557
rect 11057 8517 11069 8551
rect 11103 8517 11115 8551
rect 11057 8511 11115 8517
rect 3970 8480 3976 8492
rect 3931 8452 3976 8480
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 7374 8480 7380 8492
rect 5224 8452 7380 8480
rect 5224 8440 5230 8452
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 10502 8480 10508 8492
rect 10463 8452 10508 8480
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 11072 8480 11100 8511
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 12952 8520 14044 8548
rect 12952 8508 12958 8520
rect 11146 8480 11152 8492
rect 11072 8452 11152 8480
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11330 8440 11336 8492
rect 11388 8480 11394 8492
rect 11609 8483 11667 8489
rect 11609 8480 11621 8483
rect 11388 8452 11621 8480
rect 11388 8440 11394 8452
rect 11609 8449 11621 8452
rect 11655 8449 11667 8483
rect 13262 8480 13268 8492
rect 13223 8452 13268 8480
rect 11609 8443 11667 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 14016 8489 14044 8520
rect 15102 8508 15108 8560
rect 15160 8548 15166 8560
rect 16025 8551 16083 8557
rect 16025 8548 16037 8551
rect 15160 8520 16037 8548
rect 15160 8508 15166 8520
rect 16025 8517 16037 8520
rect 16071 8517 16083 8551
rect 16025 8511 16083 8517
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8480 13507 8483
rect 14001 8483 14059 8489
rect 13495 8452 13768 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8412 2191 8415
rect 3988 8412 4016 8440
rect 2179 8384 4016 8412
rect 4240 8415 4298 8421
rect 2179 8381 2191 8384
rect 2133 8375 2191 8381
rect 4240 8381 4252 8415
rect 4286 8412 4298 8415
rect 5258 8412 5264 8424
rect 4286 8384 5264 8412
rect 4286 8381 4298 8384
rect 4240 8375 4298 8381
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8412 5871 8415
rect 7190 8412 7196 8424
rect 5859 8384 7196 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8412 8079 8415
rect 9766 8412 9772 8424
rect 8067 8384 9772 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 10229 8415 10287 8421
rect 10229 8381 10241 8415
rect 10275 8412 10287 8415
rect 10318 8412 10324 8424
rect 10275 8384 10324 8412
rect 10275 8381 10287 8384
rect 10229 8375 10287 8381
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 10836 8384 11437 8412
rect 10836 8372 10842 8384
rect 11425 8381 11437 8384
rect 11471 8412 11483 8415
rect 13354 8412 13360 8424
rect 11471 8384 13360 8412
rect 11471 8381 11483 8384
rect 11425 8375 11483 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 13740 8356 13768 8452
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 13814 8372 13820 8424
rect 13872 8412 13878 8424
rect 15838 8412 15844 8424
rect 13872 8384 14412 8412
rect 15799 8384 15844 8412
rect 13872 8372 13878 8384
rect 2400 8347 2458 8353
rect 2400 8313 2412 8347
rect 2446 8344 2458 8347
rect 3878 8344 3884 8356
rect 2446 8316 3884 8344
rect 2446 8313 2458 8316
rect 2400 8307 2458 8313
rect 3878 8304 3884 8316
rect 3936 8304 3942 8356
rect 4356 8316 6040 8344
rect 1578 8276 1584 8288
rect 1539 8248 1584 8276
rect 1578 8236 1584 8248
rect 1636 8236 1642 8288
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 4356 8276 4384 8316
rect 6012 8285 6040 8316
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 6972 8316 7297 8344
rect 6972 8304 6978 8316
rect 7285 8313 7297 8316
rect 7331 8344 7343 8347
rect 8110 8344 8116 8356
rect 7331 8316 8116 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 8288 8347 8346 8353
rect 8288 8313 8300 8347
rect 8334 8344 8346 8347
rect 9030 8344 9036 8356
rect 8334 8316 9036 8344
rect 8334 8313 8346 8316
rect 8288 8307 8346 8313
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 9916 8316 10364 8344
rect 9916 8304 9922 8316
rect 4028 8248 4384 8276
rect 5997 8279 6055 8285
rect 4028 8236 4034 8248
rect 5997 8245 6009 8279
rect 6043 8245 6055 8279
rect 5997 8239 6055 8245
rect 7098 8236 7104 8288
rect 7156 8276 7162 8288
rect 7193 8279 7251 8285
rect 7193 8276 7205 8279
rect 7156 8248 7205 8276
rect 7156 8236 7162 8248
rect 7193 8245 7205 8248
rect 7239 8245 7251 8279
rect 7193 8239 7251 8245
rect 9401 8279 9459 8285
rect 9401 8245 9413 8279
rect 9447 8276 9459 8279
rect 9582 8276 9588 8288
rect 9447 8248 9588 8276
rect 9447 8245 9459 8248
rect 9401 8239 9459 8245
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 10336 8285 10364 8316
rect 11514 8304 11520 8356
rect 11572 8344 11578 8356
rect 11572 8316 11617 8344
rect 11572 8304 11578 8316
rect 13078 8304 13084 8356
rect 13136 8344 13142 8356
rect 13173 8347 13231 8353
rect 13173 8344 13185 8347
rect 13136 8316 13185 8344
rect 13136 8304 13142 8316
rect 13173 8313 13185 8316
rect 13219 8313 13231 8347
rect 13173 8307 13231 8313
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 14246 8347 14304 8353
rect 14246 8344 14258 8347
rect 13780 8316 14258 8344
rect 13780 8304 13786 8316
rect 14246 8313 14258 8316
rect 14292 8313 14304 8347
rect 14384 8344 14412 8384
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 16114 8344 16120 8356
rect 14384 8316 16120 8344
rect 14246 8307 14304 8313
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 10321 8279 10379 8285
rect 10321 8245 10333 8279
rect 10367 8245 10379 8279
rect 10321 8239 10379 8245
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 12618 8276 12624 8288
rect 10468 8248 12624 8276
rect 10468 8236 10474 8248
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 12802 8276 12808 8288
rect 12763 8248 12808 8276
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 15381 8279 15439 8285
rect 15381 8245 15393 8279
rect 15427 8276 15439 8279
rect 15838 8276 15844 8288
rect 15427 8248 15844 8276
rect 15427 8245 15439 8248
rect 15381 8239 15439 8245
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 1104 8186 16836 8208
rect 1104 8134 6246 8186
rect 6298 8134 6310 8186
rect 6362 8134 6374 8186
rect 6426 8134 6438 8186
rect 6490 8134 11510 8186
rect 11562 8134 11574 8186
rect 11626 8134 11638 8186
rect 11690 8134 11702 8186
rect 11754 8134 16836 8186
rect 1104 8112 16836 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 1995 8044 2789 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 3142 8072 3148 8084
rect 3103 8044 3148 8072
rect 2777 8035 2835 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 6733 8075 6791 8081
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 7282 8072 7288 8084
rect 6779 8044 7288 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7650 8072 7656 8084
rect 7524 8044 7656 8072
rect 7524 8032 7530 8044
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 8849 8075 8907 8081
rect 8849 8072 8861 8075
rect 8812 8044 8861 8072
rect 8812 8032 8818 8044
rect 8849 8041 8861 8044
rect 8895 8041 8907 8075
rect 8849 8035 8907 8041
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 10008 8044 10149 8072
rect 10008 8032 10014 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10226 8032 10232 8084
rect 10284 8072 10290 8084
rect 12434 8072 12440 8084
rect 10284 8044 10329 8072
rect 10428 8044 12440 8072
rect 10284 8032 10290 8044
rect 3237 8007 3295 8013
rect 3237 7973 3249 8007
rect 3283 8004 3295 8007
rect 10428 8004 10456 8044
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 12802 8072 12808 8084
rect 12575 8044 12808 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 13725 8075 13783 8081
rect 13725 8041 13737 8075
rect 13771 8072 13783 8075
rect 14090 8072 14096 8084
rect 13771 8044 14096 8072
rect 13771 8041 13783 8044
rect 13725 8035 13783 8041
rect 3283 7976 10456 8004
rect 3283 7973 3295 7976
rect 3237 7967 3295 7973
rect 3142 7896 3148 7948
rect 3200 7936 3206 7948
rect 4062 7936 4068 7948
rect 3200 7908 4068 7936
rect 3200 7896 3206 7908
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4890 7936 4896 7948
rect 4851 7908 4896 7936
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 5736 7945 5764 7976
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 11333 8007 11391 8013
rect 11333 8004 11345 8007
rect 11112 7976 11345 8004
rect 11112 7964 11118 7976
rect 11333 7973 11345 7976
rect 11379 8004 11391 8007
rect 11514 8004 11520 8016
rect 11379 7976 11520 8004
rect 11379 7973 11391 7976
rect 11333 7967 11391 7973
rect 11514 7964 11520 7976
rect 11572 7964 11578 8016
rect 11698 7964 11704 8016
rect 11756 8004 11762 8016
rect 12618 8004 12624 8016
rect 11756 7976 12624 8004
rect 11756 7964 11762 7976
rect 12618 7964 12624 7976
rect 12676 8004 12682 8016
rect 13740 8004 13768 8035
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 14458 8032 14464 8084
rect 14516 8072 14522 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 14516 8044 15669 8072
rect 14516 8032 14522 8044
rect 15657 8041 15669 8044
rect 15703 8041 15715 8075
rect 15657 8035 15715 8041
rect 15749 8075 15807 8081
rect 15749 8041 15761 8075
rect 15795 8072 15807 8075
rect 16114 8072 16120 8084
rect 15795 8044 16120 8072
rect 15795 8041 15807 8044
rect 15749 8035 15807 8041
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 14734 8004 14740 8016
rect 12676 7976 13768 8004
rect 13832 7976 14740 8004
rect 12676 7964 12682 7976
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7905 5779 7939
rect 6638 7936 6644 7948
rect 6599 7908 6644 7936
rect 5721 7899 5779 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 7098 7936 7104 7948
rect 7059 7908 7104 7936
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 10134 7936 10140 7948
rect 8803 7908 10140 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 10134 7896 10140 7908
rect 10192 7896 10198 7948
rect 11425 7939 11483 7945
rect 11425 7905 11437 7939
rect 11471 7936 11483 7939
rect 11606 7936 11612 7948
rect 11471 7908 11612 7936
rect 11471 7905 11483 7908
rect 11425 7899 11483 7905
rect 11606 7896 11612 7908
rect 11664 7936 11670 7948
rect 13832 7936 13860 7976
rect 14734 7964 14740 7976
rect 14792 7964 14798 8016
rect 14826 7964 14832 8016
rect 14884 8004 14890 8016
rect 15470 8004 15476 8016
rect 14884 7976 15476 8004
rect 14884 7964 14890 7976
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 11664 7908 13860 7936
rect 11664 7896 11670 7908
rect 2038 7868 2044 7880
rect 1999 7840 2044 7868
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7868 2283 7871
rect 2682 7868 2688 7880
rect 2271 7840 2688 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 3326 7868 3332 7880
rect 3287 7840 3332 7868
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 4982 7868 4988 7880
rect 4943 7840 4988 7868
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5258 7868 5264 7880
rect 5215 7840 5264 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 7190 7868 7196 7880
rect 7103 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7374 7868 7380 7880
rect 7335 7840 7380 7868
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 9030 7868 9036 7880
rect 8943 7840 9036 7868
rect 9030 7828 9036 7840
rect 9088 7868 9094 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 9088 7840 10425 7868
rect 9088 7828 9094 7840
rect 10413 7837 10425 7840
rect 10459 7868 10471 7871
rect 11330 7868 11336 7880
rect 10459 7840 11336 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 11330 7828 11336 7840
rect 11388 7868 11394 7880
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 11388 7840 11529 7868
rect 11388 7828 11394 7840
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 12621 7871 12679 7877
rect 12621 7837 12633 7871
rect 12667 7837 12679 7871
rect 12802 7868 12808 7880
rect 12763 7840 12808 7868
rect 12621 7831 12679 7837
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 5905 7803 5963 7809
rect 5905 7800 5917 7803
rect 4120 7772 5917 7800
rect 4120 7760 4126 7772
rect 5905 7769 5917 7772
rect 5951 7769 5963 7803
rect 7208 7800 7236 7828
rect 12526 7800 12532 7812
rect 7208 7772 12532 7800
rect 5905 7763 5963 7769
rect 12526 7760 12532 7772
rect 12584 7760 12590 7812
rect 12636 7800 12664 7831
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 13817 7871 13875 7877
rect 13817 7868 13829 7871
rect 13044 7840 13829 7868
rect 13044 7828 13050 7840
rect 13817 7837 13829 7840
rect 13863 7837 13875 7871
rect 13817 7831 13875 7837
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7837 13967 7871
rect 14550 7868 14556 7880
rect 14511 7840 14556 7868
rect 13909 7831 13967 7837
rect 13357 7803 13415 7809
rect 13357 7800 13369 7803
rect 12636 7772 13369 7800
rect 13357 7769 13369 7772
rect 13403 7769 13415 7803
rect 13357 7763 13415 7769
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 13924 7800 13952 7831
rect 14550 7828 14556 7840
rect 14608 7828 14614 7880
rect 15838 7868 15844 7880
rect 15799 7840 15844 7868
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 17218 7800 17224 7812
rect 13780 7772 13952 7800
rect 14016 7772 17224 7800
rect 13780 7760 13786 7772
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2314 7732 2320 7744
rect 1627 7704 2320 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2314 7692 2320 7704
rect 2372 7692 2378 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 4525 7735 4583 7741
rect 4525 7732 4537 7735
rect 4212 7704 4537 7732
rect 4212 7692 4218 7704
rect 4525 7701 4537 7704
rect 4571 7701 4583 7735
rect 4525 7695 4583 7701
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 6457 7735 6515 7741
rect 6457 7732 6469 7735
rect 5408 7704 6469 7732
rect 5408 7692 5414 7704
rect 6457 7701 6469 7704
rect 6503 7701 6515 7735
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 6457 7695 6515 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 9766 7732 9772 7744
rect 9727 7704 9772 7732
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 12161 7735 12219 7741
rect 12161 7732 12173 7735
rect 11940 7704 12173 7732
rect 11940 7692 11946 7704
rect 12161 7701 12173 7704
rect 12207 7701 12219 7735
rect 12161 7695 12219 7701
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 14016 7732 14044 7772
rect 17218 7760 17224 7772
rect 17276 7760 17282 7812
rect 12308 7704 14044 7732
rect 12308 7692 12314 7704
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 15289 7735 15347 7741
rect 15289 7732 15301 7735
rect 15252 7704 15301 7732
rect 15252 7692 15258 7704
rect 15289 7701 15301 7704
rect 15335 7701 15347 7735
rect 15289 7695 15347 7701
rect 1104 7642 16836 7664
rect 1104 7590 3614 7642
rect 3666 7590 3678 7642
rect 3730 7590 3742 7642
rect 3794 7590 3806 7642
rect 3858 7590 8878 7642
rect 8930 7590 8942 7642
rect 8994 7590 9006 7642
rect 9058 7590 9070 7642
rect 9122 7590 14142 7642
rect 14194 7590 14206 7642
rect 14258 7590 14270 7642
rect 14322 7590 14334 7642
rect 14386 7590 16836 7642
rect 1104 7568 16836 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2501 7531 2559 7537
rect 2501 7528 2513 7531
rect 2096 7500 2513 7528
rect 2096 7488 2102 7500
rect 2501 7497 2513 7500
rect 2547 7497 2559 7531
rect 4890 7528 4896 7540
rect 2501 7491 2559 7497
rect 2976 7500 4752 7528
rect 4851 7500 4896 7528
rect 2976 7460 3004 7500
rect 1504 7432 3004 7460
rect 1504 7324 1532 7432
rect 2590 7352 2596 7404
rect 2648 7392 2654 7404
rect 2976 7401 3004 7432
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 4028 7432 4292 7460
rect 4028 7420 4034 7432
rect 2961 7395 3019 7401
rect 2648 7364 2912 7392
rect 2648 7352 2654 7364
rect 2884 7333 2912 7364
rect 2961 7361 2973 7395
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 3326 7392 3332 7404
rect 3191 7364 3332 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 4154 7392 4160 7404
rect 4115 7364 4160 7392
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4264 7401 4292 7432
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 1569 7327 1627 7333
rect 1569 7324 1581 7327
rect 1504 7296 1581 7324
rect 1569 7293 1581 7296
rect 1615 7293 1627 7327
rect 1569 7287 1627 7293
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7293 2927 7327
rect 2869 7287 2927 7293
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 3970 7324 3976 7336
rect 3108 7296 3976 7324
rect 3108 7284 3114 7296
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4065 7327 4123 7333
rect 4065 7293 4077 7327
rect 4111 7324 4123 7327
rect 4338 7324 4344 7336
rect 4111 7296 4344 7324
rect 4111 7293 4123 7296
rect 4065 7287 4123 7293
rect 4338 7284 4344 7296
rect 4396 7284 4402 7336
rect 4724 7324 4752 7500
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 6638 7488 6644 7540
rect 6696 7528 6702 7540
rect 9401 7531 9459 7537
rect 9401 7528 9413 7531
rect 6696 7500 9413 7528
rect 6696 7488 6702 7500
rect 9401 7497 9413 7500
rect 9447 7528 9459 7531
rect 9674 7528 9680 7540
rect 9447 7500 9680 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 12250 7528 12256 7540
rect 9784 7500 12256 7528
rect 5810 7420 5816 7472
rect 5868 7460 5874 7472
rect 9784 7460 9812 7500
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 13817 7531 13875 7537
rect 13817 7528 13829 7531
rect 12452 7500 13829 7528
rect 5868 7432 7236 7460
rect 5868 7420 5874 7432
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 5224 7364 5457 7392
rect 5224 7352 5230 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 6089 7395 6147 7401
rect 6089 7361 6101 7395
rect 6135 7392 6147 7395
rect 7098 7392 7104 7404
rect 6135 7364 7104 7392
rect 6135 7361 6147 7364
rect 6089 7355 6147 7361
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7208 7324 7236 7432
rect 8128 7432 9812 7460
rect 11425 7463 11483 7469
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 4724 7296 6960 7324
rect 7208 7296 7297 7324
rect 5353 7259 5411 7265
rect 1780 7228 2636 7256
rect 1780 7197 1808 7228
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7157 1823 7191
rect 2608 7188 2636 7228
rect 5353 7225 5365 7259
rect 5399 7256 5411 7259
rect 6932 7256 6960 7296
rect 7285 7293 7297 7296
rect 7331 7324 7343 7327
rect 7926 7324 7932 7336
rect 7331 7296 7932 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8128 7333 8156 7432
rect 11425 7429 11437 7463
rect 11471 7460 11483 7463
rect 12342 7460 12348 7472
rect 11471 7432 12348 7460
rect 11471 7429 11483 7432
rect 11425 7423 11483 7429
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 11882 7392 11888 7404
rect 8536 7364 10088 7392
rect 11843 7364 11888 7392
rect 8536 7352 8542 7364
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7293 8171 7327
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 8113 7287 8171 7293
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 10060 7324 10088 7364
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7392 12127 7395
rect 12452 7392 12480 7500
rect 13817 7497 13829 7500
rect 13863 7528 13875 7531
rect 13906 7528 13912 7540
rect 13863 7500 13912 7528
rect 13863 7497 13875 7500
rect 13817 7491 13875 7497
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 12115 7364 12480 7392
rect 12115 7361 12127 7364
rect 12069 7355 12127 7361
rect 13722 7352 13728 7404
rect 13780 7392 13786 7404
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 13780 7364 14841 7392
rect 13780 7352 13786 7364
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 11698 7324 11704 7336
rect 10060 7296 11704 7324
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 12710 7333 12716 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12400 7296 12449 7324
rect 12400 7284 12406 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 12704 7287 12716 7333
rect 12768 7324 12774 7336
rect 12768 7296 12804 7324
rect 12710 7284 12716 7287
rect 12768 7284 12774 7296
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 15841 7327 15899 7333
rect 15841 7324 15853 7327
rect 13228 7296 15853 7324
rect 13228 7284 13234 7296
rect 15841 7293 15853 7296
rect 15887 7293 15899 7327
rect 15841 7287 15899 7293
rect 5399 7228 6868 7256
rect 6932 7228 7328 7256
rect 5399 7225 5411 7228
rect 5353 7219 5411 7225
rect 2866 7188 2872 7200
rect 2608 7160 2872 7188
rect 1765 7151 1823 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 3568 7160 3709 7188
rect 3568 7148 3574 7160
rect 3697 7157 3709 7160
rect 3743 7157 3755 7191
rect 3697 7151 3755 7157
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4764 7160 5273 7188
rect 4764 7148 4770 7160
rect 5261 7157 5273 7160
rect 5307 7188 5319 7191
rect 6730 7188 6736 7200
rect 5307 7160 6736 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 6840 7197 6868 7228
rect 6825 7191 6883 7197
rect 6825 7157 6837 7191
rect 6871 7157 6883 7191
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 6825 7151 6883 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7300 7188 7328 7228
rect 9582 7216 9588 7268
rect 9640 7256 9646 7268
rect 10198 7259 10256 7265
rect 10198 7256 10210 7259
rect 9640 7228 10210 7256
rect 9640 7216 9646 7228
rect 10198 7225 10210 7228
rect 10244 7225 10256 7259
rect 10198 7219 10256 7225
rect 11793 7259 11851 7265
rect 11793 7225 11805 7259
rect 11839 7256 11851 7259
rect 11839 7228 12112 7256
rect 11839 7225 11851 7228
rect 11793 7219 11851 7225
rect 10410 7188 10416 7200
rect 7300 7160 10416 7188
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11112 7160 11345 7188
rect 11112 7148 11118 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 12084 7188 12112 7228
rect 12526 7216 12532 7268
rect 12584 7256 12590 7268
rect 14366 7256 14372 7268
rect 12584 7228 14372 7256
rect 12584 7216 12590 7228
rect 14366 7216 14372 7228
rect 14424 7216 14430 7268
rect 14737 7259 14795 7265
rect 14737 7225 14749 7259
rect 14783 7256 14795 7259
rect 15010 7256 15016 7268
rect 14783 7228 15016 7256
rect 14783 7225 14795 7228
rect 14737 7219 14795 7225
rect 15010 7216 15016 7228
rect 15068 7216 15074 7268
rect 13170 7188 13176 7200
rect 12084 7160 13176 7188
rect 11333 7151 11391 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 14274 7188 14280 7200
rect 14235 7160 14280 7188
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 14645 7191 14703 7197
rect 14645 7157 14657 7191
rect 14691 7188 14703 7191
rect 14826 7188 14832 7200
rect 14691 7160 14832 7188
rect 14691 7157 14703 7160
rect 14645 7151 14703 7157
rect 14826 7148 14832 7160
rect 14884 7148 14890 7200
rect 16022 7188 16028 7200
rect 15983 7160 16028 7188
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 1104 7098 16836 7120
rect 1104 7046 6246 7098
rect 6298 7046 6310 7098
rect 6362 7046 6374 7098
rect 6426 7046 6438 7098
rect 6490 7046 11510 7098
rect 11562 7046 11574 7098
rect 11626 7046 11638 7098
rect 11690 7046 11702 7098
rect 11754 7046 16836 7098
rect 1104 7024 16836 7046
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 3050 6984 3056 6996
rect 2832 6956 3056 6984
rect 2832 6944 2838 6956
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5077 6987 5135 6993
rect 5077 6984 5089 6987
rect 5040 6956 5089 6984
rect 5040 6944 5046 6956
rect 5077 6953 5089 6956
rect 5123 6953 5135 6987
rect 6914 6984 6920 6996
rect 5077 6947 5135 6953
rect 5184 6956 6920 6984
rect 3326 6916 3332 6928
rect 2608 6888 3332 6916
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 2400 6851 2458 6857
rect 2400 6817 2412 6851
rect 2446 6848 2458 6851
rect 2608 6848 2636 6888
rect 3326 6876 3332 6888
rect 3384 6876 3390 6928
rect 5184 6916 5212 6956
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 7653 6987 7711 6993
rect 7653 6984 7665 6987
rect 7524 6956 7665 6984
rect 7524 6944 7530 6956
rect 7653 6953 7665 6956
rect 7699 6953 7711 6987
rect 7653 6947 7711 6953
rect 7926 6944 7932 6996
rect 7984 6984 7990 6996
rect 12894 6984 12900 6996
rect 7984 6956 12900 6984
rect 7984 6944 7990 6956
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 13170 6984 13176 6996
rect 13131 6956 13176 6984
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 14550 6944 14556 6996
rect 14608 6984 14614 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 14608 6956 15669 6984
rect 14608 6944 14614 6956
rect 15657 6953 15669 6956
rect 15703 6953 15715 6987
rect 15657 6947 15715 6953
rect 4908 6888 5212 6916
rect 5445 6919 5503 6925
rect 2446 6820 2636 6848
rect 2446 6817 2458 6820
rect 2400 6811 2458 6817
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 4065 6851 4123 6857
rect 2740 6820 3556 6848
rect 2740 6808 2746 6820
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 3528 6721 3556 6820
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4908 6848 4936 6888
rect 5445 6885 5457 6919
rect 5491 6916 5503 6919
rect 5491 6888 6868 6916
rect 5491 6885 5503 6888
rect 5445 6879 5503 6885
rect 4111 6820 4936 6848
rect 4985 6851 5043 6857
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4985 6817 4997 6851
rect 5031 6848 5043 6851
rect 5350 6848 5356 6860
rect 5031 6820 5356 6848
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 6529 6851 6587 6857
rect 6529 6848 6541 6851
rect 5868 6820 6541 6848
rect 5868 6808 5874 6820
rect 6529 6817 6541 6820
rect 6575 6817 6587 6851
rect 6840 6848 6868 6888
rect 7006 6876 7012 6928
rect 7064 6916 7070 6928
rect 13541 6919 13599 6925
rect 13541 6916 13553 6919
rect 7064 6888 13553 6916
rect 7064 6876 7070 6888
rect 13541 6885 13553 6888
rect 13587 6916 13599 6919
rect 13814 6916 13820 6928
rect 13587 6888 13820 6916
rect 13587 6885 13599 6888
rect 13541 6879 13599 6885
rect 13814 6876 13820 6888
rect 13872 6876 13878 6928
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 15749 6919 15807 6925
rect 15749 6916 15761 6919
rect 14424 6888 15761 6916
rect 14424 6876 14430 6888
rect 15749 6885 15761 6888
rect 15795 6885 15807 6919
rect 15749 6879 15807 6885
rect 6840 6820 7328 6848
rect 6529 6811 6587 6817
rect 5534 6780 5540 6792
rect 5495 6752 5540 6780
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 3513 6715 3571 6721
rect 3513 6681 3525 6715
rect 3559 6681 3571 6715
rect 3513 6675 3571 6681
rect 5166 6672 5172 6724
rect 5224 6712 5230 6724
rect 5644 6712 5672 6743
rect 5224 6684 5672 6712
rect 5224 6672 5230 6684
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2774 6644 2780 6656
rect 1627 6616 2780 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 4249 6647 4307 6653
rect 4249 6644 4261 6647
rect 4212 6616 4261 6644
rect 4212 6604 4218 6616
rect 4249 6613 4261 6616
rect 4295 6613 4307 6647
rect 4249 6607 4307 6613
rect 4430 6604 4436 6656
rect 4488 6644 4494 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4488 6616 4813 6644
rect 4488 6604 4494 6616
rect 4801 6613 4813 6616
rect 4847 6644 4859 6647
rect 5442 6644 5448 6656
rect 4847 6616 5448 6644
rect 4847 6613 4859 6616
rect 4801 6607 4859 6613
rect 5442 6604 5448 6616
rect 5500 6644 5506 6656
rect 6288 6644 6316 6743
rect 7300 6712 7328 6820
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 8260 6820 8493 6848
rect 8260 6808 8266 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 9950 6848 9956 6860
rect 8987 6820 9956 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10134 6848 10140 6860
rect 10095 6820 10140 6848
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 11054 6857 11060 6860
rect 11048 6848 11060 6857
rect 11015 6820 11060 6848
rect 11048 6811 11060 6820
rect 11054 6808 11060 6811
rect 11112 6808 11118 6860
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6848 13691 6851
rect 14274 6848 14280 6860
rect 13679 6820 14280 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 14458 6848 14464 6860
rect 14419 6820 14464 6848
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 8757 6783 8815 6789
rect 8628 6752 8673 6780
rect 8628 6740 8634 6752
rect 8757 6749 8769 6783
rect 8803 6749 8815 6783
rect 9214 6780 9220 6792
rect 9175 6752 9220 6780
rect 8757 6743 8815 6749
rect 8113 6715 8171 6721
rect 8113 6712 8125 6715
rect 7300 6684 8125 6712
rect 8113 6681 8125 6684
rect 8159 6681 8171 6715
rect 8113 6675 8171 6681
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 8772 6712 8800 6743
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10100 6752 10793 6780
rect 10100 6740 10106 6752
rect 10781 6749 10793 6752
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 12802 6740 12808 6792
rect 12860 6780 12866 6792
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 12860 6752 13829 6780
rect 12860 6740 12866 6752
rect 13817 6749 13829 6752
rect 13863 6780 13875 6783
rect 15838 6780 15844 6792
rect 13863 6752 15844 6780
rect 13863 6749 13875 6752
rect 13817 6743 13875 6749
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 14642 6712 14648 6724
rect 8720 6684 8800 6712
rect 14603 6684 14648 6712
rect 8720 6672 8726 6684
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 5500 6616 6316 6644
rect 5500 6604 5506 6616
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 9858 6644 9864 6656
rect 9456 6616 9864 6644
rect 9456 6604 9462 6616
rect 9858 6604 9864 6616
rect 9916 6644 9922 6656
rect 10410 6644 10416 6656
rect 9916 6616 10416 6644
rect 9916 6604 9922 6616
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 12161 6647 12219 6653
rect 12161 6613 12173 6647
rect 12207 6644 12219 6647
rect 12526 6644 12532 6656
rect 12207 6616 12532 6644
rect 12207 6613 12219 6616
rect 12161 6607 12219 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 15286 6644 15292 6656
rect 15247 6616 15292 6644
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 1104 6554 16836 6576
rect 1104 6502 3614 6554
rect 3666 6502 3678 6554
rect 3730 6502 3742 6554
rect 3794 6502 3806 6554
rect 3858 6502 8878 6554
rect 8930 6502 8942 6554
rect 8994 6502 9006 6554
rect 9058 6502 9070 6554
rect 9122 6502 14142 6554
rect 14194 6502 14206 6554
rect 14258 6502 14270 6554
rect 14322 6502 14334 6554
rect 14386 6502 16836 6554
rect 1104 6480 16836 6502
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 5592 6412 6837 6440
rect 5592 6400 5598 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 8478 6440 8484 6452
rect 6972 6412 8484 6440
rect 6972 6400 6978 6412
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 8680 6412 11100 6440
rect 5810 6372 5816 6384
rect 5771 6344 5816 6372
rect 5810 6332 5816 6344
rect 5868 6332 5874 6384
rect 6638 6332 6644 6384
rect 6696 6372 6702 6384
rect 8680 6372 8708 6412
rect 6696 6344 8708 6372
rect 8757 6375 8815 6381
rect 6696 6332 6702 6344
rect 8757 6341 8769 6375
rect 8803 6372 8815 6375
rect 9858 6372 9864 6384
rect 8803 6344 9864 6372
rect 8803 6341 8815 6344
rect 8757 6335 8815 6341
rect 9858 6332 9864 6344
rect 9916 6332 9922 6384
rect 5828 6304 5856 6332
rect 7374 6304 7380 6316
rect 5828 6276 7380 6304
rect 7374 6264 7380 6276
rect 7432 6304 7438 6316
rect 8662 6304 8668 6316
rect 7432 6276 8668 6304
rect 7432 6264 7438 6276
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9582 6304 9588 6316
rect 9447 6276 9588 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 11072 6304 11100 6412
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 11333 6443 11391 6449
rect 11333 6440 11345 6443
rect 11296 6412 11345 6440
rect 11296 6400 11302 6412
rect 11333 6409 11345 6412
rect 11379 6409 11391 6443
rect 11790 6440 11796 6452
rect 11751 6412 11796 6440
rect 11333 6403 11391 6409
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 16025 6443 16083 6449
rect 16025 6409 16037 6443
rect 16071 6440 16083 6443
rect 16114 6440 16120 6452
rect 16071 6412 16120 6440
rect 16071 6409 16083 6412
rect 16025 6403 16083 6409
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 9732 6276 10088 6304
rect 11072 6276 12103 6304
rect 9732 6264 9738 6276
rect 1670 6236 1676 6248
rect 1631 6208 1676 6236
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 2130 6196 2136 6248
rect 2188 6236 2194 6248
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2188 6208 2605 6236
rect 2188 6196 2194 6208
rect 2593 6205 2605 6208
rect 2639 6236 2651 6239
rect 4430 6236 4436 6248
rect 2639 6208 4436 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 9217 6239 9275 6245
rect 9217 6205 9229 6239
rect 9263 6236 9275 6239
rect 9766 6236 9772 6248
rect 9263 6208 9772 6236
rect 9263 6205 9275 6208
rect 9217 6199 9275 6205
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6205 10011 6239
rect 10060 6236 10088 6276
rect 11977 6239 12035 6245
rect 11977 6236 11989 6239
rect 10060 6208 11989 6236
rect 9953 6199 10011 6205
rect 11977 6205 11989 6208
rect 12023 6205 12035 6239
rect 11977 6199 12035 6205
rect 1949 6171 2007 6177
rect 1949 6137 1961 6171
rect 1995 6168 2007 6171
rect 2222 6168 2228 6180
rect 1995 6140 2228 6168
rect 1995 6137 2007 6140
rect 1949 6131 2007 6137
rect 2222 6128 2228 6140
rect 2280 6128 2286 6180
rect 2682 6128 2688 6180
rect 2740 6168 2746 6180
rect 2838 6171 2896 6177
rect 2838 6168 2850 6171
rect 2740 6140 2850 6168
rect 2740 6128 2746 6140
rect 2838 6137 2850 6140
rect 2884 6137 2896 6171
rect 4678 6171 4736 6177
rect 4678 6168 4690 6171
rect 2838 6131 2896 6137
rect 3988 6140 4690 6168
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 3988 6109 4016 6140
rect 4678 6137 4690 6140
rect 4724 6137 4736 6171
rect 4678 6131 4736 6137
rect 4890 6128 4896 6180
rect 4948 6168 4954 6180
rect 9398 6168 9404 6180
rect 4948 6140 9404 6168
rect 4948 6128 4954 6140
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 9968 6168 9996 6199
rect 12075 6180 12103 6276
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12492 6276 12909 6304
rect 12492 6264 12498 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6304 13139 6307
rect 13127 6276 13768 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 12342 6196 12348 6248
rect 12400 6236 12406 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 12400 6208 13645 6236
rect 12400 6196 12406 6208
rect 13633 6205 13645 6208
rect 13679 6205 13691 6239
rect 13633 6199 13691 6205
rect 10042 6168 10048 6180
rect 9548 6140 10048 6168
rect 9548 6128 9554 6140
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 10226 6177 10232 6180
rect 10220 6168 10232 6177
rect 10187 6140 10232 6168
rect 10220 6131 10232 6140
rect 10226 6128 10232 6131
rect 10284 6128 10290 6180
rect 12066 6168 12072 6180
rect 11979 6140 12072 6168
rect 12066 6128 12072 6140
rect 12124 6168 12130 6180
rect 13740 6168 13768 6276
rect 13906 6245 13912 6248
rect 13900 6236 13912 6245
rect 13867 6208 13912 6236
rect 13900 6199 13912 6208
rect 13906 6196 13912 6199
rect 13964 6196 13970 6248
rect 14182 6196 14188 6248
rect 14240 6236 14246 6248
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 14240 6208 15853 6236
rect 14240 6196 14246 6208
rect 15841 6205 15853 6208
rect 15887 6205 15899 6239
rect 15841 6199 15899 6205
rect 12124 6140 12940 6168
rect 13740 6140 15056 6168
rect 12124 6128 12130 6140
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 3476 6072 3985 6100
rect 3476 6060 3482 6072
rect 3973 6069 3985 6072
rect 4019 6069 4031 6103
rect 3973 6063 4031 6069
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7193 6103 7251 6109
rect 7193 6100 7205 6103
rect 6972 6072 7205 6100
rect 6972 6060 6978 6072
rect 7193 6069 7205 6072
rect 7239 6069 7251 6103
rect 7193 6063 7251 6069
rect 7285 6103 7343 6109
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 8294 6100 8300 6112
rect 7331 6072 8300 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 9125 6103 9183 6109
rect 9125 6069 9137 6103
rect 9171 6100 9183 6103
rect 11146 6100 11152 6112
rect 9171 6072 11152 6100
rect 9171 6069 9183 6072
rect 9125 6063 9183 6069
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12802 6100 12808 6112
rect 12492 6072 12537 6100
rect 12763 6072 12808 6100
rect 12492 6060 12498 6072
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 12912 6100 12940 6140
rect 15028 6112 15056 6140
rect 14182 6100 14188 6112
rect 12912 6072 14188 6100
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 15010 6100 15016 6112
rect 14971 6072 15016 6100
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 1104 6010 16836 6032
rect 1104 5958 6246 6010
rect 6298 5958 6310 6010
rect 6362 5958 6374 6010
rect 6426 5958 6438 6010
rect 6490 5958 11510 6010
rect 11562 5958 11574 6010
rect 11626 5958 11638 6010
rect 11690 5958 11702 6010
rect 11754 5958 16836 6010
rect 1104 5936 16836 5958
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 2777 5899 2835 5905
rect 2777 5896 2789 5899
rect 1995 5868 2789 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 2777 5865 2789 5868
rect 2823 5865 2835 5899
rect 3142 5896 3148 5908
rect 3103 5868 3148 5896
rect 2777 5859 2835 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 3283 5868 4445 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 4890 5896 4896 5908
rect 4672 5868 4896 5896
rect 4672 5856 4678 5868
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 6733 5899 6791 5905
rect 6733 5896 6745 5899
rect 6696 5868 6745 5896
rect 6696 5856 6702 5868
rect 6733 5865 6745 5868
rect 6779 5865 6791 5899
rect 6733 5859 6791 5865
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8757 5899 8815 5905
rect 8757 5896 8769 5899
rect 8444 5868 8769 5896
rect 8444 5856 8450 5868
rect 8757 5865 8769 5868
rect 8803 5865 8815 5899
rect 8757 5859 8815 5865
rect 8849 5899 8907 5905
rect 8849 5865 8861 5899
rect 8895 5896 8907 5899
rect 10962 5896 10968 5908
rect 8895 5868 10968 5896
rect 8895 5865 8907 5868
rect 8849 5859 8907 5865
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 12802 5856 12808 5908
rect 12860 5896 12866 5908
rect 14001 5899 14059 5905
rect 14001 5896 14013 5899
rect 12860 5868 14013 5896
rect 12860 5856 12866 5868
rect 14001 5865 14013 5868
rect 14047 5865 14059 5899
rect 14001 5859 14059 5865
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 15286 5896 15292 5908
rect 14415 5868 15292 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 1394 5788 1400 5840
rect 1452 5828 1458 5840
rect 6825 5831 6883 5837
rect 6825 5828 6837 5831
rect 1452 5800 6837 5828
rect 1452 5788 1458 5800
rect 6825 5797 6837 5800
rect 6871 5828 6883 5831
rect 10870 5828 10876 5840
rect 6871 5800 10876 5828
rect 6871 5797 6883 5800
rect 6825 5791 6883 5797
rect 10870 5788 10876 5800
rect 10928 5828 10934 5840
rect 11146 5828 11152 5840
rect 10928 5800 11152 5828
rect 10928 5788 10934 5800
rect 11146 5788 11152 5800
rect 11204 5788 11210 5840
rect 12060 5831 12118 5837
rect 12060 5797 12072 5831
rect 12106 5828 12118 5831
rect 12526 5828 12532 5840
rect 12106 5800 12532 5828
rect 12106 5797 12118 5800
rect 12060 5791 12118 5797
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 14461 5831 14519 5837
rect 14461 5797 14473 5831
rect 14507 5828 14519 5831
rect 15194 5828 15200 5840
rect 14507 5800 15200 5828
rect 14507 5797 14519 5800
rect 14461 5791 14519 5797
rect 15194 5788 15200 5800
rect 15252 5788 15258 5840
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5760 2099 5763
rect 2958 5760 2964 5772
rect 2087 5732 2964 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 4798 5760 4804 5772
rect 4759 5732 4804 5760
rect 4798 5720 4804 5732
rect 4856 5760 4862 5772
rect 10318 5760 10324 5772
rect 4856 5732 10324 5760
rect 4856 5720 4862 5732
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10502 5760 10508 5772
rect 10463 5732 10508 5760
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 12342 5760 12348 5772
rect 11808 5732 12348 5760
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2682 5692 2688 5704
rect 2271 5664 2688 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 3326 5692 3332 5704
rect 3287 5664 3332 5692
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 5074 5692 5080 5704
rect 5035 5664 5080 5692
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 7006 5692 7012 5704
rect 6967 5664 7012 5692
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 7558 5692 7564 5704
rect 7519 5664 7564 5692
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5692 9091 5695
rect 9582 5692 9588 5704
rect 9079 5664 9588 5692
rect 9079 5661 9091 5664
rect 9033 5655 9091 5661
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 10594 5692 10600 5704
rect 10555 5664 10600 5692
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 11238 5692 11244 5704
rect 10827 5664 11244 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 11698 5652 11704 5704
rect 11756 5692 11762 5704
rect 11808 5701 11836 5732
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 15841 5763 15899 5769
rect 15841 5760 15853 5763
rect 13872 5732 15853 5760
rect 13872 5720 13878 5732
rect 15841 5729 15853 5732
rect 15887 5729 15899 5763
rect 15841 5723 15899 5729
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11756 5664 11805 5692
rect 11756 5652 11762 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 13964 5664 14565 5692
rect 13964 5652 13970 5664
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 8389 5627 8447 5633
rect 8389 5593 8401 5627
rect 8435 5624 8447 5627
rect 10686 5624 10692 5636
rect 8435 5596 10692 5624
rect 8435 5593 8447 5596
rect 8389 5587 8447 5593
rect 10686 5584 10692 5596
rect 10744 5584 10750 5636
rect 15838 5624 15844 5636
rect 13004 5596 15844 5624
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 5994 5516 6000 5568
rect 6052 5556 6058 5568
rect 6365 5559 6423 5565
rect 6365 5556 6377 5559
rect 6052 5528 6377 5556
rect 6052 5516 6058 5528
rect 6365 5525 6377 5528
rect 6411 5525 6423 5559
rect 6365 5519 6423 5525
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 10137 5559 10195 5565
rect 10137 5556 10149 5559
rect 10100 5528 10149 5556
rect 10100 5516 10106 5528
rect 10137 5525 10149 5528
rect 10183 5525 10195 5559
rect 10137 5519 10195 5525
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 13004 5556 13032 5596
rect 15838 5584 15844 5596
rect 15896 5584 15902 5636
rect 13170 5556 13176 5568
rect 10468 5528 13032 5556
rect 13131 5528 13176 5556
rect 10468 5516 10474 5528
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 16022 5556 16028 5568
rect 15983 5528 16028 5556
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 1104 5466 16836 5488
rect 1104 5414 3614 5466
rect 3666 5414 3678 5466
rect 3730 5414 3742 5466
rect 3794 5414 3806 5466
rect 3858 5414 8878 5466
rect 8930 5414 8942 5466
rect 8994 5414 9006 5466
rect 9058 5414 9070 5466
rect 9122 5414 14142 5466
rect 14194 5414 14206 5466
rect 14258 5414 14270 5466
rect 14322 5414 14334 5466
rect 14386 5414 16836 5466
rect 1104 5392 16836 5414
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 1949 5355 2007 5361
rect 1949 5352 1961 5355
rect 1728 5324 1961 5352
rect 1728 5312 1734 5324
rect 1949 5321 1961 5324
rect 1995 5321 2007 5355
rect 1949 5315 2007 5321
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 3016 5324 3157 5352
rect 3016 5312 3022 5324
rect 3145 5321 3157 5324
rect 3191 5321 3203 5355
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 3145 5315 3203 5321
rect 6840 5324 8217 5352
rect 3326 5244 3332 5296
rect 3384 5284 3390 5296
rect 3384 5256 3740 5284
rect 3384 5244 3390 5256
rect 3712 5228 3740 5256
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 2409 5219 2467 5225
rect 2409 5216 2421 5219
rect 1636 5188 2421 5216
rect 1636 5176 1642 5188
rect 2409 5185 2421 5188
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5216 2651 5219
rect 3418 5216 3424 5228
rect 2639 5188 3424 5216
rect 2639 5185 2651 5188
rect 2593 5179 2651 5185
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 3694 5216 3700 5228
rect 3655 5188 3700 5216
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 4522 5176 4528 5228
rect 4580 5216 4586 5228
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4580 5188 4813 5216
rect 4580 5176 4586 5188
rect 4801 5185 4813 5188
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5074 5216 5080 5228
rect 5031 5188 5080 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5994 5216 6000 5228
rect 5955 5188 6000 5216
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6840 5216 6868 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 12802 5352 12808 5364
rect 9456 5324 12808 5352
rect 9456 5312 9462 5324
rect 12802 5312 12808 5324
rect 12860 5352 12866 5364
rect 13078 5352 13084 5364
rect 12860 5324 13084 5352
rect 12860 5312 12866 5324
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 10045 5287 10103 5293
rect 10045 5253 10057 5287
rect 10091 5253 10103 5287
rect 10045 5247 10103 5253
rect 6227 5188 6868 5216
rect 10060 5216 10088 5247
rect 10318 5244 10324 5296
rect 10376 5284 10382 5296
rect 10505 5287 10563 5293
rect 10505 5284 10517 5287
rect 10376 5256 10517 5284
rect 10376 5244 10382 5256
rect 10505 5253 10517 5256
rect 10551 5253 10563 5287
rect 11698 5284 11704 5296
rect 10505 5247 10563 5253
rect 11164 5256 11704 5284
rect 10226 5216 10232 5228
rect 10060 5188 10232 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 2314 5148 2320 5160
rect 2275 5120 2320 5148
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 2498 5108 2504 5160
rect 2556 5148 2562 5160
rect 4709 5151 4767 5157
rect 4709 5148 4721 5151
rect 2556 5120 4721 5148
rect 2556 5108 2562 5120
rect 4709 5117 4721 5120
rect 4755 5117 4767 5151
rect 4709 5111 4767 5117
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 6196 5148 6224 5179
rect 10226 5176 10232 5188
rect 10284 5216 10290 5228
rect 10778 5216 10784 5228
rect 10284 5188 10784 5216
rect 10284 5176 10290 5188
rect 10778 5176 10784 5188
rect 10836 5216 10842 5228
rect 11057 5219 11115 5225
rect 11057 5216 11069 5219
rect 10836 5188 11069 5216
rect 10836 5176 10842 5188
rect 11057 5185 11069 5188
rect 11103 5185 11115 5219
rect 11057 5179 11115 5185
rect 5776 5120 6224 5148
rect 6825 5151 6883 5157
rect 5776 5108 5782 5120
rect 6825 5117 6837 5151
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 5442 5040 5448 5092
rect 5500 5080 5506 5092
rect 6840 5080 6868 5111
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8628 5120 8677 5148
rect 8628 5108 8634 5120
rect 8665 5117 8677 5120
rect 8711 5148 8723 5151
rect 9490 5148 9496 5160
rect 8711 5120 9496 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 9490 5108 9496 5120
rect 9548 5148 9554 5160
rect 11164 5148 11192 5256
rect 11698 5244 11704 5256
rect 11756 5244 11762 5296
rect 12526 5176 12532 5228
rect 12584 5216 12590 5228
rect 13078 5216 13084 5228
rect 12584 5188 13084 5216
rect 12584 5176 12590 5188
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 13170 5176 13176 5228
rect 13228 5216 13234 5228
rect 14277 5219 14335 5225
rect 14277 5216 14289 5219
rect 13228 5188 14289 5216
rect 13228 5176 13234 5188
rect 14277 5185 14289 5188
rect 14323 5185 14335 5219
rect 14277 5179 14335 5185
rect 9548 5120 11192 5148
rect 9548 5108 9554 5120
rect 11790 5108 11796 5160
rect 11848 5148 11854 5160
rect 11885 5151 11943 5157
rect 11885 5148 11897 5151
rect 11848 5120 11897 5148
rect 11848 5108 11854 5120
rect 11885 5117 11897 5120
rect 11931 5117 11943 5151
rect 12986 5148 12992 5160
rect 12947 5120 12992 5148
rect 11885 5111 11943 5117
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15712 5120 15853 5148
rect 15712 5108 15718 5120
rect 15841 5117 15853 5120
rect 15887 5117 15899 5151
rect 15841 5111 15899 5117
rect 5500 5052 6868 5080
rect 5500 5040 5506 5052
rect 7006 5040 7012 5092
rect 7064 5089 7070 5092
rect 7064 5083 7128 5089
rect 7064 5049 7082 5083
rect 7116 5049 7128 5083
rect 7064 5043 7128 5049
rect 8932 5083 8990 5089
rect 8932 5049 8944 5083
rect 8978 5080 8990 5083
rect 10502 5080 10508 5092
rect 8978 5052 10508 5080
rect 8978 5049 8990 5052
rect 8932 5043 8990 5049
rect 7064 5040 7070 5043
rect 10502 5040 10508 5052
rect 10560 5040 10566 5092
rect 11330 5080 11336 5092
rect 10704 5052 11336 5080
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 3513 5015 3571 5021
rect 3513 5012 3525 5015
rect 3016 4984 3525 5012
rect 3016 4972 3022 4984
rect 3513 4981 3525 4984
rect 3559 4981 3571 5015
rect 3513 4975 3571 4981
rect 3605 5015 3663 5021
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 4341 5015 4399 5021
rect 4341 5012 4353 5015
rect 3651 4984 4353 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 4341 4981 4353 4984
rect 4387 4981 4399 5015
rect 5534 5012 5540 5024
rect 5495 4984 5540 5012
rect 4341 4975 4399 4981
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 5902 5012 5908 5024
rect 5863 4984 5908 5012
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 10704 5012 10732 5052
rect 11330 5040 11336 5052
rect 11388 5040 11394 5092
rect 14185 5083 14243 5089
rect 14185 5080 14197 5083
rect 12544 5052 14197 5080
rect 10870 5012 10876 5024
rect 9824 4984 10732 5012
rect 10831 4984 10876 5012
rect 9824 4972 9830 4984
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 10962 4972 10968 5024
rect 11020 5012 11026 5024
rect 12544 5021 12572 5052
rect 14185 5049 14197 5052
rect 14231 5049 14243 5083
rect 14185 5043 14243 5049
rect 12529 5015 12587 5021
rect 11020 4984 11065 5012
rect 11020 4972 11026 4984
rect 12529 4981 12541 5015
rect 12575 4981 12587 5015
rect 12529 4975 12587 4981
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12676 4984 12909 5012
rect 12676 4972 12682 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 13722 5012 13728 5024
rect 13683 4984 13728 5012
rect 12897 4975 12955 4981
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 14090 5012 14096 5024
rect 14051 4984 14096 5012
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 16022 5012 16028 5024
rect 15983 4984 16028 5012
rect 16022 4972 16028 4984
rect 16080 4972 16086 5024
rect 1104 4922 16836 4944
rect 1104 4870 6246 4922
rect 6298 4870 6310 4922
rect 6362 4870 6374 4922
rect 6426 4870 6438 4922
rect 6490 4870 11510 4922
rect 11562 4870 11574 4922
rect 11626 4870 11638 4922
rect 11690 4870 11702 4922
rect 11754 4870 16836 4922
rect 1104 4848 16836 4870
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 3694 4808 3700 4820
rect 3559 4780 3700 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 5534 4808 5540 4820
rect 5495 4780 5540 4808
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6365 4811 6423 4817
rect 6365 4808 6377 4811
rect 5960 4780 6377 4808
rect 5960 4768 5966 4780
rect 6365 4777 6377 4780
rect 6411 4777 6423 4811
rect 6365 4771 6423 4777
rect 6733 4811 6791 4817
rect 6733 4777 6745 4811
rect 6779 4808 6791 4811
rect 7558 4808 7564 4820
rect 6779 4780 7564 4808
rect 6779 4777 6791 4780
rect 6733 4771 6791 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7708 4780 8125 4808
rect 7708 4768 7714 4780
rect 8113 4777 8125 4780
rect 8159 4777 8171 4811
rect 8113 4771 8171 4777
rect 9953 4811 10011 4817
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10870 4808 10876 4820
rect 9999 4780 10876 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 10980 4780 11621 4808
rect 9766 4740 9772 4752
rect 1412 4712 4016 4740
rect 1412 4681 1440 4712
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4641 1455 4675
rect 2130 4672 2136 4684
rect 2091 4644 2136 4672
rect 1397 4635 1455 4641
rect 2130 4632 2136 4644
rect 2188 4632 2194 4684
rect 2400 4675 2458 4681
rect 2400 4641 2412 4675
rect 2446 4672 2458 4675
rect 3418 4672 3424 4684
rect 2446 4644 3424 4672
rect 2446 4641 2458 4644
rect 2400 4635 2458 4641
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 3988 4604 4016 4712
rect 4080 4712 9772 4740
rect 4080 4681 4108 4712
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 9858 4700 9864 4752
rect 9916 4740 9922 4752
rect 10980 4740 11008 4780
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 11609 4771 11667 4777
rect 12529 4811 12587 4817
rect 12529 4777 12541 4811
rect 12575 4808 12587 4811
rect 14090 4808 14096 4820
rect 12575 4780 14096 4808
rect 12575 4777 12587 4780
rect 12529 4771 12587 4777
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 9916 4712 11008 4740
rect 9916 4700 9922 4712
rect 12802 4700 12808 4752
rect 12860 4740 12866 4752
rect 12897 4743 12955 4749
rect 12897 4740 12909 4743
rect 12860 4712 12909 4740
rect 12860 4700 12866 4712
rect 12897 4709 12909 4712
rect 12943 4709 12955 4743
rect 12897 4703 12955 4709
rect 12989 4743 13047 4749
rect 12989 4709 13001 4743
rect 13035 4740 13047 4743
rect 13262 4740 13268 4752
rect 13035 4712 13268 4740
rect 13035 4709 13047 4712
rect 12989 4703 13047 4709
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 4065 4675 4123 4681
rect 4065 4641 4077 4675
rect 4111 4641 4123 4675
rect 4065 4635 4123 4641
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4672 5687 4675
rect 6730 4672 6736 4684
rect 5675 4644 6736 4672
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 10318 4672 10324 4684
rect 6932 4644 8432 4672
rect 10279 4644 10324 4672
rect 5810 4604 5816 4616
rect 3988 4576 5580 4604
rect 5771 4576 5816 4604
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4249 4471 4307 4477
rect 4249 4468 4261 4471
rect 4212 4440 4261 4468
rect 4212 4428 4218 4440
rect 4249 4437 4261 4440
rect 4295 4437 4307 4471
rect 5166 4468 5172 4480
rect 5127 4440 5172 4468
rect 4249 4431 4307 4437
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 5552 4468 5580 4576
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 6932 4604 6960 4644
rect 6871 4576 6960 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 5626 4496 5632 4548
rect 5684 4536 5690 4548
rect 6840 4536 6868 4567
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 8202 4604 8208 4616
rect 7064 4576 7157 4604
rect 8163 4576 8208 4604
rect 7064 4564 7070 4576
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4573 8355 4607
rect 8404 4604 8432 4644
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 10744 4644 11529 4672
rect 10744 4632 10750 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 15841 4675 15899 4681
rect 15841 4641 15853 4675
rect 15887 4641 15899 4675
rect 15841 4635 15899 4641
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 8404 4576 10425 4604
rect 8297 4567 8355 4573
rect 10413 4573 10425 4576
rect 10459 4573 10471 4607
rect 10413 4567 10471 4573
rect 5684 4508 6868 4536
rect 7024 4536 7052 4564
rect 8018 4536 8024 4548
rect 7024 4508 8024 4536
rect 5684 4496 5690 4508
rect 8018 4496 8024 4508
rect 8076 4536 8082 4548
rect 8312 4536 8340 4567
rect 8076 4508 8340 4536
rect 10428 4536 10456 4567
rect 10502 4564 10508 4616
rect 10560 4604 10566 4616
rect 10597 4607 10655 4613
rect 10597 4604 10609 4607
rect 10560 4576 10609 4604
rect 10560 4564 10566 4576
rect 10597 4573 10609 4576
rect 10643 4604 10655 4607
rect 10870 4604 10876 4616
rect 10643 4576 10876 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11793 4607 11851 4613
rect 11793 4604 11805 4607
rect 11112 4576 11805 4604
rect 11112 4564 11118 4576
rect 11793 4573 11805 4576
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 13078 4564 13084 4616
rect 13136 4604 13142 4616
rect 13136 4576 13181 4604
rect 13136 4564 13142 4576
rect 12158 4536 12164 4548
rect 10428 4508 12164 4536
rect 8076 4496 8082 4508
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 15856 4536 15884 4635
rect 12544 4508 15884 4536
rect 7466 4468 7472 4480
rect 5552 4440 7472 4468
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 7742 4468 7748 4480
rect 7703 4440 7748 4468
rect 7742 4428 7748 4440
rect 7800 4428 7806 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 11149 4471 11207 4477
rect 11149 4468 11161 4471
rect 10008 4440 11161 4468
rect 10008 4428 10014 4440
rect 11149 4437 11161 4440
rect 11195 4437 11207 4471
rect 11149 4431 11207 4437
rect 11514 4428 11520 4480
rect 11572 4468 11578 4480
rect 12544 4468 12572 4508
rect 16022 4468 16028 4480
rect 11572 4440 12572 4468
rect 15983 4440 16028 4468
rect 11572 4428 11578 4440
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 1104 4378 16836 4400
rect 1104 4326 3614 4378
rect 3666 4326 3678 4378
rect 3730 4326 3742 4378
rect 3794 4326 3806 4378
rect 3858 4326 8878 4378
rect 8930 4326 8942 4378
rect 8994 4326 9006 4378
rect 9058 4326 9070 4378
rect 9122 4326 14142 4378
rect 14194 4326 14206 4378
rect 14258 4326 14270 4378
rect 14322 4326 14334 4378
rect 14386 4326 16836 4378
rect 1104 4304 16836 4326
rect 2958 4264 2964 4276
rect 2919 4236 2964 4264
rect 2958 4224 2964 4236
rect 3016 4224 3022 4276
rect 3418 4224 3424 4276
rect 3476 4264 3482 4276
rect 5074 4264 5080 4276
rect 3476 4236 5080 4264
rect 3476 4224 3482 4236
rect 3712 4196 3740 4236
rect 5074 4224 5080 4236
rect 5132 4264 5138 4276
rect 5537 4267 5595 4273
rect 5537 4264 5549 4267
rect 5132 4236 5549 4264
rect 5132 4224 5138 4236
rect 5537 4233 5549 4236
rect 5583 4233 5595 4267
rect 5537 4227 5595 4233
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 7006 4264 7012 4276
rect 6788 4236 7012 4264
rect 6788 4224 6794 4236
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7469 4267 7527 4273
rect 7469 4233 7481 4267
rect 7515 4264 7527 4267
rect 8202 4264 8208 4276
rect 7515 4236 8208 4264
rect 7515 4233 7527 4236
rect 7469 4227 7527 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 11790 4264 11796 4276
rect 8680 4236 11100 4264
rect 11703 4236 11796 4264
rect 3620 4168 3740 4196
rect 2498 4128 2504 4140
rect 1596 4100 2504 4128
rect 1596 4069 1624 4100
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 3620 4137 3648 4168
rect 7650 4156 7656 4208
rect 7708 4196 7714 4208
rect 8680 4196 8708 4236
rect 7708 4168 8708 4196
rect 7708 4156 7714 4168
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 3108 4100 3433 4128
rect 3108 4088 3114 4100
rect 3421 4097 3433 4100
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 3605 4091 3663 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8159 4100 8800 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4029 1639 4063
rect 1581 4023 1639 4029
rect 2406 4020 2412 4072
rect 2464 4060 2470 4072
rect 3329 4063 3387 4069
rect 3329 4060 3341 4063
rect 2464 4032 3341 4060
rect 2464 4020 2470 4032
rect 3329 4029 3341 4032
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 5442 4060 5448 4072
rect 4203 4032 5448 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7892 4032 7941 4060
rect 7892 4020 7898 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8628 4032 8677 4060
rect 8628 4020 8634 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 8772 4060 8800 4100
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10376 4100 10517 4128
rect 10376 4088 10382 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 8938 4069 8944 4072
rect 8921 4063 8944 4069
rect 8921 4060 8933 4063
rect 8772 4032 8933 4060
rect 8665 4023 8723 4029
rect 8921 4029 8933 4032
rect 8996 4060 9002 4072
rect 11072 4060 11100 4236
rect 11716 4137 11744 4236
rect 11790 4224 11796 4236
rect 11848 4264 11854 4276
rect 13170 4264 13176 4276
rect 11848 4236 13176 4264
rect 11848 4224 11854 4236
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 13078 4196 13084 4208
rect 13004 4168 13084 4196
rect 13004 4137 13032 4168
rect 13078 4156 13084 4168
rect 13136 4156 13142 4208
rect 13354 4156 13360 4208
rect 13412 4196 13418 4208
rect 13412 4168 15884 4196
rect 13412 4156 13418 4168
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 15010 4088 15016 4140
rect 15068 4128 15074 4140
rect 15746 4128 15752 4140
rect 15068 4100 15752 4128
rect 15068 4088 15074 4100
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 11514 4060 11520 4072
rect 8996 4032 9069 4060
rect 11072 4032 11520 4060
rect 8921 4023 8944 4029
rect 8938 4020 8944 4023
rect 8996 4020 9002 4032
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 14369 4063 14427 4069
rect 14369 4029 14381 4063
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 4424 3995 4482 4001
rect 4424 3961 4436 3995
rect 4470 3992 4482 3995
rect 5810 3992 5816 4004
rect 4470 3964 5816 3992
rect 4470 3961 4482 3964
rect 4424 3955 4482 3961
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 7190 3952 7196 4004
rect 7248 3992 7254 4004
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 7248 3964 12817 3992
rect 7248 3952 7254 3964
rect 12805 3961 12817 3964
rect 12851 3992 12863 3995
rect 13630 3992 13636 4004
rect 12851 3964 13636 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 13630 3952 13636 3964
rect 13688 3952 13694 4004
rect 14384 3992 14412 4023
rect 14918 4020 14924 4072
rect 14976 4060 14982 4072
rect 15856 4069 15884 4168
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14976 4032 15117 4060
rect 14976 4020 14982 4032
rect 15105 4029 15117 4032
rect 15151 4029 15163 4063
rect 15105 4023 15163 4029
rect 15841 4063 15899 4069
rect 15841 4029 15853 4063
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 15378 3992 15384 4004
rect 14384 3964 15384 3992
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 3142 3924 3148 3936
rect 1811 3896 3148 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 7834 3924 7840 3936
rect 7795 3896 7840 3924
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 10045 3927 10103 3933
rect 10045 3924 10057 3927
rect 8076 3896 10057 3924
rect 8076 3884 8082 3896
rect 10045 3893 10057 3896
rect 10091 3893 10103 3927
rect 10045 3887 10103 3893
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 11330 3924 11336 3936
rect 11195 3896 11336 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11609 3927 11667 3933
rect 11609 3893 11621 3927
rect 11655 3924 11667 3927
rect 12437 3927 12495 3933
rect 12437 3924 12449 3927
rect 11655 3896 12449 3924
rect 11655 3893 11667 3896
rect 11609 3887 11667 3893
rect 12437 3893 12449 3896
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 14550 3924 14556 3936
rect 12952 3896 12997 3924
rect 14511 3896 14556 3924
rect 12952 3884 12958 3896
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 15160 3896 15301 3924
rect 15160 3884 15166 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 16022 3924 16028 3936
rect 15983 3896 16028 3924
rect 15289 3887 15347 3893
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 1104 3834 16836 3856
rect 1104 3782 6246 3834
rect 6298 3782 6310 3834
rect 6362 3782 6374 3834
rect 6426 3782 6438 3834
rect 6490 3782 11510 3834
rect 11562 3782 11574 3834
rect 11626 3782 11638 3834
rect 11690 3782 11702 3834
rect 11754 3782 16836 3834
rect 1104 3760 16836 3782
rect 5166 3720 5172 3732
rect 1504 3692 5172 3720
rect 1504 3593 1532 3692
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 5868 3692 6837 3720
rect 5868 3680 5874 3692
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8757 3723 8815 3729
rect 8757 3720 8769 3723
rect 8352 3692 8769 3720
rect 8352 3680 8358 3692
rect 8757 3689 8769 3692
rect 8803 3689 8815 3723
rect 8757 3683 8815 3689
rect 5718 3661 5724 3664
rect 5712 3652 5724 3661
rect 3160 3624 5580 3652
rect 5679 3624 5724 3652
rect 3160 3593 3188 3624
rect 1489 3587 1547 3593
rect 1489 3553 1501 3587
rect 1535 3553 1547 3587
rect 1489 3547 1547 3553
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3553 2467 3587
rect 2409 3547 2467 3553
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3553 3203 3587
rect 3145 3547 3203 3553
rect 750 3476 756 3528
rect 808 3516 814 3528
rect 1673 3519 1731 3525
rect 1673 3516 1685 3519
rect 808 3488 1685 3516
rect 808 3476 814 3488
rect 1673 3485 1685 3488
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 2424 3448 2452 3547
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 4028 3556 4077 3584
rect 4028 3544 4034 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 5442 3584 5448 3596
rect 5403 3556 5448 3584
rect 4065 3547 4123 3553
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 5552 3584 5580 3624
rect 5712 3615 5724 3624
rect 5718 3612 5724 3615
rect 5776 3612 5782 3664
rect 8772 3652 8800 3683
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 10137 3723 10195 3729
rect 10137 3720 10149 3723
rect 8904 3692 10149 3720
rect 8904 3680 8910 3692
rect 10137 3689 10149 3692
rect 10183 3720 10195 3723
rect 10873 3723 10931 3729
rect 10183 3692 10456 3720
rect 10183 3689 10195 3692
rect 10137 3683 10195 3689
rect 8772 3624 10364 3652
rect 7190 3584 7196 3596
rect 5552 3556 7196 3584
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3553 8723 3587
rect 9398 3584 9404 3596
rect 8665 3547 8723 3553
rect 8772 3556 9404 3584
rect 6822 3476 6828 3528
rect 6880 3516 6886 3528
rect 8680 3516 8708 3547
rect 6880 3488 8708 3516
rect 6880 3476 6886 3488
rect 2424 3420 5488 3448
rect 2593 3383 2651 3389
rect 2593 3349 2605 3383
rect 2639 3380 2651 3383
rect 2958 3380 2964 3392
rect 2639 3352 2964 3380
rect 2639 3349 2651 3352
rect 2593 3343 2651 3349
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 3326 3380 3332 3392
rect 3287 3352 3332 3380
rect 3326 3340 3332 3352
rect 3384 3340 3390 3392
rect 3418 3340 3424 3392
rect 3476 3380 3482 3392
rect 4249 3383 4307 3389
rect 4249 3380 4261 3383
rect 3476 3352 4261 3380
rect 3476 3340 3482 3352
rect 4249 3349 4261 3352
rect 4295 3349 4307 3383
rect 5460 3380 5488 3420
rect 7374 3408 7380 3460
rect 7432 3448 7438 3460
rect 8772 3448 8800 3556
rect 9398 3544 9404 3556
rect 9456 3584 9462 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9456 3556 10057 3584
rect 9456 3544 9462 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 8938 3516 8944 3528
rect 8899 3488 8944 3516
rect 8938 3476 8944 3488
rect 8996 3516 9002 3528
rect 9582 3516 9588 3528
rect 8996 3488 9588 3516
rect 8996 3476 9002 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 7432 3420 8800 3448
rect 9600 3448 9628 3476
rect 10244 3448 10272 3479
rect 9600 3420 10272 3448
rect 10336 3448 10364 3624
rect 10428 3584 10456 3692
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 10962 3720 10968 3732
rect 10919 3692 10968 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 11204 3692 11345 3720
rect 11204 3680 11210 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 11333 3683 11391 3689
rect 11241 3655 11299 3661
rect 11241 3621 11253 3655
rect 11287 3652 11299 3655
rect 12066 3652 12072 3664
rect 11287 3624 12072 3652
rect 11287 3621 11299 3624
rect 11241 3615 11299 3621
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 13262 3584 13268 3596
rect 10428 3556 13268 3584
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 14461 3587 14519 3593
rect 14461 3553 14473 3587
rect 14507 3584 14519 3587
rect 15562 3584 15568 3596
rect 14507 3556 15568 3584
rect 14507 3553 14519 3556
rect 14461 3547 14519 3553
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 15841 3587 15899 3593
rect 15841 3553 15853 3587
rect 15887 3584 15899 3587
rect 16298 3584 16304 3596
rect 15887 3556 16304 3584
rect 15887 3553 15899 3556
rect 15841 3547 15899 3553
rect 16298 3544 16304 3556
rect 16356 3544 16362 3596
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 11517 3519 11575 3525
rect 11517 3516 11529 3519
rect 10928 3488 11529 3516
rect 10928 3476 10934 3488
rect 11517 3485 11529 3488
rect 11563 3516 11575 3519
rect 11790 3516 11796 3528
rect 11563 3488 11796 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 12986 3448 12992 3460
rect 10336 3420 12992 3448
rect 7432 3408 7438 3420
rect 12986 3408 12992 3420
rect 13044 3408 13050 3460
rect 7098 3380 7104 3392
rect 5460 3352 7104 3380
rect 4249 3343 4307 3349
rect 7098 3340 7104 3352
rect 7156 3380 7162 3392
rect 7834 3380 7840 3392
rect 7156 3352 7840 3380
rect 7156 3340 7162 3352
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 8294 3380 8300 3392
rect 8255 3352 8300 3380
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 9677 3383 9735 3389
rect 9677 3380 9689 3383
rect 8444 3352 9689 3380
rect 8444 3340 8450 3352
rect 9677 3349 9689 3352
rect 9723 3349 9735 3383
rect 14642 3380 14648 3392
rect 14603 3352 14648 3380
rect 9677 3343 9735 3349
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 16022 3380 16028 3392
rect 15983 3352 16028 3380
rect 16022 3340 16028 3352
rect 16080 3340 16086 3392
rect 1104 3290 16836 3312
rect 1104 3238 3614 3290
rect 3666 3238 3678 3290
rect 3730 3238 3742 3290
rect 3794 3238 3806 3290
rect 3858 3238 8878 3290
rect 8930 3238 8942 3290
rect 8994 3238 9006 3290
rect 9058 3238 9070 3290
rect 9122 3238 14142 3290
rect 14194 3238 14206 3290
rect 14258 3238 14270 3290
rect 14322 3238 14334 3290
rect 14386 3238 16836 3290
rect 1104 3216 16836 3238
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3176 2007 3179
rect 2774 3176 2780 3188
rect 1995 3148 2780 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 6822 3176 6828 3188
rect 5644 3148 6828 3176
rect 5644 3108 5672 3148
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 8570 3176 8576 3188
rect 8220 3148 8576 3176
rect 1780 3080 5672 3108
rect 1780 2981 1808 3080
rect 5718 3068 5724 3120
rect 5776 3108 5782 3120
rect 5776 3080 7604 3108
rect 5776 3068 5782 3080
rect 3234 3000 3240 3052
rect 3292 3040 3298 3052
rect 6086 3040 6092 3052
rect 3292 3012 4752 3040
rect 3292 3000 3298 3012
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2941 1823 2975
rect 1765 2935 1823 2941
rect 2501 2975 2559 2981
rect 2501 2941 2513 2975
rect 2547 2941 2559 2975
rect 2501 2935 2559 2941
rect 2516 2904 2544 2935
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 4724 2981 4752 3012
rect 5828 3012 6092 3040
rect 5828 2981 5856 3012
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 7576 3049 7604 3080
rect 8220 3049 8248 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 9582 3176 9588 3188
rect 9543 3148 9588 3176
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10652 3148 10977 3176
rect 10652 3136 10658 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 10965 3139 11023 3145
rect 13722 3108 13728 3120
rect 11440 3080 13728 3108
rect 11440 3049 11468 3080
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 11425 3043 11483 3049
rect 11425 3009 11437 3043
rect 11471 3009 11483 3043
rect 11425 3003 11483 3009
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 3789 2975 3847 2981
rect 3789 2972 3801 2975
rect 3568 2944 3801 2972
rect 3568 2932 3574 2944
rect 3789 2941 3801 2944
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2941 5871 2975
rect 5813 2935 5871 2941
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2972 7435 2975
rect 7742 2972 7748 2984
rect 7423 2944 7748 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 10042 2972 10048 2984
rect 10003 2944 10048 2972
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 11330 2972 11336 2984
rect 11291 2944 11336 2972
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 2516 2876 3924 2904
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2836 2743 2839
rect 3050 2836 3056 2848
rect 2731 2808 3056 2836
rect 2731 2805 2743 2808
rect 2685 2799 2743 2805
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 3896 2836 3924 2876
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 4065 2907 4123 2913
rect 4065 2904 4077 2907
rect 4028 2876 4077 2904
rect 4028 2864 4034 2876
rect 4065 2873 4077 2876
rect 4111 2873 4123 2907
rect 4065 2867 4123 2873
rect 4985 2907 5043 2913
rect 4985 2873 4997 2907
rect 5031 2904 5043 2907
rect 5258 2904 5264 2916
rect 5031 2876 5264 2904
rect 5031 2873 5043 2876
rect 4985 2867 5043 2873
rect 5258 2864 5264 2876
rect 5316 2864 5322 2916
rect 6089 2907 6147 2913
rect 6089 2873 6101 2907
rect 6135 2904 6147 2907
rect 6730 2904 6736 2916
rect 6135 2876 6736 2904
rect 6135 2873 6147 2876
rect 6089 2867 6147 2873
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 8472 2907 8530 2913
rect 8472 2873 8484 2907
rect 8518 2904 8530 2907
rect 8518 2876 9720 2904
rect 8518 2873 8530 2876
rect 8472 2867 8530 2873
rect 7374 2836 7380 2848
rect 3896 2808 7380 2836
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 9692 2836 9720 2876
rect 9766 2864 9772 2916
rect 9824 2904 9830 2916
rect 10321 2907 10379 2913
rect 10321 2904 10333 2907
rect 9824 2876 10333 2904
rect 9824 2864 9830 2876
rect 10321 2873 10333 2876
rect 10367 2873 10379 2907
rect 10321 2867 10379 2873
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 11532 2904 11560 3003
rect 12894 3000 12900 3052
rect 12952 3040 12958 3052
rect 12952 3012 15884 3040
rect 12952 3000 12958 3012
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 12492 2944 12817 2972
rect 12492 2932 12498 2944
rect 12805 2941 12817 2944
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 15856 2981 15884 3012
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13044 2944 14197 2972
rect 13044 2932 13050 2944
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 14921 2975 14979 2981
rect 14921 2941 14933 2975
rect 14967 2941 14979 2975
rect 14921 2935 14979 2941
rect 15841 2975 15899 2981
rect 15841 2941 15853 2975
rect 15887 2941 15899 2975
rect 15841 2935 15899 2941
rect 10836 2876 11560 2904
rect 10836 2864 10842 2876
rect 12710 2864 12716 2916
rect 12768 2904 12774 2916
rect 13081 2907 13139 2913
rect 13081 2904 13093 2907
rect 12768 2876 13093 2904
rect 12768 2864 12774 2876
rect 13081 2873 13093 2876
rect 13127 2873 13139 2907
rect 13081 2867 13139 2873
rect 13262 2864 13268 2916
rect 13320 2904 13326 2916
rect 14936 2904 14964 2935
rect 13320 2876 14964 2904
rect 13320 2864 13326 2876
rect 13998 2836 14004 2848
rect 7524 2808 7569 2836
rect 9692 2808 14004 2836
rect 7524 2796 7530 2808
rect 13998 2796 14004 2808
rect 14056 2796 14062 2848
rect 14369 2839 14427 2845
rect 14369 2805 14381 2839
rect 14415 2836 14427 2839
rect 14918 2836 14924 2848
rect 14415 2808 14924 2836
rect 14415 2805 14427 2808
rect 14369 2799 14427 2805
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 15102 2836 15108 2848
rect 15063 2808 15108 2836
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 16022 2836 16028 2848
rect 15983 2808 16028 2836
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 1104 2746 16836 2768
rect 1104 2694 6246 2746
rect 6298 2694 6310 2746
rect 6362 2694 6374 2746
rect 6426 2694 6438 2746
rect 6490 2694 11510 2746
rect 11562 2694 11574 2746
rect 11626 2694 11638 2746
rect 11690 2694 11702 2746
rect 11754 2694 16836 2746
rect 1104 2672 16836 2694
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 7653 2635 7711 2641
rect 7653 2632 7665 2635
rect 7524 2604 7665 2632
rect 7524 2592 7530 2604
rect 7653 2601 7665 2604
rect 7699 2601 7711 2635
rect 7653 2595 7711 2601
rect 8113 2635 8171 2641
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 8294 2632 8300 2644
rect 8159 2604 8300 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8021 2567 8079 2573
rect 8021 2533 8033 2567
rect 8067 2564 8079 2567
rect 8386 2564 8392 2576
rect 8067 2536 8392 2564
rect 8067 2533 8079 2536
rect 8021 2527 8079 2533
rect 8386 2524 8392 2536
rect 8444 2524 8450 2576
rect 8487 2536 14688 2564
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2406 2496 2412 2508
rect 1995 2468 2412 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2406 2456 2412 2468
rect 2464 2456 2470 2508
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2496 2743 2499
rect 4798 2496 4804 2508
rect 2731 2468 4804 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 7926 2456 7932 2508
rect 7984 2496 7990 2508
rect 8487 2496 8515 2536
rect 7984 2468 8515 2496
rect 11333 2499 11391 2505
rect 7984 2456 7990 2468
rect 11333 2465 11345 2499
rect 11379 2496 11391 2499
rect 11974 2496 11980 2508
rect 11379 2468 11980 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 14660 2505 14688 2536
rect 14645 2499 14703 2505
rect 14645 2465 14657 2499
rect 14691 2465 14703 2499
rect 15838 2496 15844 2508
rect 15799 2468 15844 2496
rect 14645 2459 14703 2465
rect 15838 2456 15844 2468
rect 15896 2456 15902 2508
rect 8018 2388 8024 2440
rect 8076 2428 8082 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 8076 2400 8217 2428
rect 8076 2388 8082 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11296 2400 11529 2428
rect 11296 2388 11302 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 2130 2292 2136 2304
rect 2091 2264 2136 2292
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 2866 2292 2872 2304
rect 2827 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 9214 2292 9220 2304
rect 8260 2264 9220 2292
rect 8260 2252 8266 2264
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 14826 2292 14832 2304
rect 14787 2264 14832 2292
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 16022 2292 16028 2304
rect 15983 2264 16028 2292
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 1104 2202 16836 2224
rect 1104 2150 3614 2202
rect 3666 2150 3678 2202
rect 3730 2150 3742 2202
rect 3794 2150 3806 2202
rect 3858 2150 8878 2202
rect 8930 2150 8942 2202
rect 8994 2150 9006 2202
rect 9058 2150 9070 2202
rect 9122 2150 14142 2202
rect 14194 2150 14206 2202
rect 14258 2150 14270 2202
rect 14322 2150 14334 2202
rect 14386 2150 16836 2202
rect 1104 2128 16836 2150
<< via1 >>
rect 3884 15240 3936 15292
rect 6552 15240 6604 15292
rect 11888 15172 11940 15224
rect 14924 15172 14976 15224
rect 3516 14764 3568 14816
rect 10324 14764 10376 14816
rect 6246 14662 6298 14714
rect 6310 14662 6362 14714
rect 6374 14662 6426 14714
rect 6438 14662 6490 14714
rect 11510 14662 11562 14714
rect 11574 14662 11626 14714
rect 11638 14662 11690 14714
rect 11702 14662 11754 14714
rect 3614 14118 3666 14170
rect 3678 14118 3730 14170
rect 3742 14118 3794 14170
rect 3806 14118 3858 14170
rect 8878 14118 8930 14170
rect 8942 14118 8994 14170
rect 9006 14118 9058 14170
rect 9070 14118 9122 14170
rect 14142 14118 14194 14170
rect 14206 14118 14258 14170
rect 14270 14118 14322 14170
rect 14334 14118 14386 14170
rect 6246 13574 6298 13626
rect 6310 13574 6362 13626
rect 6374 13574 6426 13626
rect 6438 13574 6490 13626
rect 11510 13574 11562 13626
rect 11574 13574 11626 13626
rect 11638 13574 11690 13626
rect 11702 13574 11754 13626
rect 3614 13030 3666 13082
rect 3678 13030 3730 13082
rect 3742 13030 3794 13082
rect 3806 13030 3858 13082
rect 8878 13030 8930 13082
rect 8942 13030 8994 13082
rect 9006 13030 9058 13082
rect 9070 13030 9122 13082
rect 14142 13030 14194 13082
rect 14206 13030 14258 13082
rect 14270 13030 14322 13082
rect 14334 13030 14386 13082
rect 3516 12656 3568 12708
rect 7656 12656 7708 12708
rect 4068 12588 4120 12640
rect 10784 12588 10836 12640
rect 6246 12486 6298 12538
rect 6310 12486 6362 12538
rect 6374 12486 6426 12538
rect 6438 12486 6490 12538
rect 11510 12486 11562 12538
rect 11574 12486 11626 12538
rect 11638 12486 11690 12538
rect 11702 12486 11754 12538
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 13820 12384 13872 12436
rect 2872 12316 2924 12368
rect 9220 12316 9272 12368
rect 1952 12248 2004 12300
rect 3976 12248 4028 12300
rect 6644 12291 6696 12300
rect 6644 12257 6653 12291
rect 6653 12257 6687 12291
rect 6687 12257 6696 12291
rect 6644 12248 6696 12257
rect 7380 12248 7432 12300
rect 7656 12248 7708 12300
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 3332 12180 3384 12232
rect 4252 12180 4304 12232
rect 5540 12180 5592 12232
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 8208 12180 8260 12232
rect 15660 12180 15712 12232
rect 7840 12112 7892 12164
rect 3240 12044 3292 12096
rect 6092 12044 6144 12096
rect 7472 12087 7524 12096
rect 7472 12053 7481 12087
rect 7481 12053 7515 12087
rect 7515 12053 7524 12087
rect 7472 12044 7524 12053
rect 7656 12044 7708 12096
rect 9312 12044 9364 12096
rect 14832 12044 14884 12096
rect 16212 12044 16264 12096
rect 3614 11942 3666 11994
rect 3678 11942 3730 11994
rect 3742 11942 3794 11994
rect 3806 11942 3858 11994
rect 8878 11942 8930 11994
rect 8942 11942 8994 11994
rect 9006 11942 9058 11994
rect 9070 11942 9122 11994
rect 14142 11942 14194 11994
rect 14206 11942 14258 11994
rect 14270 11942 14322 11994
rect 14334 11942 14386 11994
rect 1952 11883 2004 11892
rect 1952 11849 1961 11883
rect 1961 11849 1995 11883
rect 1995 11849 2004 11883
rect 1952 11840 2004 11849
rect 2964 11840 3016 11892
rect 3516 11840 3568 11892
rect 3976 11883 4028 11892
rect 3976 11849 3985 11883
rect 3985 11849 4019 11883
rect 4019 11849 4028 11883
rect 3976 11840 4028 11849
rect 6644 11840 6696 11892
rect 3424 11772 3476 11824
rect 6000 11772 6052 11824
rect 7840 11772 7892 11824
rect 9036 11772 9088 11824
rect 12164 11772 12216 11824
rect 14556 11772 14608 11824
rect 2228 11704 2280 11756
rect 3332 11704 3384 11756
rect 7656 11704 7708 11756
rect 8024 11747 8076 11756
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 8852 11704 8904 11756
rect 11336 11704 11388 11756
rect 13452 11704 13504 11756
rect 14280 11704 14332 11756
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 2320 11679 2372 11688
rect 2320 11645 2329 11679
rect 2329 11645 2363 11679
rect 2363 11645 2372 11679
rect 2320 11636 2372 11645
rect 4988 11636 5040 11688
rect 5816 11636 5868 11688
rect 7840 11636 7892 11688
rect 9404 11636 9456 11688
rect 15844 11636 15896 11688
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 2780 11500 2832 11552
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 4436 11543 4488 11552
rect 4436 11509 4445 11543
rect 4445 11509 4479 11543
rect 4479 11509 4488 11543
rect 4436 11500 4488 11509
rect 4896 11500 4948 11552
rect 15660 11568 15712 11620
rect 7564 11500 7616 11552
rect 9312 11500 9364 11552
rect 12440 11543 12492 11552
rect 12440 11509 12449 11543
rect 12449 11509 12483 11543
rect 12483 11509 12492 11543
rect 12808 11543 12860 11552
rect 12440 11500 12492 11509
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 14924 11543 14976 11552
rect 12900 11500 12952 11509
rect 14924 11509 14933 11543
rect 14933 11509 14967 11543
rect 14967 11509 14976 11543
rect 14924 11500 14976 11509
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 6246 11398 6298 11450
rect 6310 11398 6362 11450
rect 6374 11398 6426 11450
rect 6438 11398 6490 11450
rect 11510 11398 11562 11450
rect 11574 11398 11626 11450
rect 11638 11398 11690 11450
rect 11702 11398 11754 11450
rect 3332 11339 3384 11348
rect 3332 11305 3341 11339
rect 3341 11305 3375 11339
rect 3375 11305 3384 11339
rect 3332 11296 3384 11305
rect 4344 11296 4396 11348
rect 4896 11339 4948 11348
rect 4896 11305 4905 11339
rect 4905 11305 4939 11339
rect 4939 11305 4948 11339
rect 4896 11296 4948 11305
rect 8760 11296 8812 11348
rect 9036 11296 9088 11348
rect 14280 11339 14332 11348
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 15384 11339 15436 11348
rect 15384 11305 15393 11339
rect 15393 11305 15427 11339
rect 15427 11305 15436 11339
rect 15384 11296 15436 11305
rect 15752 11339 15804 11348
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 15752 11296 15804 11305
rect 4988 11271 5040 11280
rect 4988 11237 4997 11271
rect 4997 11237 5031 11271
rect 5031 11237 5040 11271
rect 4988 11228 5040 11237
rect 2228 11203 2280 11212
rect 2228 11169 2262 11203
rect 2262 11169 2280 11203
rect 2228 11160 2280 11169
rect 6736 11228 6788 11280
rect 8852 11228 8904 11280
rect 9220 11228 9272 11280
rect 6644 11160 6696 11212
rect 8300 11160 8352 11212
rect 11888 11160 11940 11212
rect 12992 11160 13044 11212
rect 13544 11160 13596 11212
rect 14004 11228 14056 11280
rect 16304 11160 16356 11212
rect 1952 11135 2004 11144
rect 1952 11101 1961 11135
rect 1961 11101 1995 11135
rect 1995 11101 2004 11135
rect 1952 11092 2004 11101
rect 5264 11092 5316 11144
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 4068 11024 4120 11076
rect 5816 11024 5868 11076
rect 6828 11024 6880 11076
rect 2596 10956 2648 11008
rect 3148 10956 3200 11008
rect 13268 10956 13320 11008
rect 3614 10854 3666 10906
rect 3678 10854 3730 10906
rect 3742 10854 3794 10906
rect 3806 10854 3858 10906
rect 8878 10854 8930 10906
rect 8942 10854 8994 10906
rect 9006 10854 9058 10906
rect 9070 10854 9122 10906
rect 14142 10854 14194 10906
rect 14206 10854 14258 10906
rect 14270 10854 14322 10906
rect 14334 10854 14386 10906
rect 2136 10752 2188 10804
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 4436 10752 4488 10804
rect 4804 10752 4856 10804
rect 11888 10752 11940 10804
rect 12900 10795 12952 10804
rect 12900 10761 12909 10795
rect 12909 10761 12943 10795
rect 12943 10761 12952 10795
rect 12900 10752 12952 10761
rect 12992 10752 13044 10804
rect 15568 10795 15620 10804
rect 4068 10684 4120 10736
rect 8208 10684 8260 10736
rect 2228 10616 2280 10668
rect 1952 10548 2004 10600
rect 4804 10616 4856 10668
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 6644 10616 6696 10668
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 2964 10480 3016 10532
rect 3332 10480 3384 10532
rect 4712 10480 4764 10532
rect 6000 10548 6052 10600
rect 7380 10548 7432 10600
rect 7012 10480 7064 10532
rect 8760 10548 8812 10600
rect 9220 10548 9272 10600
rect 9772 10548 9824 10600
rect 14004 10684 14056 10736
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 15568 10761 15577 10795
rect 15577 10761 15611 10795
rect 15611 10761 15620 10795
rect 15568 10752 15620 10761
rect 13544 10616 13596 10625
rect 11888 10548 11940 10600
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 2136 10412 2188 10421
rect 5264 10412 5316 10464
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 8116 10412 8168 10464
rect 8760 10412 8812 10464
rect 9312 10480 9364 10532
rect 10600 10480 10652 10532
rect 11336 10480 11388 10532
rect 13820 10480 13872 10532
rect 15200 10480 15252 10532
rect 9772 10412 9824 10464
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 12716 10412 12768 10464
rect 13268 10455 13320 10464
rect 13268 10421 13277 10455
rect 13277 10421 13311 10455
rect 13311 10421 13320 10455
rect 13268 10412 13320 10421
rect 14556 10412 14608 10464
rect 6246 10310 6298 10362
rect 6310 10310 6362 10362
rect 6374 10310 6426 10362
rect 6438 10310 6490 10362
rect 11510 10310 11562 10362
rect 11574 10310 11626 10362
rect 11638 10310 11690 10362
rect 11702 10310 11754 10362
rect 2412 10208 2464 10260
rect 2688 10251 2740 10260
rect 2688 10217 2697 10251
rect 2697 10217 2731 10251
rect 2731 10217 2740 10251
rect 2688 10208 2740 10217
rect 2872 10208 2924 10260
rect 3148 10208 3200 10260
rect 4620 10208 4672 10260
rect 5080 10208 5132 10260
rect 5264 10208 5316 10260
rect 2688 10072 2740 10124
rect 2964 10072 3016 10124
rect 4252 10140 4304 10192
rect 7380 10140 7432 10192
rect 10048 10183 10100 10192
rect 2688 9936 2740 9988
rect 4068 9868 4120 9920
rect 7104 9936 7156 9988
rect 4804 9868 4856 9920
rect 6920 9868 6972 9920
rect 8668 10072 8720 10124
rect 8760 10115 8812 10124
rect 8760 10081 8769 10115
rect 8769 10081 8803 10115
rect 8803 10081 8812 10115
rect 10048 10149 10082 10183
rect 10082 10149 10100 10183
rect 10048 10140 10100 10149
rect 12440 10208 12492 10260
rect 12624 10208 12676 10260
rect 13084 10208 13136 10260
rect 13360 10208 13412 10260
rect 13728 10140 13780 10192
rect 8760 10072 8812 10081
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 8116 10004 8168 10056
rect 8484 10004 8536 10056
rect 9220 10004 9272 10056
rect 8760 9868 8812 9920
rect 9312 9868 9364 9920
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 14004 10072 14056 10124
rect 12716 10004 12768 10056
rect 13360 10047 13412 10056
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 15108 10140 15160 10192
rect 15292 10140 15344 10192
rect 15384 10072 15436 10124
rect 15568 10004 15620 10056
rect 11244 9868 11296 9920
rect 11980 9868 12032 9920
rect 13636 9936 13688 9988
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 16028 9936 16080 9988
rect 13912 9868 13964 9920
rect 15752 9868 15804 9920
rect 3614 9766 3666 9818
rect 3678 9766 3730 9818
rect 3742 9766 3794 9818
rect 3806 9766 3858 9818
rect 8878 9766 8930 9818
rect 8942 9766 8994 9818
rect 9006 9766 9058 9818
rect 9070 9766 9122 9818
rect 14142 9766 14194 9818
rect 14206 9766 14258 9818
rect 14270 9766 14322 9818
rect 14334 9766 14386 9818
rect 2044 9707 2096 9716
rect 2044 9673 2053 9707
rect 2053 9673 2087 9707
rect 2087 9673 2096 9707
rect 2044 9664 2096 9673
rect 2964 9664 3016 9716
rect 4068 9664 4120 9716
rect 4712 9707 4764 9716
rect 4712 9673 4721 9707
rect 4721 9673 4755 9707
rect 4755 9673 4764 9707
rect 4712 9664 4764 9673
rect 4804 9664 4856 9716
rect 6736 9664 6788 9716
rect 7104 9664 7156 9716
rect 2320 9596 2372 9648
rect 5540 9639 5592 9648
rect 2688 9571 2740 9580
rect 2688 9537 2697 9571
rect 2697 9537 2731 9571
rect 2731 9537 2740 9571
rect 5540 9605 5549 9639
rect 5549 9605 5583 9639
rect 5583 9605 5592 9639
rect 5540 9596 5592 9605
rect 6828 9596 6880 9648
rect 7840 9664 7892 9716
rect 8668 9639 8720 9648
rect 2688 9528 2740 9537
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 5356 9503 5408 9512
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 8668 9605 8677 9639
rect 8677 9605 8711 9639
rect 8711 9605 8720 9639
rect 8668 9596 8720 9605
rect 10324 9596 10376 9648
rect 14648 9664 14700 9716
rect 16396 9664 16448 9716
rect 15016 9596 15068 9648
rect 15384 9639 15436 9648
rect 15384 9605 15393 9639
rect 15393 9605 15427 9639
rect 15427 9605 15436 9639
rect 15384 9596 15436 9605
rect 9220 9571 9272 9580
rect 6736 9460 6788 9512
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 10048 9528 10100 9580
rect 10508 9528 10560 9580
rect 10876 9528 10928 9580
rect 3516 9392 3568 9444
rect 4160 9392 4212 9444
rect 5632 9392 5684 9444
rect 6920 9392 6972 9444
rect 7104 9503 7156 9512
rect 7104 9469 7138 9503
rect 7138 9469 7156 9503
rect 7104 9460 7156 9469
rect 7380 9460 7432 9512
rect 11796 9460 11848 9512
rect 14464 9528 14516 9580
rect 14832 9528 14884 9580
rect 15200 9528 15252 9580
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 10692 9435 10744 9444
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2412 9324 2464 9333
rect 2872 9324 2924 9376
rect 5724 9324 5776 9376
rect 7288 9324 7340 9376
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 9128 9367 9180 9376
rect 9128 9333 9137 9367
rect 9137 9333 9171 9367
rect 9171 9333 9180 9367
rect 10232 9367 10284 9376
rect 9128 9324 9180 9333
rect 10232 9333 10241 9367
rect 10241 9333 10275 9367
rect 10275 9333 10284 9367
rect 10232 9324 10284 9333
rect 10692 9401 10701 9435
rect 10701 9401 10735 9435
rect 10735 9401 10744 9435
rect 10692 9392 10744 9401
rect 13820 9460 13872 9512
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 10968 9324 11020 9376
rect 12707 9435 12759 9444
rect 12707 9401 12739 9435
rect 12739 9401 12759 9435
rect 12707 9392 12759 9401
rect 13636 9392 13688 9444
rect 15384 9392 15436 9444
rect 12900 9324 12952 9376
rect 13728 9324 13780 9376
rect 14832 9367 14884 9376
rect 14832 9333 14841 9367
rect 14841 9333 14875 9367
rect 14875 9333 14884 9367
rect 14832 9324 14884 9333
rect 15936 9324 15988 9376
rect 6246 9222 6298 9274
rect 6310 9222 6362 9274
rect 6374 9222 6426 9274
rect 6438 9222 6490 9274
rect 11510 9222 11562 9274
rect 11574 9222 11626 9274
rect 11638 9222 11690 9274
rect 11702 9222 11754 9274
rect 2136 9120 2188 9172
rect 2320 8984 2372 9036
rect 4252 9120 4304 9172
rect 4344 9120 4396 9172
rect 7288 9163 7340 9172
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 7656 9120 7708 9172
rect 8208 9120 8260 9172
rect 12440 9120 12492 9172
rect 3148 9052 3200 9104
rect 7104 9052 7156 9104
rect 3332 8984 3384 9036
rect 4160 8984 4212 9036
rect 4252 8984 4304 9036
rect 4896 8984 4948 9036
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 3516 8916 3568 8968
rect 3976 8916 4028 8968
rect 4804 8916 4856 8968
rect 5172 8984 5224 9036
rect 5724 8984 5776 9036
rect 3148 8848 3200 8900
rect 3332 8848 3384 8900
rect 5080 8848 5132 8900
rect 6828 8916 6880 8968
rect 7748 9052 7800 9104
rect 10416 9052 10468 9104
rect 12808 9120 12860 9172
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 14924 9120 14976 9172
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 15752 9120 15804 9129
rect 15200 9052 15252 9104
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 9772 8984 9824 9036
rect 10968 8984 11020 9036
rect 11244 8984 11296 9036
rect 13360 8984 13412 9036
rect 14464 9027 14516 9036
rect 14464 8993 14473 9027
rect 14473 8993 14507 9027
rect 14507 8993 14516 9027
rect 14464 8984 14516 8993
rect 8300 8916 8352 8968
rect 9220 8916 9272 8968
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 12440 8916 12492 8968
rect 13176 8916 13228 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 2320 8780 2372 8832
rect 2504 8780 2556 8832
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 4252 8823 4304 8832
rect 4252 8789 4261 8823
rect 4261 8789 4295 8823
rect 4295 8789 4304 8823
rect 4252 8780 4304 8789
rect 5264 8780 5316 8832
rect 9956 8823 10008 8832
rect 9956 8789 9965 8823
rect 9965 8789 9999 8823
rect 9999 8789 10008 8823
rect 9956 8780 10008 8789
rect 12532 8848 12584 8900
rect 13820 8848 13872 8900
rect 13268 8780 13320 8832
rect 13452 8780 13504 8832
rect 14004 8848 14056 8900
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 3614 8678 3666 8730
rect 3678 8678 3730 8730
rect 3742 8678 3794 8730
rect 3806 8678 3858 8730
rect 8878 8678 8930 8730
rect 8942 8678 8994 8730
rect 9006 8678 9058 8730
rect 9070 8678 9122 8730
rect 14142 8678 14194 8730
rect 14206 8678 14258 8730
rect 14270 8678 14322 8730
rect 14334 8678 14386 8730
rect 3332 8576 3384 8628
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 7104 8576 7156 8628
rect 13360 8576 13412 8628
rect 3884 8508 3936 8560
rect 4988 8508 5040 8560
rect 7932 8508 7984 8560
rect 9864 8551 9916 8560
rect 9864 8517 9873 8551
rect 9873 8517 9907 8551
rect 9907 8517 9916 8551
rect 9864 8508 9916 8517
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 5172 8440 5224 8492
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 12900 8508 12952 8560
rect 11152 8440 11204 8492
rect 11336 8440 11388 8492
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 13268 8440 13320 8449
rect 15108 8508 15160 8560
rect 5264 8372 5316 8424
rect 7196 8372 7248 8424
rect 9772 8372 9824 8424
rect 10324 8372 10376 8424
rect 10784 8372 10836 8424
rect 13360 8372 13412 8424
rect 13820 8372 13872 8424
rect 15844 8415 15896 8424
rect 3884 8304 3936 8356
rect 1584 8279 1636 8288
rect 1584 8245 1593 8279
rect 1593 8245 1627 8279
rect 1627 8245 1636 8279
rect 1584 8236 1636 8245
rect 3976 8236 4028 8288
rect 6920 8304 6972 8356
rect 8116 8304 8168 8356
rect 9036 8304 9088 8356
rect 9864 8304 9916 8356
rect 7104 8236 7156 8288
rect 9588 8236 9640 8288
rect 11520 8347 11572 8356
rect 11520 8313 11529 8347
rect 11529 8313 11563 8347
rect 11563 8313 11572 8347
rect 11520 8304 11572 8313
rect 13084 8304 13136 8356
rect 13728 8304 13780 8356
rect 15844 8381 15853 8415
rect 15853 8381 15887 8415
rect 15887 8381 15896 8415
rect 15844 8372 15896 8381
rect 16120 8304 16172 8356
rect 10416 8236 10468 8288
rect 12624 8236 12676 8288
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 15844 8236 15896 8288
rect 6246 8134 6298 8186
rect 6310 8134 6362 8186
rect 6374 8134 6426 8186
rect 6438 8134 6490 8186
rect 11510 8134 11562 8186
rect 11574 8134 11626 8186
rect 11638 8134 11690 8186
rect 11702 8134 11754 8186
rect 3148 8075 3200 8084
rect 3148 8041 3157 8075
rect 3157 8041 3191 8075
rect 3191 8041 3200 8075
rect 3148 8032 3200 8041
rect 7288 8032 7340 8084
rect 7472 8032 7524 8084
rect 7656 8032 7708 8084
rect 8760 8032 8812 8084
rect 9956 8032 10008 8084
rect 10232 8075 10284 8084
rect 10232 8041 10241 8075
rect 10241 8041 10275 8075
rect 10275 8041 10284 8075
rect 10232 8032 10284 8041
rect 12440 8032 12492 8084
rect 12808 8032 12860 8084
rect 3148 7896 3200 7948
rect 4068 7896 4120 7948
rect 4896 7939 4948 7948
rect 4896 7905 4905 7939
rect 4905 7905 4939 7939
rect 4939 7905 4948 7939
rect 4896 7896 4948 7905
rect 11060 7964 11112 8016
rect 11520 7964 11572 8016
rect 11704 7964 11756 8016
rect 12624 7964 12676 8016
rect 14096 8032 14148 8084
rect 14464 8032 14516 8084
rect 16120 8032 16172 8084
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 7104 7939 7156 7948
rect 7104 7905 7113 7939
rect 7113 7905 7147 7939
rect 7147 7905 7156 7939
rect 7104 7896 7156 7905
rect 10140 7896 10192 7948
rect 11612 7896 11664 7948
rect 14740 7964 14792 8016
rect 14832 7964 14884 8016
rect 15476 7964 15528 8016
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2688 7828 2740 7880
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3332 7828 3384 7837
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 5264 7828 5316 7880
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 9036 7871 9088 7880
rect 9036 7837 9045 7871
rect 9045 7837 9079 7871
rect 9079 7837 9088 7871
rect 9036 7828 9088 7837
rect 11336 7828 11388 7880
rect 12808 7871 12860 7880
rect 4068 7760 4120 7812
rect 12532 7760 12584 7812
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 12992 7828 13044 7880
rect 14556 7871 14608 7880
rect 13728 7760 13780 7812
rect 14556 7837 14565 7871
rect 14565 7837 14599 7871
rect 14599 7837 14608 7871
rect 14556 7828 14608 7837
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 2320 7692 2372 7744
rect 4160 7692 4212 7744
rect 5356 7692 5408 7744
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 11888 7692 11940 7744
rect 12256 7692 12308 7744
rect 17224 7760 17276 7812
rect 15200 7692 15252 7744
rect 3614 7590 3666 7642
rect 3678 7590 3730 7642
rect 3742 7590 3794 7642
rect 3806 7590 3858 7642
rect 8878 7590 8930 7642
rect 8942 7590 8994 7642
rect 9006 7590 9058 7642
rect 9070 7590 9122 7642
rect 14142 7590 14194 7642
rect 14206 7590 14258 7642
rect 14270 7590 14322 7642
rect 14334 7590 14386 7642
rect 2044 7488 2096 7540
rect 4896 7531 4948 7540
rect 2596 7352 2648 7404
rect 3976 7420 4028 7472
rect 3332 7352 3384 7404
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 3056 7284 3108 7336
rect 3976 7284 4028 7336
rect 4344 7284 4396 7336
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 6644 7488 6696 7540
rect 9680 7488 9732 7540
rect 5816 7420 5868 7472
rect 12256 7488 12308 7540
rect 5172 7352 5224 7404
rect 7104 7352 7156 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 7932 7284 7984 7336
rect 12348 7420 12400 7472
rect 8484 7352 8536 7404
rect 11888 7395 11940 7404
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 13912 7488 13964 7540
rect 13728 7352 13780 7404
rect 11704 7284 11756 7336
rect 12348 7284 12400 7336
rect 12716 7327 12768 7336
rect 12716 7293 12750 7327
rect 12750 7293 12768 7327
rect 12716 7284 12768 7293
rect 13176 7284 13228 7336
rect 2872 7148 2924 7200
rect 3516 7148 3568 7200
rect 4712 7148 4764 7200
rect 6736 7148 6788 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 9588 7216 9640 7268
rect 10416 7148 10468 7200
rect 11060 7148 11112 7200
rect 12532 7216 12584 7268
rect 14372 7216 14424 7268
rect 15016 7216 15068 7268
rect 13176 7148 13228 7200
rect 14280 7191 14332 7200
rect 14280 7157 14289 7191
rect 14289 7157 14323 7191
rect 14323 7157 14332 7191
rect 14280 7148 14332 7157
rect 14832 7148 14884 7200
rect 16028 7191 16080 7200
rect 16028 7157 16037 7191
rect 16037 7157 16071 7191
rect 16071 7157 16080 7191
rect 16028 7148 16080 7157
rect 6246 7046 6298 7098
rect 6310 7046 6362 7098
rect 6374 7046 6426 7098
rect 6438 7046 6490 7098
rect 11510 7046 11562 7098
rect 11574 7046 11626 7098
rect 11638 7046 11690 7098
rect 11702 7046 11754 7098
rect 2780 6944 2832 6996
rect 3056 6944 3108 6996
rect 4988 6944 5040 6996
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 3332 6876 3384 6928
rect 6920 6944 6972 6996
rect 7472 6944 7524 6996
rect 7932 6944 7984 6996
rect 12900 6944 12952 6996
rect 13176 6987 13228 6996
rect 13176 6953 13185 6987
rect 13185 6953 13219 6987
rect 13219 6953 13228 6987
rect 13176 6944 13228 6953
rect 14556 6944 14608 6996
rect 2688 6808 2740 6860
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 5356 6808 5408 6860
rect 5816 6808 5868 6860
rect 7012 6876 7064 6928
rect 13820 6876 13872 6928
rect 14372 6876 14424 6928
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 5172 6672 5224 6724
rect 2780 6604 2832 6656
rect 4160 6604 4212 6656
rect 4436 6604 4488 6656
rect 5448 6604 5500 6656
rect 8208 6808 8260 6860
rect 9956 6808 10008 6860
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 11060 6851 11112 6860
rect 11060 6817 11094 6851
rect 11094 6817 11112 6851
rect 11060 6808 11112 6817
rect 14280 6808 14332 6860
rect 14464 6851 14516 6860
rect 14464 6817 14473 6851
rect 14473 6817 14507 6851
rect 14507 6817 14516 6851
rect 14464 6808 14516 6817
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 9220 6783 9272 6792
rect 8668 6672 8720 6724
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 10048 6740 10100 6792
rect 12808 6740 12860 6792
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 14648 6715 14700 6724
rect 14648 6681 14657 6715
rect 14657 6681 14691 6715
rect 14691 6681 14700 6715
rect 14648 6672 14700 6681
rect 9404 6604 9456 6656
rect 9864 6604 9916 6656
rect 10416 6604 10468 6656
rect 12532 6604 12584 6656
rect 15292 6647 15344 6656
rect 15292 6613 15301 6647
rect 15301 6613 15335 6647
rect 15335 6613 15344 6647
rect 15292 6604 15344 6613
rect 3614 6502 3666 6554
rect 3678 6502 3730 6554
rect 3742 6502 3794 6554
rect 3806 6502 3858 6554
rect 8878 6502 8930 6554
rect 8942 6502 8994 6554
rect 9006 6502 9058 6554
rect 9070 6502 9122 6554
rect 14142 6502 14194 6554
rect 14206 6502 14258 6554
rect 14270 6502 14322 6554
rect 14334 6502 14386 6554
rect 5540 6400 5592 6452
rect 6920 6400 6972 6452
rect 8484 6400 8536 6452
rect 5816 6375 5868 6384
rect 5816 6341 5825 6375
rect 5825 6341 5859 6375
rect 5859 6341 5868 6375
rect 5816 6332 5868 6341
rect 6644 6332 6696 6384
rect 9864 6332 9916 6384
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 8668 6264 8720 6316
rect 9588 6264 9640 6316
rect 9680 6264 9732 6316
rect 11244 6400 11296 6452
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 16120 6400 16172 6452
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 2136 6196 2188 6248
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 9772 6196 9824 6248
rect 2228 6128 2280 6180
rect 2688 6128 2740 6180
rect 3424 6060 3476 6112
rect 4896 6128 4948 6180
rect 9404 6128 9456 6180
rect 9496 6128 9548 6180
rect 12440 6264 12492 6316
rect 12348 6196 12400 6248
rect 10048 6128 10100 6180
rect 10232 6171 10284 6180
rect 10232 6137 10266 6171
rect 10266 6137 10284 6171
rect 10232 6128 10284 6137
rect 12072 6128 12124 6180
rect 13912 6239 13964 6248
rect 13912 6205 13946 6239
rect 13946 6205 13964 6239
rect 13912 6196 13964 6205
rect 14188 6196 14240 6248
rect 6920 6060 6972 6112
rect 8300 6060 8352 6112
rect 11152 6060 11204 6112
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12808 6103 12860 6112
rect 12440 6060 12492 6069
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 14188 6060 14240 6112
rect 15016 6103 15068 6112
rect 15016 6069 15025 6103
rect 15025 6069 15059 6103
rect 15059 6069 15068 6103
rect 15016 6060 15068 6069
rect 6246 5958 6298 6010
rect 6310 5958 6362 6010
rect 6374 5958 6426 6010
rect 6438 5958 6490 6010
rect 11510 5958 11562 6010
rect 11574 5958 11626 6010
rect 11638 5958 11690 6010
rect 11702 5958 11754 6010
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 4620 5856 4672 5908
rect 4896 5899 4948 5908
rect 4896 5865 4905 5899
rect 4905 5865 4939 5899
rect 4939 5865 4948 5899
rect 4896 5856 4948 5865
rect 6644 5856 6696 5908
rect 8392 5856 8444 5908
rect 10968 5856 11020 5908
rect 12808 5856 12860 5908
rect 15292 5856 15344 5908
rect 1400 5788 1452 5840
rect 10876 5788 10928 5840
rect 11152 5788 11204 5840
rect 12532 5788 12584 5840
rect 15200 5788 15252 5840
rect 2964 5720 3016 5772
rect 4804 5763 4856 5772
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 4804 5720 4856 5729
rect 10324 5720 10376 5772
rect 10508 5763 10560 5772
rect 10508 5729 10517 5763
rect 10517 5729 10551 5763
rect 10551 5729 10560 5763
rect 10508 5720 10560 5729
rect 2688 5652 2740 5704
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 9588 5652 9640 5704
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 11244 5652 11296 5704
rect 11704 5652 11756 5704
rect 12348 5720 12400 5772
rect 13820 5720 13872 5772
rect 13912 5652 13964 5704
rect 10692 5584 10744 5636
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 6000 5516 6052 5568
rect 10048 5516 10100 5568
rect 10416 5516 10468 5568
rect 15844 5584 15896 5636
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 16028 5559 16080 5568
rect 16028 5525 16037 5559
rect 16037 5525 16071 5559
rect 16071 5525 16080 5559
rect 16028 5516 16080 5525
rect 3614 5414 3666 5466
rect 3678 5414 3730 5466
rect 3742 5414 3794 5466
rect 3806 5414 3858 5466
rect 8878 5414 8930 5466
rect 8942 5414 8994 5466
rect 9006 5414 9058 5466
rect 9070 5414 9122 5466
rect 14142 5414 14194 5466
rect 14206 5414 14258 5466
rect 14270 5414 14322 5466
rect 14334 5414 14386 5466
rect 1676 5312 1728 5364
rect 2964 5312 3016 5364
rect 3332 5244 3384 5296
rect 1584 5176 1636 5228
rect 3424 5176 3476 5228
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 4528 5176 4580 5228
rect 5080 5176 5132 5228
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 9404 5312 9456 5364
rect 12808 5312 12860 5364
rect 13084 5312 13136 5364
rect 10324 5244 10376 5296
rect 11704 5287 11756 5296
rect 2320 5151 2372 5160
rect 2320 5117 2329 5151
rect 2329 5117 2363 5151
rect 2363 5117 2372 5151
rect 2320 5108 2372 5117
rect 2504 5108 2556 5160
rect 5724 5108 5776 5160
rect 10232 5176 10284 5228
rect 10784 5176 10836 5228
rect 5448 5040 5500 5092
rect 8576 5108 8628 5160
rect 9496 5108 9548 5160
rect 11704 5253 11713 5287
rect 11713 5253 11747 5287
rect 11747 5253 11756 5287
rect 11704 5244 11756 5253
rect 12532 5176 12584 5228
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 13176 5176 13228 5228
rect 11796 5108 11848 5160
rect 12992 5151 13044 5160
rect 12992 5117 13001 5151
rect 13001 5117 13035 5151
rect 13035 5117 13044 5151
rect 12992 5108 13044 5117
rect 15660 5108 15712 5160
rect 7012 5040 7064 5092
rect 10508 5040 10560 5092
rect 2964 4972 3016 5024
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 5908 5015 5960 5024
rect 5908 4981 5917 5015
rect 5917 4981 5951 5015
rect 5951 4981 5960 5015
rect 5908 4972 5960 4981
rect 9772 4972 9824 5024
rect 11336 5040 11388 5092
rect 10876 5015 10928 5024
rect 10876 4981 10885 5015
rect 10885 4981 10919 5015
rect 10919 4981 10928 5015
rect 10876 4972 10928 4981
rect 10968 5015 11020 5024
rect 10968 4981 10977 5015
rect 10977 4981 11011 5015
rect 11011 4981 11020 5015
rect 10968 4972 11020 4981
rect 12624 4972 12676 5024
rect 13728 5015 13780 5024
rect 13728 4981 13737 5015
rect 13737 4981 13771 5015
rect 13771 4981 13780 5015
rect 13728 4972 13780 4981
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 16028 5015 16080 5024
rect 16028 4981 16037 5015
rect 16037 4981 16071 5015
rect 16071 4981 16080 5015
rect 16028 4972 16080 4981
rect 6246 4870 6298 4922
rect 6310 4870 6362 4922
rect 6374 4870 6426 4922
rect 6438 4870 6490 4922
rect 11510 4870 11562 4922
rect 11574 4870 11626 4922
rect 11638 4870 11690 4922
rect 11702 4870 11754 4922
rect 3700 4768 3752 4820
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 5908 4768 5960 4820
rect 7564 4768 7616 4820
rect 7656 4768 7708 4820
rect 10876 4768 10928 4820
rect 2136 4675 2188 4684
rect 2136 4641 2145 4675
rect 2145 4641 2179 4675
rect 2179 4641 2188 4675
rect 2136 4632 2188 4641
rect 3424 4632 3476 4684
rect 9772 4700 9824 4752
rect 9864 4700 9916 4752
rect 14096 4768 14148 4820
rect 12808 4700 12860 4752
rect 13268 4700 13320 4752
rect 6736 4632 6788 4684
rect 10324 4675 10376 4684
rect 5816 4607 5868 4616
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 4160 4428 4212 4480
rect 5172 4471 5224 4480
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 5632 4496 5684 4548
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 8208 4607 8260 4616
rect 7012 4564 7064 4573
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 10324 4641 10333 4675
rect 10333 4641 10367 4675
rect 10367 4641 10376 4675
rect 10324 4632 10376 4641
rect 10692 4632 10744 4684
rect 8024 4496 8076 4548
rect 10508 4564 10560 4616
rect 10876 4564 10928 4616
rect 11060 4564 11112 4616
rect 13084 4607 13136 4616
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 12164 4496 12216 4548
rect 7472 4428 7524 4480
rect 7748 4471 7800 4480
rect 7748 4437 7757 4471
rect 7757 4437 7791 4471
rect 7791 4437 7800 4471
rect 7748 4428 7800 4437
rect 9956 4428 10008 4480
rect 11520 4428 11572 4480
rect 16028 4471 16080 4480
rect 16028 4437 16037 4471
rect 16037 4437 16071 4471
rect 16071 4437 16080 4471
rect 16028 4428 16080 4437
rect 3614 4326 3666 4378
rect 3678 4326 3730 4378
rect 3742 4326 3794 4378
rect 3806 4326 3858 4378
rect 8878 4326 8930 4378
rect 8942 4326 8994 4378
rect 9006 4326 9058 4378
rect 9070 4326 9122 4378
rect 14142 4326 14194 4378
rect 14206 4326 14258 4378
rect 14270 4326 14322 4378
rect 14334 4326 14386 4378
rect 2964 4267 3016 4276
rect 2964 4233 2973 4267
rect 2973 4233 3007 4267
rect 3007 4233 3016 4267
rect 2964 4224 3016 4233
rect 3424 4224 3476 4276
rect 5080 4224 5132 4276
rect 6736 4224 6788 4276
rect 7012 4224 7064 4276
rect 8208 4224 8260 4276
rect 2504 4088 2556 4140
rect 3056 4088 3108 4140
rect 7656 4156 7708 4208
rect 2412 4020 2464 4072
rect 5448 4020 5500 4072
rect 7840 4020 7892 4072
rect 8576 4020 8628 4072
rect 10324 4088 10376 4140
rect 8944 4063 8996 4072
rect 8944 4029 8967 4063
rect 8967 4029 8996 4063
rect 11796 4224 11848 4276
rect 13176 4224 13228 4276
rect 13084 4156 13136 4208
rect 13360 4156 13412 4208
rect 15016 4088 15068 4140
rect 15752 4088 15804 4140
rect 11520 4063 11572 4072
rect 8944 4020 8996 4029
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 5816 3952 5868 4004
rect 7196 3952 7248 4004
rect 13636 3952 13688 4004
rect 14924 4020 14976 4072
rect 15384 3952 15436 4004
rect 3148 3884 3200 3936
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 8024 3884 8076 3936
rect 11336 3884 11388 3936
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 14556 3927 14608 3936
rect 12900 3884 12952 3893
rect 14556 3893 14565 3927
rect 14565 3893 14599 3927
rect 14599 3893 14608 3927
rect 14556 3884 14608 3893
rect 15108 3884 15160 3936
rect 16028 3927 16080 3936
rect 16028 3893 16037 3927
rect 16037 3893 16071 3927
rect 16071 3893 16080 3927
rect 16028 3884 16080 3893
rect 6246 3782 6298 3834
rect 6310 3782 6362 3834
rect 6374 3782 6426 3834
rect 6438 3782 6490 3834
rect 11510 3782 11562 3834
rect 11574 3782 11626 3834
rect 11638 3782 11690 3834
rect 11702 3782 11754 3834
rect 5172 3680 5224 3732
rect 5816 3680 5868 3732
rect 8300 3680 8352 3732
rect 5724 3655 5776 3664
rect 756 3476 808 3528
rect 3976 3544 4028 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 5724 3621 5758 3655
rect 5758 3621 5776 3655
rect 5724 3612 5776 3621
rect 8852 3680 8904 3732
rect 7196 3544 7248 3596
rect 6828 3476 6880 3528
rect 2964 3340 3016 3392
rect 3332 3383 3384 3392
rect 3332 3349 3341 3383
rect 3341 3349 3375 3383
rect 3375 3349 3384 3383
rect 3332 3340 3384 3349
rect 3424 3340 3476 3392
rect 7380 3408 7432 3460
rect 9404 3544 9456 3596
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9588 3476 9640 3528
rect 10968 3680 11020 3732
rect 11152 3680 11204 3732
rect 12072 3612 12124 3664
rect 13268 3544 13320 3596
rect 15568 3544 15620 3596
rect 16304 3544 16356 3596
rect 10876 3476 10928 3528
rect 11796 3476 11848 3528
rect 12992 3408 13044 3460
rect 7104 3340 7156 3392
rect 7840 3340 7892 3392
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 8392 3340 8444 3392
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 16028 3383 16080 3392
rect 16028 3349 16037 3383
rect 16037 3349 16071 3383
rect 16071 3349 16080 3383
rect 16028 3340 16080 3349
rect 3614 3238 3666 3290
rect 3678 3238 3730 3290
rect 3742 3238 3794 3290
rect 3806 3238 3858 3290
rect 8878 3238 8930 3290
rect 8942 3238 8994 3290
rect 9006 3238 9058 3290
rect 9070 3238 9122 3290
rect 14142 3238 14194 3290
rect 14206 3238 14258 3290
rect 14270 3238 14322 3290
rect 14334 3238 14386 3290
rect 2780 3136 2832 3188
rect 6828 3136 6880 3188
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 5724 3068 5776 3120
rect 3240 3000 3292 3052
rect 3516 2932 3568 2984
rect 6092 3000 6144 3052
rect 8576 3136 8628 3188
rect 9588 3179 9640 3188
rect 9588 3145 9597 3179
rect 9597 3145 9631 3179
rect 9631 3145 9640 3179
rect 9588 3136 9640 3145
rect 10600 3136 10652 3188
rect 13728 3068 13780 3120
rect 7748 2932 7800 2984
rect 10048 2975 10100 2984
rect 10048 2941 10057 2975
rect 10057 2941 10091 2975
rect 10091 2941 10100 2975
rect 10048 2932 10100 2941
rect 11336 2975 11388 2984
rect 11336 2941 11345 2975
rect 11345 2941 11379 2975
rect 11379 2941 11388 2975
rect 11336 2932 11388 2941
rect 3056 2796 3108 2848
rect 3976 2864 4028 2916
rect 5264 2864 5316 2916
rect 6736 2864 6788 2916
rect 7380 2796 7432 2848
rect 7472 2839 7524 2848
rect 7472 2805 7481 2839
rect 7481 2805 7515 2839
rect 7515 2805 7524 2839
rect 9772 2864 9824 2916
rect 10784 2864 10836 2916
rect 12900 3000 12952 3052
rect 12440 2932 12492 2984
rect 12992 2932 13044 2984
rect 12716 2864 12768 2916
rect 13268 2864 13320 2916
rect 7472 2796 7524 2805
rect 14004 2796 14056 2848
rect 14924 2796 14976 2848
rect 15108 2839 15160 2848
rect 15108 2805 15117 2839
rect 15117 2805 15151 2839
rect 15151 2805 15160 2839
rect 15108 2796 15160 2805
rect 16028 2839 16080 2848
rect 16028 2805 16037 2839
rect 16037 2805 16071 2839
rect 16071 2805 16080 2839
rect 16028 2796 16080 2805
rect 6246 2694 6298 2746
rect 6310 2694 6362 2746
rect 6374 2694 6426 2746
rect 6438 2694 6490 2746
rect 11510 2694 11562 2746
rect 11574 2694 11626 2746
rect 11638 2694 11690 2746
rect 11702 2694 11754 2746
rect 7472 2592 7524 2644
rect 8300 2592 8352 2644
rect 8392 2524 8444 2576
rect 2412 2456 2464 2508
rect 4804 2456 4856 2508
rect 7932 2456 7984 2508
rect 11980 2456 12032 2508
rect 15844 2499 15896 2508
rect 15844 2465 15853 2499
rect 15853 2465 15887 2499
rect 15887 2465 15896 2499
rect 15844 2456 15896 2465
rect 8024 2388 8076 2440
rect 11244 2388 11296 2440
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 8208 2252 8260 2304
rect 9220 2252 9272 2304
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 14832 2252 14884 2261
rect 16028 2295 16080 2304
rect 16028 2261 16037 2295
rect 16037 2261 16071 2295
rect 16071 2261 16080 2295
rect 16028 2252 16080 2261
rect 3614 2150 3666 2202
rect 3678 2150 3730 2202
rect 3742 2150 3794 2202
rect 3806 2150 3858 2202
rect 8878 2150 8930 2202
rect 8942 2150 8994 2202
rect 9006 2150 9058 2202
rect 9070 2150 9122 2202
rect 14142 2150 14194 2202
rect 14206 2150 14258 2202
rect 14270 2150 14322 2202
rect 14334 2150 14386 2202
<< metal2 >>
rect 4802 16688 4858 16697
rect 4802 16623 4858 16632
rect 14922 16688 14978 16697
rect 14922 16623 14978 16632
rect 3054 16280 3110 16289
rect 3054 16215 3110 16224
rect 2318 14240 2374 14249
rect 2318 14175 2374 14184
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 1964 11898 1992 12242
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1964 10606 1992 11086
rect 2148 10810 2176 12174
rect 2332 11801 2360 14175
rect 2962 13832 3018 13841
rect 2962 13767 3018 13776
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2318 11792 2374 11801
rect 2228 11756 2280 11762
rect 2318 11727 2374 11736
rect 2228 11698 2280 11704
rect 2240 11218 2268 11698
rect 2332 11694 2360 11727
rect 2320 11688 2372 11694
rect 2884 11665 2912 12310
rect 2976 11898 3004 13767
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2320 11630 2372 11636
rect 2870 11656 2926 11665
rect 2870 11591 2926 11600
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2240 10674 2268 11154
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2056 9722 2084 10406
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2148 9178 2176 10406
rect 2424 10266 2452 11494
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2332 9042 2360 9590
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2424 9081 2452 9318
rect 2410 9072 2466 9081
rect 2320 9036 2372 9042
rect 2410 9007 2466 9016
rect 2320 8978 2372 8984
rect 2332 8838 2360 8978
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 5846 1440 6802
rect 1400 5840 1452 5846
rect 1400 5782 1452 5788
rect 1596 5681 1624 8230
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7546 2084 7822
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6254 2176 6734
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1596 5234 1624 5510
rect 1688 5370 1716 6190
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 2148 4690 2176 6190
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 3641 1624 4422
rect 1582 3632 1638 3641
rect 1582 3567 1638 3576
rect 756 3528 808 3534
rect 756 3470 808 3476
rect 768 480 796 3470
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 1465 2176 2246
rect 2134 1456 2190 1465
rect 2134 1391 2190 1400
rect 2240 480 2268 6122
rect 2332 5166 2360 7686
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2424 4078 2452 9007
rect 2504 8968 2556 8974
rect 2502 8936 2504 8945
rect 2556 8936 2558 8945
rect 2502 8871 2558 8880
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2516 5166 2544 8774
rect 2608 7410 2636 10950
rect 2686 10568 2742 10577
rect 2686 10503 2742 10512
rect 2700 10266 2728 10503
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2700 10130 2728 10202
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2700 9586 2728 9930
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2792 8537 2820 11494
rect 2884 10266 2912 11591
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2976 10305 3004 10474
rect 2962 10296 3018 10305
rect 2872 10260 2924 10266
rect 2962 10231 3018 10240
rect 2872 10202 2924 10208
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2976 9976 3004 10066
rect 3068 10044 3096 16215
rect 3146 15872 3202 15881
rect 3146 15807 3202 15816
rect 3160 11014 3188 15807
rect 3882 15464 3938 15473
rect 3882 15399 3938 15408
rect 3896 15298 3924 15399
rect 3884 15292 3936 15298
rect 3884 15234 3936 15240
rect 3514 15056 3570 15065
rect 3514 14991 3570 15000
rect 3528 14822 3556 14991
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3588 14172 3884 14192
rect 3644 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3666 14118 3668 14170
rect 3730 14118 3742 14170
rect 3804 14118 3806 14170
rect 3644 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3588 14096 3884 14116
rect 4158 13288 4214 13297
rect 4158 13223 4214 13232
rect 3588 13084 3884 13104
rect 3644 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3666 13030 3668 13082
rect 3730 13030 3742 13082
rect 3804 13030 3806 13082
rect 3644 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3588 13008 3884 13028
rect 3514 12880 3570 12889
rect 3514 12815 3570 12824
rect 3528 12714 3556 12815
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 12481 4108 12582
rect 4066 12472 4122 12481
rect 4066 12407 4122 12416
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3146 10840 3202 10849
rect 3146 10775 3202 10784
rect 3160 10266 3188 10775
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3068 10016 3188 10044
rect 2976 9948 3096 9976
rect 2870 9888 2926 9897
rect 2870 9823 2926 9832
rect 2884 9382 2912 9823
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2778 8528 2834 8537
rect 2778 8463 2834 8472
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2700 6866 2728 7822
rect 2884 7290 2912 9318
rect 2792 7262 2912 7290
rect 2792 7002 2820 7262
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 6186 2728 6802
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2700 5710 2728 6122
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2516 4146 2544 5102
rect 2792 4457 2820 6598
rect 2884 4865 2912 7142
rect 2976 6497 3004 9658
rect 3068 7342 3096 9948
rect 3160 9110 3188 10016
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3160 8090 3188 8842
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 2962 6488 3018 6497
rect 2962 6423 3018 6432
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2976 5370 3004 5714
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2870 4856 2926 4865
rect 2870 4791 2926 4800
rect 2778 4448 2834 4457
rect 2778 4383 2834 4392
rect 2976 4282 3004 4966
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 3068 4146 3096 6938
rect 3160 5914 3188 7890
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2424 2514 2452 4014
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 754 0 810 480
rect 2226 0 2282 480
rect 2792 241 2820 3130
rect 2872 2304 2924 2310
rect 2870 2272 2872 2281
rect 2924 2272 2926 2281
rect 2870 2207 2926 2216
rect 2976 1873 3004 3334
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2962 1864 3018 1873
rect 2962 1799 3018 1808
rect 3068 1057 3096 2790
rect 3054 1048 3110 1057
rect 3054 983 3110 992
rect 3160 649 3188 3878
rect 3252 3058 3280 12038
rect 3344 11762 3372 12174
rect 3422 12064 3478 12073
rect 3422 11999 3478 12008
rect 3436 11830 3464 11999
rect 3588 11996 3884 12016
rect 3644 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3666 11942 3668 11994
rect 3730 11942 3742 11994
rect 3804 11942 3806 11994
rect 3644 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3588 11920 3884 11940
rect 3988 11898 4016 12242
rect 4172 12209 4200 13223
rect 4252 12232 4304 12238
rect 4158 12200 4214 12209
rect 4252 12174 4304 12180
rect 4158 12135 4214 12144
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3344 11354 3372 11698
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3344 10538 3372 11290
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3330 10296 3386 10305
rect 3330 10231 3386 10240
rect 3344 9518 3372 10231
rect 3528 9625 3556 11834
rect 4172 11744 4200 12135
rect 3988 11716 4200 11744
rect 3588 10908 3884 10928
rect 3644 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3666 10854 3668 10906
rect 3730 10854 3742 10906
rect 3804 10854 3806 10906
rect 3644 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3588 10832 3884 10852
rect 3588 9820 3884 9840
rect 3644 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3666 9766 3668 9818
rect 3730 9766 3742 9818
rect 3804 9766 3806 9818
rect 3644 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3588 9744 3884 9764
rect 3514 9616 3570 9625
rect 3514 9551 3570 9560
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3344 9042 3372 9454
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3528 8974 3556 9386
rect 3988 9058 4016 11716
rect 4066 11248 4122 11257
rect 4066 11183 4122 11192
rect 4080 11082 4108 11183
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4264 10810 4292 12174
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4356 11354 4384 11494
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4448 10810 4476 11494
rect 4816 10810 4844 16623
rect 13174 15872 13230 15881
rect 13174 15807 13230 15816
rect 6552 15292 6604 15298
rect 6552 15234 6604 15240
rect 6220 14716 6516 14736
rect 6276 14714 6300 14716
rect 6356 14714 6380 14716
rect 6436 14714 6460 14716
rect 6298 14662 6300 14714
rect 6362 14662 6374 14714
rect 6436 14662 6438 14714
rect 6276 14660 6300 14662
rect 6356 14660 6380 14662
rect 6436 14660 6460 14662
rect 5814 14648 5870 14657
rect 6220 14640 6516 14660
rect 5814 14583 5870 14592
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 11354 4936 11494
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5000 11286 5028 11630
rect 4988 11280 5040 11286
rect 4986 11248 4988 11257
rect 5040 11248 5042 11257
rect 4986 11183 5042 11192
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4080 10441 4108 10678
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4264 10198 4292 10746
rect 4816 10674 4844 10746
rect 5276 10674 5304 11086
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4080 9722 4108 9862
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 3988 9030 4108 9058
rect 4172 9042 4200 9386
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4264 9042 4292 9114
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3344 8634 3372 8842
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3344 7410 3372 7822
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3344 6934 3372 7346
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3344 5710 3372 6870
rect 3436 6225 3464 8774
rect 3528 8634 3556 8910
rect 3588 8732 3884 8752
rect 3644 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3666 8678 3668 8730
rect 3730 8678 3742 8730
rect 3804 8678 3806 8730
rect 3644 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3588 8656 3884 8676
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3896 8362 3924 8502
rect 3988 8498 4016 8910
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3896 7732 3924 8298
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 7857 4016 8230
rect 4080 7954 4108 9030
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3974 7848 4030 7857
rect 3974 7783 4030 7792
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3896 7704 4016 7732
rect 3588 7644 3884 7664
rect 3644 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3666 7590 3668 7642
rect 3730 7590 3742 7642
rect 3804 7590 3806 7642
rect 3644 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3588 7568 3884 7588
rect 3988 7478 4016 7704
rect 3976 7472 4028 7478
rect 4080 7449 4108 7754
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 3976 7414 4028 7420
rect 4066 7440 4122 7449
rect 4172 7410 4200 7686
rect 4066 7375 4122 7384
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3422 6216 3478 6225
rect 3422 6151 3478 6160
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3344 5302 3372 5646
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 3436 5234 3464 6054
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3436 4282 3464 4626
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3344 2689 3372 3334
rect 3436 3097 3464 3334
rect 3422 3088 3478 3097
rect 3422 3023 3478 3032
rect 3528 2990 3556 7142
rect 3588 6556 3884 6576
rect 3644 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3666 6502 3668 6554
rect 3730 6502 3742 6554
rect 3804 6502 3806 6554
rect 3644 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3588 6480 3884 6500
rect 3588 5468 3884 5488
rect 3644 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3666 5414 3668 5466
rect 3730 5414 3742 5466
rect 3804 5414 3806 5466
rect 3644 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3588 5392 3884 5412
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3712 4826 3740 5170
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3588 4380 3884 4400
rect 3644 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3666 4326 3668 4378
rect 3730 4326 3742 4378
rect 3804 4326 3806 4378
rect 3644 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3588 4304 3884 4324
rect 3988 3602 4016 7278
rect 4264 7256 4292 8774
rect 4356 7342 4384 9114
rect 4526 8936 4582 8945
rect 4526 8871 4582 8880
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4080 7228 4292 7256
rect 4080 7177 4108 7228
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4066 5264 4122 5273
rect 4172 5250 4200 6598
rect 4448 6254 4476 6598
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4122 5222 4200 5250
rect 4540 5234 4568 8871
rect 4632 5914 4660 10202
rect 4724 9722 4752 10474
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 10266 5304 10406
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4816 9722 4844 9862
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4710 9616 4766 9625
rect 4710 9551 4766 9560
rect 4724 7206 4752 9551
rect 4816 8974 4844 9658
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4908 8650 4936 8978
rect 5092 8906 5120 10202
rect 5552 9654 5580 12174
rect 5828 11694 5856 14583
rect 6220 13628 6516 13648
rect 6276 13626 6300 13628
rect 6356 13626 6380 13628
rect 6436 13626 6460 13628
rect 6298 13574 6300 13626
rect 6362 13574 6374 13626
rect 6436 13574 6438 13626
rect 6276 13572 6300 13574
rect 6356 13572 6380 13574
rect 6436 13572 6460 13574
rect 6220 13552 6516 13572
rect 6220 12540 6516 12560
rect 6276 12538 6300 12540
rect 6356 12538 6380 12540
rect 6436 12538 6460 12540
rect 6298 12486 6300 12538
rect 6362 12486 6374 12538
rect 6436 12486 6438 12538
rect 6276 12484 6300 12486
rect 6356 12484 6380 12486
rect 6436 12484 6460 12486
rect 6220 12464 6516 12484
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4908 8622 5028 8650
rect 5000 8566 5028 8622
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5184 8498 5212 8978
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4908 7546 4936 7890
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 5000 7002 5028 7822
rect 5184 7410 5212 8434
rect 5276 8430 5304 8774
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5276 7886 5304 8366
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5368 7750 5396 9454
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5184 6730 5212 7346
rect 5368 6866 5396 7686
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 4908 5914 4936 6122
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4528 5228 4580 5234
rect 4066 5199 4122 5208
rect 4528 5170 4580 5176
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4066 4040 4122 4049
rect 4172 4026 4200 4422
rect 4122 3998 4200 4026
rect 4066 3975 4122 3984
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3588 3292 3884 3312
rect 3644 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3666 3238 3668 3290
rect 3730 3238 3742 3290
rect 3804 3238 3806 3290
rect 3644 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3588 3216 3884 3236
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3330 2680 3386 2689
rect 3330 2615 3386 2624
rect 3588 2204 3884 2224
rect 3644 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3666 2150 3668 2202
rect 3730 2150 3742 2202
rect 3804 2150 3806 2202
rect 3644 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3588 2128 3884 2148
rect 3988 1442 4016 2858
rect 4816 2514 4844 5714
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5092 5234 5120 5646
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5092 4282 5120 5170
rect 5460 5098 5488 6598
rect 5552 6458 5580 6734
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5184 3738 5212 4422
rect 5460 4078 5488 5034
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4826 5580 4966
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5644 4554 5672 9386
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5736 9042 5764 9318
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5828 7478 5856 11018
rect 6012 10606 6040 11766
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5828 6390 5856 6802
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6012 5234 6040 5510
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5460 3602 5488 4014
rect 5736 3670 5764 5102
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4826 5948 4966
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5828 4010 5856 4558
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5828 3738 5856 3946
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5736 3126 5764 3606
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 6104 3058 6132 12038
rect 6220 11452 6516 11472
rect 6276 11450 6300 11452
rect 6356 11450 6380 11452
rect 6436 11450 6460 11452
rect 6298 11398 6300 11450
rect 6362 11398 6374 11450
rect 6436 11398 6438 11450
rect 6276 11396 6300 11398
rect 6356 11396 6380 11398
rect 6436 11396 6460 11398
rect 6220 11376 6516 11396
rect 6220 10364 6516 10384
rect 6276 10362 6300 10364
rect 6356 10362 6380 10364
rect 6436 10362 6460 10364
rect 6298 10310 6300 10362
rect 6362 10310 6374 10362
rect 6436 10310 6438 10362
rect 6276 10308 6300 10310
rect 6356 10308 6380 10310
rect 6436 10308 6460 10310
rect 6220 10288 6516 10308
rect 6220 9276 6516 9296
rect 6276 9274 6300 9276
rect 6356 9274 6380 9276
rect 6436 9274 6460 9276
rect 6298 9222 6300 9274
rect 6362 9222 6374 9274
rect 6436 9222 6438 9274
rect 6276 9220 6300 9222
rect 6356 9220 6380 9222
rect 6436 9220 6460 9222
rect 6220 9200 6516 9220
rect 6220 8188 6516 8208
rect 6276 8186 6300 8188
rect 6356 8186 6380 8188
rect 6436 8186 6460 8188
rect 6298 8134 6300 8186
rect 6362 8134 6374 8186
rect 6436 8134 6438 8186
rect 6276 8132 6300 8134
rect 6356 8132 6380 8134
rect 6436 8132 6460 8134
rect 6220 8112 6516 8132
rect 6220 7100 6516 7120
rect 6276 7098 6300 7100
rect 6356 7098 6380 7100
rect 6436 7098 6460 7100
rect 6298 7046 6300 7098
rect 6362 7046 6374 7098
rect 6436 7046 6438 7098
rect 6276 7044 6300 7046
rect 6356 7044 6380 7046
rect 6436 7044 6460 7046
rect 6220 7024 6516 7044
rect 6564 7018 6592 15234
rect 11888 15224 11940 15230
rect 11888 15166 11940 15172
rect 10598 15056 10654 15065
rect 10598 14991 10654 15000
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 8852 14172 9148 14192
rect 8908 14170 8932 14172
rect 8988 14170 9012 14172
rect 9068 14170 9092 14172
rect 8930 14118 8932 14170
rect 8994 14118 9006 14170
rect 9068 14118 9070 14170
rect 8908 14116 8932 14118
rect 8988 14116 9012 14118
rect 9068 14116 9092 14118
rect 8852 14096 9148 14116
rect 8852 13084 9148 13104
rect 8908 13082 8932 13084
rect 8988 13082 9012 13084
rect 9068 13082 9092 13084
rect 8930 13030 8932 13082
rect 8994 13030 9006 13082
rect 9068 13030 9070 13082
rect 8908 13028 8932 13030
rect 8988 13028 9012 13030
rect 9068 13028 9092 13030
rect 8852 13008 9148 13028
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7668 12306 7696 12650
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 6656 11898 6684 12242
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6656 10674 6684 11154
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6748 9722 6776 11222
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6748 9518 6776 9658
rect 6840 9654 6868 11018
rect 7392 10690 7420 12242
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7484 11642 7512 12038
rect 7668 11762 7696 12038
rect 7852 11830 7880 12106
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7840 11688 7892 11694
rect 7484 11636 7840 11642
rect 7484 11630 7892 11636
rect 7484 11614 7880 11630
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7838 11520 7894 11529
rect 7392 10662 7512 10690
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6932 9450 6960 9862
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6840 8634 6868 8910
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 7546 6684 7890
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6564 6990 6684 7018
rect 6656 6390 6684 6990
rect 6748 6882 6776 7142
rect 6932 7002 6960 8298
rect 7024 7290 7052 10474
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7116 9722 7144 9930
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7116 9518 7144 9658
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7300 9382 7328 10406
rect 7392 10198 7420 10542
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7116 8634 7144 9046
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7116 8294 7144 8570
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7116 7410 7144 7890
rect 7208 7886 7236 8366
rect 7300 8090 7328 9114
rect 7392 8945 7420 9454
rect 7378 8936 7434 8945
rect 7378 8871 7434 8880
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7392 7886 7420 8434
rect 7484 8090 7512 10662
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7380 7880 7432 7886
rect 7432 7840 7512 7868
rect 7380 7822 7432 7828
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7024 7262 7144 7290
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7012 6928 7064 6934
rect 6748 6876 7012 6882
rect 6748 6870 7064 6876
rect 6748 6854 7052 6870
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6220 6012 6516 6032
rect 6276 6010 6300 6012
rect 6356 6010 6380 6012
rect 6436 6010 6460 6012
rect 6298 5958 6300 6010
rect 6362 5958 6374 6010
rect 6436 5958 6438 6010
rect 6276 5956 6300 5958
rect 6356 5956 6380 5958
rect 6436 5956 6460 5958
rect 6220 5936 6516 5956
rect 6656 5914 6684 6326
rect 6932 6118 6960 6394
rect 6920 6112 6972 6118
rect 6840 6072 6920 6100
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6220 4924 6516 4944
rect 6276 4922 6300 4924
rect 6356 4922 6380 4924
rect 6436 4922 6460 4924
rect 6298 4870 6300 4922
rect 6362 4870 6374 4922
rect 6436 4870 6438 4922
rect 6276 4868 6300 4870
rect 6356 4868 6380 4870
rect 6436 4868 6460 4870
rect 6220 4848 6516 4868
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6748 4282 6776 4626
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6220 3836 6516 3856
rect 6276 3834 6300 3836
rect 6356 3834 6380 3836
rect 6436 3834 6460 3836
rect 6298 3782 6300 3834
rect 6362 3782 6374 3834
rect 6436 3782 6438 3834
rect 6276 3780 6300 3782
rect 6356 3780 6380 3782
rect 6436 3780 6460 3782
rect 6220 3760 6516 3780
rect 6840 3534 6868 6072
rect 6920 6054 6972 6060
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7024 5098 7052 5646
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 7024 4622 7052 5034
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6840 3194 6868 3470
rect 7024 3194 7052 4218
rect 7116 3398 7144 7262
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 4010 7236 7142
rect 7392 6322 7420 7346
rect 7484 7002 7512 7840
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7576 6882 7604 11494
rect 7838 11455 7894 11464
rect 7852 10674 7880 11455
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7852 10062 7880 10610
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7668 9178 7696 9998
rect 7852 9722 7880 9998
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7748 9104 7800 9110
rect 7746 9072 7748 9081
rect 7800 9072 7802 9081
rect 7746 9007 7802 9016
rect 7944 8566 7972 12378
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 8024 12232 8076 12238
rect 8208 12232 8260 12238
rect 8024 12174 8076 12180
rect 8206 12200 8208 12209
rect 8260 12200 8262 12209
rect 8036 11762 8064 12174
rect 8206 12135 8262 12144
rect 8852 11996 9148 12016
rect 8908 11994 8932 11996
rect 8988 11994 9012 11996
rect 9068 11994 9092 11996
rect 8930 11942 8932 11994
rect 8994 11942 9006 11994
rect 9068 11942 9070 11994
rect 8908 11940 8932 11942
rect 8988 11940 9012 11942
rect 9068 11940 9092 11942
rect 8852 11920 9148 11940
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8036 11529 8064 11698
rect 8022 11520 8078 11529
rect 8022 11455 8078 11464
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8298 11248 8354 11257
rect 8298 11183 8300 11192
rect 8352 11183 8354 11192
rect 8300 11154 8352 11160
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8128 10062 8156 10406
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8220 10044 8248 10678
rect 8772 10606 8800 11290
rect 8864 11286 8892 11698
rect 9048 11354 9076 11766
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9232 11286 9260 12310
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9324 11558 9352 12038
rect 9402 11792 9458 11801
rect 9402 11727 9458 11736
rect 9416 11694 9444 11727
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 8852 10908 9148 10928
rect 8908 10906 8932 10908
rect 8988 10906 9012 10908
rect 9068 10906 9092 10908
rect 8930 10854 8932 10906
rect 8994 10854 9006 10906
rect 9068 10854 9070 10906
rect 8908 10852 8932 10854
rect 8988 10852 9012 10854
rect 9068 10852 9092 10854
rect 8852 10832 9148 10852
rect 8760 10600 8812 10606
rect 9220 10600 9272 10606
rect 8760 10542 8812 10548
rect 9218 10568 9220 10577
rect 9772 10600 9824 10606
rect 9272 10568 9274 10577
rect 9772 10542 9824 10548
rect 9218 10503 9274 10512
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8772 10130 8800 10406
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8484 10056 8536 10062
rect 8220 10016 8484 10044
rect 8220 9330 8248 10016
rect 8484 9998 8536 10004
rect 8680 9654 8708 10066
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8574 9480 8630 9489
rect 8574 9415 8630 9424
rect 8036 9302 8248 9330
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7484 6854 7604 6882
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7484 4486 7512 6854
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7576 4826 7604 5646
rect 7668 4826 7696 8026
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7944 7002 7972 7278
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 8036 6746 8064 9302
rect 8208 9172 8260 9178
rect 8128 9132 8208 9160
rect 8128 8362 8156 9132
rect 8208 9114 8260 9120
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8537 8340 8910
rect 8298 8528 8354 8537
rect 8298 8463 8354 8472
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8220 6769 8248 6802
rect 7852 6718 8064 6746
rect 8206 6760 8262 6769
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7668 4214 7696 4762
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7208 3602 7236 3946
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 3712 1414 4016 1442
rect 3146 640 3202 649
rect 3146 575 3202 584
rect 3712 480 3740 1414
rect 5276 480 5304 2858
rect 6220 2748 6516 2768
rect 6276 2746 6300 2748
rect 6356 2746 6380 2748
rect 6436 2746 6460 2748
rect 6298 2694 6300 2746
rect 6362 2694 6374 2746
rect 6436 2694 6438 2746
rect 6276 2692 6300 2694
rect 6356 2692 6380 2694
rect 6436 2692 6460 2694
rect 6220 2672 6516 2692
rect 6748 480 6776 2858
rect 7392 2854 7420 3402
rect 7760 2990 7788 4422
rect 7852 4078 7880 6718
rect 8206 6695 8262 6704
rect 8312 6118 8340 8463
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 7840 4072 7892 4078
rect 7892 4032 7972 4060
rect 7840 4014 7892 4020
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 3398 7880 3878
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7484 2650 7512 2790
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7944 2514 7972 4032
rect 8036 3942 8064 4490
rect 8220 4282 8248 4558
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8036 2446 8064 3878
rect 8312 3738 8340 6054
rect 8404 5914 8432 7686
rect 8496 7410 8524 8978
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8496 6458 8524 7346
rect 8588 6798 8616 9415
rect 8772 8090 8800 9862
rect 8852 9820 9148 9840
rect 8908 9818 8932 9820
rect 8988 9818 9012 9820
rect 9068 9818 9092 9820
rect 8930 9766 8932 9818
rect 8994 9766 9006 9818
rect 9068 9766 9070 9818
rect 8908 9764 8932 9766
rect 8988 9764 9012 9766
rect 9068 9764 9092 9766
rect 8852 9744 9148 9764
rect 9232 9586 9260 9998
rect 9324 9926 9352 10474
rect 9784 10470 9812 10542
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9784 10062 9812 10406
rect 10060 10198 10088 10406
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9126 9480 9182 9489
rect 9126 9415 9182 9424
rect 9140 9382 9168 9415
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9048 8820 9076 9318
rect 9232 8974 9260 9522
rect 9784 9042 9812 9998
rect 10060 9586 10088 10134
rect 10336 9761 10364 14758
rect 10612 10538 10640 14991
rect 11484 14716 11780 14736
rect 11540 14714 11564 14716
rect 11620 14714 11644 14716
rect 11700 14714 11724 14716
rect 11562 14662 11564 14714
rect 11626 14662 11638 14714
rect 11700 14662 11702 14714
rect 11540 14660 11564 14662
rect 11620 14660 11644 14662
rect 11700 14660 11724 14662
rect 11484 14640 11780 14660
rect 11484 13628 11780 13648
rect 11540 13626 11564 13628
rect 11620 13626 11644 13628
rect 11700 13626 11724 13628
rect 11562 13574 11564 13626
rect 11626 13574 11638 13626
rect 11700 13574 11702 13626
rect 11540 13572 11564 13574
rect 11620 13572 11644 13574
rect 11700 13572 11724 13574
rect 11484 13552 11780 13572
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10414 9616 10470 9625
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9048 8792 9352 8820
rect 8852 8732 9148 8752
rect 8908 8730 8932 8732
rect 8988 8730 9012 8732
rect 9068 8730 9092 8732
rect 8930 8678 8932 8730
rect 8994 8678 9006 8730
rect 9068 8678 9070 8730
rect 8908 8676 8932 8678
rect 8988 8676 9012 8678
rect 9068 8676 9092 8678
rect 8852 8656 9148 8676
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 9048 7886 9076 8298
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8852 7644 9148 7664
rect 8908 7642 8932 7644
rect 8988 7642 9012 7644
rect 9068 7642 9092 7644
rect 8930 7590 8932 7642
rect 8994 7590 9006 7642
rect 9068 7590 9070 7642
rect 8908 7588 8932 7590
rect 8988 7588 9012 7590
rect 9068 7588 9092 7590
rect 8852 7568 9148 7588
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 9220 6792 9272 6798
rect 9324 6769 9352 8792
rect 9784 8430 9812 8978
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9864 8560 9916 8566
rect 9862 8528 9864 8537
rect 9916 8528 9918 8537
rect 9862 8463 9918 8472
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9600 7274 9628 8230
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9220 6734 9272 6740
rect 9310 6760 9366 6769
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8588 5386 8616 6734
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8680 6322 8708 6666
rect 8852 6556 9148 6576
rect 8908 6554 8932 6556
rect 8988 6554 9012 6556
rect 9068 6554 9092 6556
rect 8930 6502 8932 6554
rect 8994 6502 9006 6554
rect 9068 6502 9070 6554
rect 8908 6500 8932 6502
rect 8988 6500 9012 6502
rect 9068 6500 9092 6502
rect 8852 6480 9148 6500
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8852 5468 9148 5488
rect 8908 5466 8932 5468
rect 8988 5466 9012 5468
rect 9068 5466 9092 5468
rect 8930 5414 8932 5466
rect 8994 5414 9006 5466
rect 9068 5414 9070 5466
rect 8908 5412 8932 5414
rect 8988 5412 9012 5414
rect 9068 5412 9092 5414
rect 8852 5392 9148 5412
rect 8588 5358 8708 5386
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8588 4078 8616 5102
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8312 2650 8340 3334
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2582 8432 3334
rect 8588 3194 8616 4014
rect 8680 3720 8708 5358
rect 8852 4380 9148 4400
rect 8908 4378 8932 4380
rect 8988 4378 9012 4380
rect 9068 4378 9092 4380
rect 8930 4326 8932 4378
rect 8994 4326 9006 4378
rect 9068 4326 9070 4378
rect 8908 4324 8932 4326
rect 8988 4324 9012 4326
rect 9068 4324 9092 4326
rect 8852 4304 9148 4324
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8852 3732 8904 3738
rect 8680 3692 8852 3720
rect 8852 3674 8904 3680
rect 8956 3534 8984 4014
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8852 3292 9148 3312
rect 8908 3290 8932 3292
rect 8988 3290 9012 3292
rect 9068 3290 9092 3292
rect 8930 3238 8932 3290
rect 8994 3238 9006 3290
rect 9068 3238 9070 3290
rect 8908 3236 8932 3238
rect 8988 3236 9012 3238
rect 9068 3236 9092 3238
rect 8852 3216 9148 3236
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 9232 2310 9260 6734
rect 9310 6695 9366 6704
rect 9324 5352 9352 6695
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9416 6186 9444 6598
rect 9600 6322 9628 7210
rect 9692 6322 9720 7482
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9404 5364 9456 5370
rect 9324 5324 9404 5352
rect 9404 5306 9456 5312
rect 9416 3602 9444 5306
rect 9508 5166 9536 6122
rect 9600 5710 9628 6258
rect 9784 6254 9812 7686
rect 9876 6662 9904 8298
rect 9968 8090 9996 8774
rect 10244 8090 10272 9318
rect 10336 8430 10364 9590
rect 10414 9551 10470 9560
rect 10508 9580 10560 9586
rect 10428 9110 10456 9551
rect 10508 9522 10560 9528
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10520 8974 10548 9522
rect 10690 9480 10746 9489
rect 10690 9415 10692 9424
rect 10744 9415 10746 9424
rect 10692 9386 10744 9392
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9081 10640 9318
rect 10598 9072 10654 9081
rect 10598 9007 10654 9016
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10520 8498 10548 8910
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10796 8430 10824 12582
rect 11484 12540 11780 12560
rect 11540 12538 11564 12540
rect 11620 12538 11644 12540
rect 11700 12538 11724 12540
rect 11562 12486 11564 12538
rect 11626 12486 11638 12538
rect 11700 12486 11702 12538
rect 11540 12484 11564 12486
rect 11620 12484 11644 12486
rect 11700 12484 11724 12486
rect 11484 12464 11780 12484
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11348 10538 11376 11698
rect 11484 11452 11780 11472
rect 11540 11450 11564 11452
rect 11620 11450 11644 11452
rect 11700 11450 11724 11452
rect 11562 11398 11564 11450
rect 11626 11398 11638 11450
rect 11700 11398 11702 11450
rect 11540 11396 11564 11398
rect 11620 11396 11644 11398
rect 11700 11396 11724 11398
rect 11484 11376 11780 11396
rect 11900 11218 11928 15166
rect 13082 13288 13138 13297
rect 13082 13223 13138 13232
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11900 10606 11928 10746
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11484 10364 11780 10384
rect 11540 10362 11564 10364
rect 11620 10362 11644 10364
rect 11700 10362 11724 10364
rect 11562 10310 11564 10362
rect 11626 10310 11638 10362
rect 11700 10310 11702 10362
rect 11540 10308 11564 10310
rect 11620 10308 11644 10310
rect 11700 10308 11724 10310
rect 11484 10288 11780 10308
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11058 9752 11114 9761
rect 11058 9687 11114 9696
rect 11072 9636 11100 9687
rect 10980 9608 11100 9636
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 9956 7336 10008 7342
rect 10008 7296 10088 7324
rect 9956 7278 10008 7284
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9784 4758 9812 4966
rect 9876 4758 9904 6326
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9968 4486 9996 6802
rect 10060 6798 10088 7296
rect 10152 6866 10180 7890
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6186 10088 6734
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9600 3194 9628 3470
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 10060 2990 10088 5510
rect 10244 5234 10272 6122
rect 10336 5778 10364 8366
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 7206 10456 8230
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10428 5574 10456 6598
rect 10888 5846 10916 9522
rect 10980 9500 11008 9608
rect 10980 9472 11100 9500
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 9042 11008 9318
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 11072 8022 11100 9472
rect 11256 9160 11284 9862
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11484 9276 11780 9296
rect 11540 9274 11564 9276
rect 11620 9274 11644 9276
rect 11700 9274 11724 9276
rect 11562 9222 11564 9274
rect 11626 9222 11638 9274
rect 11700 9222 11702 9274
rect 11540 9220 11564 9222
rect 11620 9220 11644 9222
rect 11700 9220 11724 9222
rect 11484 9200 11780 9220
rect 11256 9132 11376 9160
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 5914 11008 7686
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6866 11100 7142
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10520 5386 10548 5714
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10336 5358 10548 5386
rect 10336 5302 10364 5358
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10336 4146 10364 4626
rect 10520 4622 10548 5034
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10612 3194 10640 5646
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10704 4690 10732 5578
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10796 2922 10824 5170
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10888 4826 10916 4966
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 3534 10916 4558
rect 10980 3738 11008 4966
rect 11072 4622 11100 6802
rect 11164 6118 11192 8434
rect 11256 6458 11284 8978
rect 11348 8498 11376 9132
rect 11518 8528 11574 8537
rect 11336 8492 11388 8498
rect 11518 8463 11574 8472
rect 11336 8434 11388 8440
rect 11348 7886 11376 8434
rect 11532 8362 11560 8463
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11484 8188 11780 8208
rect 11540 8186 11564 8188
rect 11620 8186 11644 8188
rect 11700 8186 11724 8188
rect 11562 8134 11564 8186
rect 11626 8134 11638 8186
rect 11700 8134 11702 8186
rect 11540 8132 11564 8134
rect 11620 8132 11644 8134
rect 11700 8132 11724 8134
rect 11484 8112 11780 8132
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11336 7880 11388 7886
rect 11532 7857 11560 7958
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11336 7822 11388 7828
rect 11518 7848 11574 7857
rect 11518 7783 11574 7792
rect 11624 7256 11652 7890
rect 11716 7342 11744 7958
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11348 7228 11652 7256
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11164 3738 11192 5782
rect 11256 5710 11284 6394
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11348 5098 11376 7228
rect 11484 7100 11780 7120
rect 11540 7098 11564 7100
rect 11620 7098 11644 7100
rect 11700 7098 11724 7100
rect 11562 7046 11564 7098
rect 11626 7046 11638 7098
rect 11700 7046 11702 7098
rect 11540 7044 11564 7046
rect 11620 7044 11644 7046
rect 11700 7044 11724 7046
rect 11484 7024 11780 7044
rect 11808 6458 11836 9454
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 7410 11928 7686
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11484 6012 11780 6032
rect 11540 6010 11564 6012
rect 11620 6010 11644 6012
rect 11700 6010 11724 6012
rect 11562 5958 11564 6010
rect 11626 5958 11638 6010
rect 11700 5958 11702 6010
rect 11540 5956 11564 5958
rect 11620 5956 11644 5958
rect 11700 5956 11724 5958
rect 11484 5936 11780 5956
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11716 5302 11744 5646
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11808 5166 11836 6394
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 11484 4924 11780 4944
rect 11540 4922 11564 4924
rect 11620 4922 11644 4924
rect 11700 4922 11724 4924
rect 11562 4870 11564 4922
rect 11626 4870 11638 4922
rect 11700 4870 11702 4922
rect 11540 4868 11564 4870
rect 11620 4868 11644 4870
rect 11700 4868 11724 4870
rect 11484 4848 11780 4868
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11532 4078 11560 4422
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 11348 2990 11376 3878
rect 11484 3836 11780 3856
rect 11540 3834 11564 3836
rect 11620 3834 11644 3836
rect 11700 3834 11724 3836
rect 11562 3782 11564 3834
rect 11626 3782 11638 3834
rect 11700 3782 11702 3834
rect 11540 3780 11564 3782
rect 11620 3780 11644 3782
rect 11700 3780 11724 3782
rect 11484 3760 11780 3780
rect 11808 3534 11836 4218
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 8220 480 8248 2246
rect 8852 2204 9148 2224
rect 8908 2202 8932 2204
rect 8988 2202 9012 2204
rect 9068 2202 9092 2204
rect 8930 2150 8932 2202
rect 8994 2150 9006 2202
rect 9068 2150 9070 2202
rect 8908 2148 8932 2150
rect 8988 2148 9012 2150
rect 9068 2148 9092 2150
rect 8852 2128 9148 2148
rect 9784 480 9812 2858
rect 11484 2748 11780 2768
rect 11540 2746 11564 2748
rect 11620 2746 11644 2748
rect 11700 2746 11724 2748
rect 11562 2694 11564 2746
rect 11626 2694 11638 2746
rect 11700 2694 11702 2746
rect 11540 2692 11564 2694
rect 11620 2692 11644 2694
rect 11700 2692 11724 2694
rect 11484 2672 11780 2692
rect 11992 2514 12020 9862
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12084 3670 12112 6122
rect 12176 4554 12204 11766
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12452 10266 12480 11494
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12452 9058 12480 9114
rect 12452 9030 12572 9058
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12452 8090 12480 8910
rect 12544 8906 12572 9030
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12636 8294 12664 10202
rect 12728 10062 12756 10406
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12728 9450 12756 9998
rect 12707 9444 12759 9450
rect 12707 9386 12759 9392
rect 12820 9178 12848 11494
rect 12912 10810 12940 11494
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 13004 10810 13032 11154
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13004 10690 13032 10746
rect 12912 10662 13032 10690
rect 12912 9382 12940 10662
rect 13096 10266 13124 13223
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13082 9480 13138 9489
rect 13082 9415 13138 9424
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12912 8566 12940 9318
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 8090 12848 8230
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 7546 12296 7686
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12348 7472 12400 7478
rect 12400 7420 12480 7426
rect 12348 7414 12480 7420
rect 12360 7398 12480 7414
rect 12348 7336 12400 7342
rect 12346 7304 12348 7313
rect 12400 7304 12402 7313
rect 12346 7239 12402 7248
rect 12452 6322 12480 7398
rect 12544 7274 12572 7754
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12360 5778 12388 6190
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 12452 2990 12480 6054
rect 12544 5846 12572 6598
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12544 5234 12572 5782
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12636 5030 12664 7958
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12716 7336 12768 7342
rect 12820 7324 12848 7822
rect 12768 7296 12848 7324
rect 12912 7313 12940 8502
rect 13096 8362 13124 9415
rect 13188 8974 13216 15807
rect 14554 15464 14610 15473
rect 14554 15399 14610 15408
rect 13818 14648 13874 14657
rect 13818 14583 13874 14592
rect 13832 12442 13860 14583
rect 14116 14172 14412 14192
rect 14172 14170 14196 14172
rect 14252 14170 14276 14172
rect 14332 14170 14356 14172
rect 14194 14118 14196 14170
rect 14258 14118 14270 14170
rect 14332 14118 14334 14170
rect 14172 14116 14196 14118
rect 14252 14116 14276 14118
rect 14332 14116 14356 14118
rect 14116 14096 14412 14116
rect 13910 13968 13966 13977
rect 13910 13903 13966 13912
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13280 10470 13308 10950
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13372 10266 13400 10610
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13266 9208 13322 9217
rect 13372 9178 13400 9998
rect 13266 9143 13322 9152
rect 13360 9172 13412 9178
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13280 8838 13308 9143
rect 13360 9114 13412 9120
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13372 8634 13400 8978
rect 13464 8838 13492 11698
rect 13924 11506 13952 13903
rect 14116 13084 14412 13104
rect 14172 13082 14196 13084
rect 14252 13082 14276 13084
rect 14332 13082 14356 13084
rect 14194 13030 14196 13082
rect 14258 13030 14270 13082
rect 14332 13030 14334 13082
rect 14172 13028 14196 13030
rect 14252 13028 14276 13030
rect 14332 13028 14356 13030
rect 14116 13008 14412 13028
rect 14462 12880 14518 12889
rect 14462 12815 14518 12824
rect 14116 11996 14412 12016
rect 14172 11994 14196 11996
rect 14252 11994 14276 11996
rect 14332 11994 14356 11996
rect 14194 11942 14196 11994
rect 14258 11942 14270 11994
rect 14332 11942 14334 11994
rect 14172 11940 14196 11942
rect 14252 11940 14276 11942
rect 14332 11940 14356 11942
rect 14116 11920 14412 11940
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 13832 11478 13952 11506
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 10674 13584 11154
rect 13832 10690 13860 11478
rect 14292 11354 14320 11698
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 14016 10742 14044 11222
rect 14116 10908 14412 10928
rect 14172 10906 14196 10908
rect 14252 10906 14276 10908
rect 14332 10906 14356 10908
rect 14194 10854 14196 10906
rect 14258 10854 14270 10906
rect 14332 10854 14334 10906
rect 14172 10852 14196 10854
rect 14252 10852 14276 10854
rect 14332 10852 14356 10854
rect 14116 10832 14412 10852
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13740 10662 13860 10690
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 13556 8974 13584 10610
rect 13740 10198 13768 10662
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13648 9625 13676 9930
rect 13634 9616 13690 9625
rect 13634 9551 13690 9560
rect 13832 9518 13860 10474
rect 13910 10432 13966 10441
rect 13910 10367 13966 10376
rect 13924 9926 13952 10367
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12716 7278 12768 7284
rect 12820 6798 12848 7296
rect 12898 7304 12954 7313
rect 12898 7239 12954 7248
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5914 12848 6054
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12820 4758 12848 5306
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12912 3942 12940 6938
rect 13004 5166 13032 7822
rect 13096 5370 13124 8298
rect 13174 7848 13230 7857
rect 13174 7783 13230 7792
rect 13188 7342 13216 7783
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 7002 13216 7142
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13188 5234 13216 5510
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3058 12940 3878
rect 13004 3466 13032 5102
rect 13096 4622 13124 5170
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13096 4214 13124 4558
rect 13188 4282 13216 5170
rect 13280 4758 13308 8434
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 13280 3602 13308 4694
rect 13372 4214 13400 8366
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13648 4010 13676 9386
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 8362 13768 9318
rect 14016 8906 14044 10066
rect 14116 9820 14412 9840
rect 14172 9818 14196 9820
rect 14252 9818 14276 9820
rect 14332 9818 14356 9820
rect 14194 9766 14196 9818
rect 14258 9766 14270 9818
rect 14332 9766 14334 9818
rect 14172 9764 14196 9766
rect 14252 9764 14276 9766
rect 14332 9764 14356 9766
rect 14116 9744 14412 9764
rect 14476 9586 14504 12815
rect 14568 11830 14596 15399
rect 14936 15230 14964 16623
rect 16394 16280 16450 16289
rect 16394 16215 16450 16224
rect 14924 15224 14976 15230
rect 14924 15166 14976 15172
rect 16118 13832 16174 13841
rect 16118 13767 16174 13776
rect 15014 12472 15070 12481
rect 15014 12407 15070 12416
rect 14832 12096 14884 12102
rect 14830 12064 14832 12073
rect 14884 12064 14886 12073
rect 14830 11999 14886 12008
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 15028 11642 15056 12407
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15106 12064 15162 12073
rect 15106 11999 15162 12008
rect 14752 11614 15056 11642
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13832 8430 13860 8842
rect 14116 8732 14412 8752
rect 14172 8730 14196 8732
rect 14252 8730 14276 8732
rect 14332 8730 14356 8732
rect 14194 8678 14196 8730
rect 14258 8678 14270 8730
rect 14332 8678 14334 8730
rect 14172 8676 14196 8678
rect 14252 8676 14276 8678
rect 14332 8676 14356 8678
rect 14116 8656 14412 8676
rect 14094 8528 14150 8537
rect 14094 8463 14150 8472
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13740 7818 13768 8298
rect 14108 8090 14136 8463
rect 14476 8090 14504 8978
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14568 7970 14596 10406
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14660 9625 14688 9658
rect 14646 9616 14702 9625
rect 14646 9551 14702 9560
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14476 7942 14596 7970
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13740 7410 13768 7754
rect 14116 7644 14412 7664
rect 14172 7642 14196 7644
rect 14252 7642 14276 7644
rect 14332 7642 14356 7644
rect 14194 7590 14196 7642
rect 14258 7590 14270 7642
rect 14332 7590 14334 7642
rect 14172 7588 14196 7590
rect 14252 7588 14276 7590
rect 14332 7588 14356 7590
rect 14116 7568 14412 7588
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13832 5778 13860 6870
rect 13924 6254 13952 7482
rect 14370 7304 14426 7313
rect 14370 7239 14372 7248
rect 14424 7239 14426 7248
rect 14372 7210 14424 7216
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14292 6866 14320 7142
rect 14384 6934 14412 7210
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14476 6866 14504 7942
rect 14556 7880 14608 7886
rect 14660 7857 14688 8774
rect 14752 8022 14780 11614
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14830 11248 14886 11257
rect 14830 11183 14886 11192
rect 14844 9586 14872 11183
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14844 8265 14872 9318
rect 14936 9178 14964 11494
rect 15014 10840 15070 10849
rect 15014 10775 15070 10784
rect 15028 9654 15056 10775
rect 15120 10690 15148 11999
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 11354 15424 11494
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15580 10810 15608 11698
rect 15672 11626 15700 12174
rect 15844 11688 15896 11694
rect 15750 11656 15806 11665
rect 15660 11620 15712 11626
rect 15844 11630 15896 11636
rect 15750 11591 15806 11600
rect 15660 11562 15712 11568
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15120 10662 15516 10690
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15120 8650 15148 10134
rect 15212 9586 15240 10474
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15212 9110 15240 9522
rect 15304 9217 15332 10134
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15396 9654 15424 10066
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15384 9444 15436 9450
rect 15384 9386 15436 9392
rect 15396 9353 15424 9386
rect 15382 9344 15438 9353
rect 15382 9279 15438 9288
rect 15290 9208 15346 9217
rect 15290 9143 15346 9152
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15028 8622 15148 8650
rect 14830 8256 14886 8265
rect 14830 8191 14886 8200
rect 14740 8016 14792 8022
rect 14740 7958 14792 7964
rect 14832 8016 14884 8022
rect 14832 7958 14884 7964
rect 14556 7822 14608 7828
rect 14646 7848 14702 7857
rect 14568 7002 14596 7822
rect 14646 7783 14702 7792
rect 14646 7440 14702 7449
rect 14646 7375 14702 7384
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14660 6730 14688 7375
rect 14844 7206 14872 7958
rect 15028 7274 15056 8622
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15016 7268 15068 7274
rect 15016 7210 15068 7216
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14116 6556 14412 6576
rect 14172 6554 14196 6556
rect 14252 6554 14276 6556
rect 14332 6554 14356 6556
rect 14194 6502 14196 6554
rect 14258 6502 14270 6554
rect 14332 6502 14334 6554
rect 14172 6500 14196 6502
rect 14252 6500 14276 6502
rect 14332 6500 14356 6502
rect 14116 6480 14412 6500
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 14188 6248 14240 6254
rect 15028 6236 15056 7210
rect 14188 6190 14240 6196
rect 14936 6208 15056 6236
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13924 5710 13952 6190
rect 14200 6118 14228 6190
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 14116 5468 14412 5488
rect 14172 5466 14196 5468
rect 14252 5466 14276 5468
rect 14332 5466 14356 5468
rect 14194 5414 14196 5466
rect 14258 5414 14270 5466
rect 14332 5414 14334 5466
rect 14172 5412 14196 5414
rect 14252 5412 14276 5414
rect 14332 5412 14356 5414
rect 14116 5392 14412 5412
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 12992 3460 13044 3466
rect 12992 3402 13044 3408
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 13004 2990 13032 3402
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 13280 2922 13308 3538
rect 13740 3126 13768 4966
rect 14108 4826 14136 4966
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14116 4380 14412 4400
rect 14172 4378 14196 4380
rect 14252 4378 14276 4380
rect 14332 4378 14356 4380
rect 14194 4326 14196 4378
rect 14258 4326 14270 4378
rect 14332 4326 14334 4378
rect 14172 4324 14196 4326
rect 14252 4324 14276 4326
rect 14332 4324 14356 4326
rect 14116 4304 14412 4324
rect 14936 4078 14964 6208
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15028 4146 15056 6054
rect 15120 5681 15148 8502
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15212 5846 15240 7686
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 5914 15332 6598
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15106 5672 15162 5681
rect 15106 5607 15162 5616
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 15396 4010 15424 9279
rect 15488 8022 15516 10662
rect 15580 10062 15608 10746
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15566 9208 15622 9217
rect 15566 9143 15622 9152
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 14116 3292 14412 3312
rect 14172 3290 14196 3292
rect 14252 3290 14276 3292
rect 14332 3290 14356 3292
rect 14194 3238 14196 3290
rect 14258 3238 14270 3290
rect 14332 3238 14334 3290
rect 14172 3236 14196 3238
rect 14252 3236 14276 3238
rect 14332 3236 14356 3238
rect 14116 3216 14412 3236
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11256 480 11284 2382
rect 12728 480 12756 2858
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14016 1442 14044 2790
rect 14116 2204 14412 2224
rect 14172 2202 14196 2204
rect 14252 2202 14276 2204
rect 14332 2202 14356 2204
rect 14194 2150 14196 2202
rect 14258 2150 14270 2202
rect 14332 2150 14334 2202
rect 14172 2148 14196 2150
rect 14252 2148 14276 2150
rect 14332 2148 14356 2150
rect 14116 2128 14412 2148
rect 14016 1414 14320 1442
rect 14292 480 14320 1414
rect 14568 649 14596 3878
rect 15120 3641 15148 3878
rect 15106 3632 15162 3641
rect 15580 3602 15608 9143
rect 15672 5166 15700 11562
rect 15764 11354 15792 11591
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15764 9178 15792 9862
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15856 8430 15884 11630
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15948 10062 15976 11086
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15948 9586 15976 9998
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 16040 9897 16068 9930
rect 16026 9888 16082 9897
rect 16026 9823 16082 9832
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15948 9081 15976 9318
rect 15934 9072 15990 9081
rect 15934 9007 15990 9016
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 16132 8362 16160 13767
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15856 7886 15884 8230
rect 16132 8090 16160 8298
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15856 6798 15884 7822
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 16040 6497 16068 7142
rect 16118 7032 16174 7041
rect 16118 6967 16174 6976
rect 16026 6488 16082 6497
rect 16132 6458 16160 6967
rect 16026 6423 16082 6432
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16224 6089 16252 12038
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16210 6080 16266 6089
rect 16210 6015 16266 6024
rect 15844 5636 15896 5642
rect 15844 5578 15896 5584
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15106 3567 15162 3576
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14660 1465 14688 3334
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 1873 14872 2246
rect 14830 1864 14886 1873
rect 14830 1799 14886 1808
rect 14646 1456 14702 1465
rect 14646 1391 14702 1400
rect 14554 640 14610 649
rect 14554 575 14610 584
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 3698 0 3754 480
rect 5262 0 5318 480
rect 6734 0 6790 480
rect 8206 0 8262 480
rect 9770 0 9826 480
rect 11242 0 11298 480
rect 12714 0 12770 480
rect 14278 0 14334 480
rect 14936 241 14964 2790
rect 15120 1057 15148 2790
rect 15106 1048 15162 1057
rect 15106 983 15162 992
rect 15764 480 15792 4082
rect 15856 2514 15884 5578
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 16040 5273 16068 5510
rect 16026 5264 16082 5273
rect 16026 5199 16082 5208
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16040 4865 16068 4966
rect 16026 4856 16082 4865
rect 16026 4791 16082 4800
rect 16028 4480 16080 4486
rect 16026 4448 16028 4457
rect 16080 4448 16082 4457
rect 16026 4383 16082 4392
rect 16026 4040 16082 4049
rect 16026 3975 16082 3984
rect 16040 3942 16068 3975
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16316 3602 16344 11154
rect 16408 9722 16436 16215
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16040 3097 16068 3334
rect 16026 3088 16082 3097
rect 16026 3023 16082 3032
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 16040 2689 16068 2790
rect 16026 2680 16082 2689
rect 16026 2615 16082 2624
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 16028 2304 16080 2310
rect 16026 2272 16028 2281
rect 16080 2272 16082 2281
rect 16026 2207 16082 2216
rect 17236 480 17264 7754
rect 14922 232 14978 241
rect 14922 167 14978 176
rect 15750 0 15806 480
rect 17222 0 17278 480
<< via2 >>
rect 4802 16632 4858 16688
rect 14922 16632 14978 16688
rect 3054 16224 3110 16280
rect 2318 14184 2374 14240
rect 2962 13776 3018 13832
rect 2318 11736 2374 11792
rect 2870 11600 2926 11656
rect 2410 9016 2466 9072
rect 1582 5616 1638 5672
rect 1582 3576 1638 3632
rect 2134 1400 2190 1456
rect 2502 8916 2504 8936
rect 2504 8916 2556 8936
rect 2556 8916 2558 8936
rect 2502 8880 2558 8916
rect 2686 10512 2742 10568
rect 2962 10240 3018 10296
rect 3146 15816 3202 15872
rect 3882 15408 3938 15464
rect 3514 15000 3570 15056
rect 3588 14170 3644 14172
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3588 14118 3614 14170
rect 3614 14118 3644 14170
rect 3668 14118 3678 14170
rect 3678 14118 3724 14170
rect 3748 14118 3794 14170
rect 3794 14118 3804 14170
rect 3828 14118 3858 14170
rect 3858 14118 3884 14170
rect 3588 14116 3644 14118
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 4158 13232 4214 13288
rect 3588 13082 3644 13084
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3588 13030 3614 13082
rect 3614 13030 3644 13082
rect 3668 13030 3678 13082
rect 3678 13030 3724 13082
rect 3748 13030 3794 13082
rect 3794 13030 3804 13082
rect 3828 13030 3858 13082
rect 3858 13030 3884 13082
rect 3588 13028 3644 13030
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3514 12824 3570 12880
rect 4066 12416 4122 12472
rect 3146 10784 3202 10840
rect 2870 9832 2926 9888
rect 2778 8472 2834 8528
rect 2962 6432 3018 6488
rect 2870 4800 2926 4856
rect 2778 4392 2834 4448
rect 2870 2252 2872 2272
rect 2872 2252 2924 2272
rect 2924 2252 2926 2272
rect 2870 2216 2926 2252
rect 2962 1808 3018 1864
rect 3054 992 3110 1048
rect 3422 12008 3478 12064
rect 3588 11994 3644 11996
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3588 11942 3614 11994
rect 3614 11942 3644 11994
rect 3668 11942 3678 11994
rect 3678 11942 3724 11994
rect 3748 11942 3794 11994
rect 3794 11942 3804 11994
rect 3828 11942 3858 11994
rect 3858 11942 3884 11994
rect 3588 11940 3644 11942
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 4158 12144 4214 12200
rect 3330 10240 3386 10296
rect 3588 10906 3644 10908
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3588 10854 3614 10906
rect 3614 10854 3644 10906
rect 3668 10854 3678 10906
rect 3678 10854 3724 10906
rect 3748 10854 3794 10906
rect 3794 10854 3804 10906
rect 3828 10854 3858 10906
rect 3858 10854 3884 10906
rect 3588 10852 3644 10854
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3588 9818 3644 9820
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3588 9766 3614 9818
rect 3614 9766 3644 9818
rect 3668 9766 3678 9818
rect 3678 9766 3724 9818
rect 3748 9766 3794 9818
rect 3794 9766 3804 9818
rect 3828 9766 3858 9818
rect 3858 9766 3884 9818
rect 3588 9764 3644 9766
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3514 9560 3570 9616
rect 4066 11192 4122 11248
rect 13174 15816 13230 15872
rect 6220 14714 6276 14716
rect 6300 14714 6356 14716
rect 6380 14714 6436 14716
rect 6460 14714 6516 14716
rect 6220 14662 6246 14714
rect 6246 14662 6276 14714
rect 6300 14662 6310 14714
rect 6310 14662 6356 14714
rect 6380 14662 6426 14714
rect 6426 14662 6436 14714
rect 6460 14662 6490 14714
rect 6490 14662 6516 14714
rect 6220 14660 6276 14662
rect 6300 14660 6356 14662
rect 6380 14660 6436 14662
rect 6460 14660 6516 14662
rect 5814 14592 5870 14648
rect 4986 11228 4988 11248
rect 4988 11228 5040 11248
rect 5040 11228 5042 11248
rect 4986 11192 5042 11228
rect 4066 10376 4122 10432
rect 3588 8730 3644 8732
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3588 8678 3614 8730
rect 3614 8678 3644 8730
rect 3668 8678 3678 8730
rect 3678 8678 3724 8730
rect 3748 8678 3794 8730
rect 3794 8678 3804 8730
rect 3828 8678 3858 8730
rect 3858 8678 3884 8730
rect 3588 8676 3644 8678
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3974 7792 4030 7848
rect 3588 7642 3644 7644
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3588 7590 3614 7642
rect 3614 7590 3644 7642
rect 3668 7590 3678 7642
rect 3678 7590 3724 7642
rect 3748 7590 3794 7642
rect 3794 7590 3804 7642
rect 3828 7590 3858 7642
rect 3858 7590 3884 7642
rect 3588 7588 3644 7590
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 4066 7384 4122 7440
rect 3422 6160 3478 6216
rect 3422 3032 3478 3088
rect 3588 6554 3644 6556
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3588 6502 3614 6554
rect 3614 6502 3644 6554
rect 3668 6502 3678 6554
rect 3678 6502 3724 6554
rect 3748 6502 3794 6554
rect 3794 6502 3804 6554
rect 3828 6502 3858 6554
rect 3858 6502 3884 6554
rect 3588 6500 3644 6502
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3588 5466 3644 5468
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3588 5414 3614 5466
rect 3614 5414 3644 5466
rect 3668 5414 3678 5466
rect 3678 5414 3724 5466
rect 3748 5414 3794 5466
rect 3794 5414 3804 5466
rect 3828 5414 3858 5466
rect 3858 5414 3884 5466
rect 3588 5412 3644 5414
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3588 4378 3644 4380
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3588 4326 3614 4378
rect 3614 4326 3644 4378
rect 3668 4326 3678 4378
rect 3678 4326 3724 4378
rect 3748 4326 3794 4378
rect 3794 4326 3804 4378
rect 3828 4326 3858 4378
rect 3858 4326 3884 4378
rect 3588 4324 3644 4326
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 4526 8880 4582 8936
rect 4066 7112 4122 7168
rect 4066 5208 4122 5264
rect 4710 9560 4766 9616
rect 6220 13626 6276 13628
rect 6300 13626 6356 13628
rect 6380 13626 6436 13628
rect 6460 13626 6516 13628
rect 6220 13574 6246 13626
rect 6246 13574 6276 13626
rect 6300 13574 6310 13626
rect 6310 13574 6356 13626
rect 6380 13574 6426 13626
rect 6426 13574 6436 13626
rect 6460 13574 6490 13626
rect 6490 13574 6516 13626
rect 6220 13572 6276 13574
rect 6300 13572 6356 13574
rect 6380 13572 6436 13574
rect 6460 13572 6516 13574
rect 6220 12538 6276 12540
rect 6300 12538 6356 12540
rect 6380 12538 6436 12540
rect 6460 12538 6516 12540
rect 6220 12486 6246 12538
rect 6246 12486 6276 12538
rect 6300 12486 6310 12538
rect 6310 12486 6356 12538
rect 6380 12486 6426 12538
rect 6426 12486 6436 12538
rect 6460 12486 6490 12538
rect 6490 12486 6516 12538
rect 6220 12484 6276 12486
rect 6300 12484 6356 12486
rect 6380 12484 6436 12486
rect 6460 12484 6516 12486
rect 4066 3984 4122 4040
rect 3588 3290 3644 3292
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3588 3238 3614 3290
rect 3614 3238 3644 3290
rect 3668 3238 3678 3290
rect 3678 3238 3724 3290
rect 3748 3238 3794 3290
rect 3794 3238 3804 3290
rect 3828 3238 3858 3290
rect 3858 3238 3884 3290
rect 3588 3236 3644 3238
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3330 2624 3386 2680
rect 3588 2202 3644 2204
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3588 2150 3614 2202
rect 3614 2150 3644 2202
rect 3668 2150 3678 2202
rect 3678 2150 3724 2202
rect 3748 2150 3794 2202
rect 3794 2150 3804 2202
rect 3828 2150 3858 2202
rect 3858 2150 3884 2202
rect 3588 2148 3644 2150
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 6220 11450 6276 11452
rect 6300 11450 6356 11452
rect 6380 11450 6436 11452
rect 6460 11450 6516 11452
rect 6220 11398 6246 11450
rect 6246 11398 6276 11450
rect 6300 11398 6310 11450
rect 6310 11398 6356 11450
rect 6380 11398 6426 11450
rect 6426 11398 6436 11450
rect 6460 11398 6490 11450
rect 6490 11398 6516 11450
rect 6220 11396 6276 11398
rect 6300 11396 6356 11398
rect 6380 11396 6436 11398
rect 6460 11396 6516 11398
rect 6220 10362 6276 10364
rect 6300 10362 6356 10364
rect 6380 10362 6436 10364
rect 6460 10362 6516 10364
rect 6220 10310 6246 10362
rect 6246 10310 6276 10362
rect 6300 10310 6310 10362
rect 6310 10310 6356 10362
rect 6380 10310 6426 10362
rect 6426 10310 6436 10362
rect 6460 10310 6490 10362
rect 6490 10310 6516 10362
rect 6220 10308 6276 10310
rect 6300 10308 6356 10310
rect 6380 10308 6436 10310
rect 6460 10308 6516 10310
rect 6220 9274 6276 9276
rect 6300 9274 6356 9276
rect 6380 9274 6436 9276
rect 6460 9274 6516 9276
rect 6220 9222 6246 9274
rect 6246 9222 6276 9274
rect 6300 9222 6310 9274
rect 6310 9222 6356 9274
rect 6380 9222 6426 9274
rect 6426 9222 6436 9274
rect 6460 9222 6490 9274
rect 6490 9222 6516 9274
rect 6220 9220 6276 9222
rect 6300 9220 6356 9222
rect 6380 9220 6436 9222
rect 6460 9220 6516 9222
rect 6220 8186 6276 8188
rect 6300 8186 6356 8188
rect 6380 8186 6436 8188
rect 6460 8186 6516 8188
rect 6220 8134 6246 8186
rect 6246 8134 6276 8186
rect 6300 8134 6310 8186
rect 6310 8134 6356 8186
rect 6380 8134 6426 8186
rect 6426 8134 6436 8186
rect 6460 8134 6490 8186
rect 6490 8134 6516 8186
rect 6220 8132 6276 8134
rect 6300 8132 6356 8134
rect 6380 8132 6436 8134
rect 6460 8132 6516 8134
rect 6220 7098 6276 7100
rect 6300 7098 6356 7100
rect 6380 7098 6436 7100
rect 6460 7098 6516 7100
rect 6220 7046 6246 7098
rect 6246 7046 6276 7098
rect 6300 7046 6310 7098
rect 6310 7046 6356 7098
rect 6380 7046 6426 7098
rect 6426 7046 6436 7098
rect 6460 7046 6490 7098
rect 6490 7046 6516 7098
rect 6220 7044 6276 7046
rect 6300 7044 6356 7046
rect 6380 7044 6436 7046
rect 6460 7044 6516 7046
rect 10598 15000 10654 15056
rect 8852 14170 8908 14172
rect 8932 14170 8988 14172
rect 9012 14170 9068 14172
rect 9092 14170 9148 14172
rect 8852 14118 8878 14170
rect 8878 14118 8908 14170
rect 8932 14118 8942 14170
rect 8942 14118 8988 14170
rect 9012 14118 9058 14170
rect 9058 14118 9068 14170
rect 9092 14118 9122 14170
rect 9122 14118 9148 14170
rect 8852 14116 8908 14118
rect 8932 14116 8988 14118
rect 9012 14116 9068 14118
rect 9092 14116 9148 14118
rect 8852 13082 8908 13084
rect 8932 13082 8988 13084
rect 9012 13082 9068 13084
rect 9092 13082 9148 13084
rect 8852 13030 8878 13082
rect 8878 13030 8908 13082
rect 8932 13030 8942 13082
rect 8942 13030 8988 13082
rect 9012 13030 9058 13082
rect 9058 13030 9068 13082
rect 9092 13030 9122 13082
rect 9122 13030 9148 13082
rect 8852 13028 8908 13030
rect 8932 13028 8988 13030
rect 9012 13028 9068 13030
rect 9092 13028 9148 13030
rect 7378 8880 7434 8936
rect 6220 6010 6276 6012
rect 6300 6010 6356 6012
rect 6380 6010 6436 6012
rect 6460 6010 6516 6012
rect 6220 5958 6246 6010
rect 6246 5958 6276 6010
rect 6300 5958 6310 6010
rect 6310 5958 6356 6010
rect 6380 5958 6426 6010
rect 6426 5958 6436 6010
rect 6460 5958 6490 6010
rect 6490 5958 6516 6010
rect 6220 5956 6276 5958
rect 6300 5956 6356 5958
rect 6380 5956 6436 5958
rect 6460 5956 6516 5958
rect 6220 4922 6276 4924
rect 6300 4922 6356 4924
rect 6380 4922 6436 4924
rect 6460 4922 6516 4924
rect 6220 4870 6246 4922
rect 6246 4870 6276 4922
rect 6300 4870 6310 4922
rect 6310 4870 6356 4922
rect 6380 4870 6426 4922
rect 6426 4870 6436 4922
rect 6460 4870 6490 4922
rect 6490 4870 6516 4922
rect 6220 4868 6276 4870
rect 6300 4868 6356 4870
rect 6380 4868 6436 4870
rect 6460 4868 6516 4870
rect 6220 3834 6276 3836
rect 6300 3834 6356 3836
rect 6380 3834 6436 3836
rect 6460 3834 6516 3836
rect 6220 3782 6246 3834
rect 6246 3782 6276 3834
rect 6300 3782 6310 3834
rect 6310 3782 6356 3834
rect 6380 3782 6426 3834
rect 6426 3782 6436 3834
rect 6460 3782 6490 3834
rect 6490 3782 6516 3834
rect 6220 3780 6276 3782
rect 6300 3780 6356 3782
rect 6380 3780 6436 3782
rect 6460 3780 6516 3782
rect 7838 11464 7894 11520
rect 7746 9052 7748 9072
rect 7748 9052 7800 9072
rect 7800 9052 7802 9072
rect 7746 9016 7802 9052
rect 8206 12180 8208 12200
rect 8208 12180 8260 12200
rect 8260 12180 8262 12200
rect 8206 12144 8262 12180
rect 8852 11994 8908 11996
rect 8932 11994 8988 11996
rect 9012 11994 9068 11996
rect 9092 11994 9148 11996
rect 8852 11942 8878 11994
rect 8878 11942 8908 11994
rect 8932 11942 8942 11994
rect 8942 11942 8988 11994
rect 9012 11942 9058 11994
rect 9058 11942 9068 11994
rect 9092 11942 9122 11994
rect 9122 11942 9148 11994
rect 8852 11940 8908 11942
rect 8932 11940 8988 11942
rect 9012 11940 9068 11942
rect 9092 11940 9148 11942
rect 8022 11464 8078 11520
rect 8298 11212 8354 11248
rect 8298 11192 8300 11212
rect 8300 11192 8352 11212
rect 8352 11192 8354 11212
rect 9402 11736 9458 11792
rect 8852 10906 8908 10908
rect 8932 10906 8988 10908
rect 9012 10906 9068 10908
rect 9092 10906 9148 10908
rect 8852 10854 8878 10906
rect 8878 10854 8908 10906
rect 8932 10854 8942 10906
rect 8942 10854 8988 10906
rect 9012 10854 9058 10906
rect 9058 10854 9068 10906
rect 9092 10854 9122 10906
rect 9122 10854 9148 10906
rect 8852 10852 8908 10854
rect 8932 10852 8988 10854
rect 9012 10852 9068 10854
rect 9092 10852 9148 10854
rect 9218 10548 9220 10568
rect 9220 10548 9272 10568
rect 9272 10548 9274 10568
rect 9218 10512 9274 10548
rect 8574 9424 8630 9480
rect 8298 8472 8354 8528
rect 3146 584 3202 640
rect 6220 2746 6276 2748
rect 6300 2746 6356 2748
rect 6380 2746 6436 2748
rect 6460 2746 6516 2748
rect 6220 2694 6246 2746
rect 6246 2694 6276 2746
rect 6300 2694 6310 2746
rect 6310 2694 6356 2746
rect 6380 2694 6426 2746
rect 6426 2694 6436 2746
rect 6460 2694 6490 2746
rect 6490 2694 6516 2746
rect 6220 2692 6276 2694
rect 6300 2692 6356 2694
rect 6380 2692 6436 2694
rect 6460 2692 6516 2694
rect 8206 6704 8262 6760
rect 8852 9818 8908 9820
rect 8932 9818 8988 9820
rect 9012 9818 9068 9820
rect 9092 9818 9148 9820
rect 8852 9766 8878 9818
rect 8878 9766 8908 9818
rect 8932 9766 8942 9818
rect 8942 9766 8988 9818
rect 9012 9766 9058 9818
rect 9058 9766 9068 9818
rect 9092 9766 9122 9818
rect 9122 9766 9148 9818
rect 8852 9764 8908 9766
rect 8932 9764 8988 9766
rect 9012 9764 9068 9766
rect 9092 9764 9148 9766
rect 9126 9424 9182 9480
rect 11484 14714 11540 14716
rect 11564 14714 11620 14716
rect 11644 14714 11700 14716
rect 11724 14714 11780 14716
rect 11484 14662 11510 14714
rect 11510 14662 11540 14714
rect 11564 14662 11574 14714
rect 11574 14662 11620 14714
rect 11644 14662 11690 14714
rect 11690 14662 11700 14714
rect 11724 14662 11754 14714
rect 11754 14662 11780 14714
rect 11484 14660 11540 14662
rect 11564 14660 11620 14662
rect 11644 14660 11700 14662
rect 11724 14660 11780 14662
rect 11484 13626 11540 13628
rect 11564 13626 11620 13628
rect 11644 13626 11700 13628
rect 11724 13626 11780 13628
rect 11484 13574 11510 13626
rect 11510 13574 11540 13626
rect 11564 13574 11574 13626
rect 11574 13574 11620 13626
rect 11644 13574 11690 13626
rect 11690 13574 11700 13626
rect 11724 13574 11754 13626
rect 11754 13574 11780 13626
rect 11484 13572 11540 13574
rect 11564 13572 11620 13574
rect 11644 13572 11700 13574
rect 11724 13572 11780 13574
rect 10322 9696 10378 9752
rect 8852 8730 8908 8732
rect 8932 8730 8988 8732
rect 9012 8730 9068 8732
rect 9092 8730 9148 8732
rect 8852 8678 8878 8730
rect 8878 8678 8908 8730
rect 8932 8678 8942 8730
rect 8942 8678 8988 8730
rect 9012 8678 9058 8730
rect 9058 8678 9068 8730
rect 9092 8678 9122 8730
rect 9122 8678 9148 8730
rect 8852 8676 8908 8678
rect 8932 8676 8988 8678
rect 9012 8676 9068 8678
rect 9092 8676 9148 8678
rect 8852 7642 8908 7644
rect 8932 7642 8988 7644
rect 9012 7642 9068 7644
rect 9092 7642 9148 7644
rect 8852 7590 8878 7642
rect 8878 7590 8908 7642
rect 8932 7590 8942 7642
rect 8942 7590 8988 7642
rect 9012 7590 9058 7642
rect 9058 7590 9068 7642
rect 9092 7590 9122 7642
rect 9122 7590 9148 7642
rect 8852 7588 8908 7590
rect 8932 7588 8988 7590
rect 9012 7588 9068 7590
rect 9092 7588 9148 7590
rect 9862 8508 9864 8528
rect 9864 8508 9916 8528
rect 9916 8508 9918 8528
rect 9862 8472 9918 8508
rect 8852 6554 8908 6556
rect 8932 6554 8988 6556
rect 9012 6554 9068 6556
rect 9092 6554 9148 6556
rect 8852 6502 8878 6554
rect 8878 6502 8908 6554
rect 8932 6502 8942 6554
rect 8942 6502 8988 6554
rect 9012 6502 9058 6554
rect 9058 6502 9068 6554
rect 9092 6502 9122 6554
rect 9122 6502 9148 6554
rect 8852 6500 8908 6502
rect 8932 6500 8988 6502
rect 9012 6500 9068 6502
rect 9092 6500 9148 6502
rect 8852 5466 8908 5468
rect 8932 5466 8988 5468
rect 9012 5466 9068 5468
rect 9092 5466 9148 5468
rect 8852 5414 8878 5466
rect 8878 5414 8908 5466
rect 8932 5414 8942 5466
rect 8942 5414 8988 5466
rect 9012 5414 9058 5466
rect 9058 5414 9068 5466
rect 9092 5414 9122 5466
rect 9122 5414 9148 5466
rect 8852 5412 8908 5414
rect 8932 5412 8988 5414
rect 9012 5412 9068 5414
rect 9092 5412 9148 5414
rect 8852 4378 8908 4380
rect 8932 4378 8988 4380
rect 9012 4378 9068 4380
rect 9092 4378 9148 4380
rect 8852 4326 8878 4378
rect 8878 4326 8908 4378
rect 8932 4326 8942 4378
rect 8942 4326 8988 4378
rect 9012 4326 9058 4378
rect 9058 4326 9068 4378
rect 9092 4326 9122 4378
rect 9122 4326 9148 4378
rect 8852 4324 8908 4326
rect 8932 4324 8988 4326
rect 9012 4324 9068 4326
rect 9092 4324 9148 4326
rect 8852 3290 8908 3292
rect 8932 3290 8988 3292
rect 9012 3290 9068 3292
rect 9092 3290 9148 3292
rect 8852 3238 8878 3290
rect 8878 3238 8908 3290
rect 8932 3238 8942 3290
rect 8942 3238 8988 3290
rect 9012 3238 9058 3290
rect 9058 3238 9068 3290
rect 9092 3238 9122 3290
rect 9122 3238 9148 3290
rect 8852 3236 8908 3238
rect 8932 3236 8988 3238
rect 9012 3236 9068 3238
rect 9092 3236 9148 3238
rect 9310 6704 9366 6760
rect 10414 9560 10470 9616
rect 10690 9444 10746 9480
rect 10690 9424 10692 9444
rect 10692 9424 10744 9444
rect 10744 9424 10746 9444
rect 10598 9016 10654 9072
rect 11484 12538 11540 12540
rect 11564 12538 11620 12540
rect 11644 12538 11700 12540
rect 11724 12538 11780 12540
rect 11484 12486 11510 12538
rect 11510 12486 11540 12538
rect 11564 12486 11574 12538
rect 11574 12486 11620 12538
rect 11644 12486 11690 12538
rect 11690 12486 11700 12538
rect 11724 12486 11754 12538
rect 11754 12486 11780 12538
rect 11484 12484 11540 12486
rect 11564 12484 11620 12486
rect 11644 12484 11700 12486
rect 11724 12484 11780 12486
rect 11484 11450 11540 11452
rect 11564 11450 11620 11452
rect 11644 11450 11700 11452
rect 11724 11450 11780 11452
rect 11484 11398 11510 11450
rect 11510 11398 11540 11450
rect 11564 11398 11574 11450
rect 11574 11398 11620 11450
rect 11644 11398 11690 11450
rect 11690 11398 11700 11450
rect 11724 11398 11754 11450
rect 11754 11398 11780 11450
rect 11484 11396 11540 11398
rect 11564 11396 11620 11398
rect 11644 11396 11700 11398
rect 11724 11396 11780 11398
rect 13082 13232 13138 13288
rect 11484 10362 11540 10364
rect 11564 10362 11620 10364
rect 11644 10362 11700 10364
rect 11724 10362 11780 10364
rect 11484 10310 11510 10362
rect 11510 10310 11540 10362
rect 11564 10310 11574 10362
rect 11574 10310 11620 10362
rect 11644 10310 11690 10362
rect 11690 10310 11700 10362
rect 11724 10310 11754 10362
rect 11754 10310 11780 10362
rect 11484 10308 11540 10310
rect 11564 10308 11620 10310
rect 11644 10308 11700 10310
rect 11724 10308 11780 10310
rect 11058 9696 11114 9752
rect 11484 9274 11540 9276
rect 11564 9274 11620 9276
rect 11644 9274 11700 9276
rect 11724 9274 11780 9276
rect 11484 9222 11510 9274
rect 11510 9222 11540 9274
rect 11564 9222 11574 9274
rect 11574 9222 11620 9274
rect 11644 9222 11690 9274
rect 11690 9222 11700 9274
rect 11724 9222 11754 9274
rect 11754 9222 11780 9274
rect 11484 9220 11540 9222
rect 11564 9220 11620 9222
rect 11644 9220 11700 9222
rect 11724 9220 11780 9222
rect 11518 8472 11574 8528
rect 11484 8186 11540 8188
rect 11564 8186 11620 8188
rect 11644 8186 11700 8188
rect 11724 8186 11780 8188
rect 11484 8134 11510 8186
rect 11510 8134 11540 8186
rect 11564 8134 11574 8186
rect 11574 8134 11620 8186
rect 11644 8134 11690 8186
rect 11690 8134 11700 8186
rect 11724 8134 11754 8186
rect 11754 8134 11780 8186
rect 11484 8132 11540 8134
rect 11564 8132 11620 8134
rect 11644 8132 11700 8134
rect 11724 8132 11780 8134
rect 11518 7792 11574 7848
rect 11484 7098 11540 7100
rect 11564 7098 11620 7100
rect 11644 7098 11700 7100
rect 11724 7098 11780 7100
rect 11484 7046 11510 7098
rect 11510 7046 11540 7098
rect 11564 7046 11574 7098
rect 11574 7046 11620 7098
rect 11644 7046 11690 7098
rect 11690 7046 11700 7098
rect 11724 7046 11754 7098
rect 11754 7046 11780 7098
rect 11484 7044 11540 7046
rect 11564 7044 11620 7046
rect 11644 7044 11700 7046
rect 11724 7044 11780 7046
rect 11484 6010 11540 6012
rect 11564 6010 11620 6012
rect 11644 6010 11700 6012
rect 11724 6010 11780 6012
rect 11484 5958 11510 6010
rect 11510 5958 11540 6010
rect 11564 5958 11574 6010
rect 11574 5958 11620 6010
rect 11644 5958 11690 6010
rect 11690 5958 11700 6010
rect 11724 5958 11754 6010
rect 11754 5958 11780 6010
rect 11484 5956 11540 5958
rect 11564 5956 11620 5958
rect 11644 5956 11700 5958
rect 11724 5956 11780 5958
rect 11484 4922 11540 4924
rect 11564 4922 11620 4924
rect 11644 4922 11700 4924
rect 11724 4922 11780 4924
rect 11484 4870 11510 4922
rect 11510 4870 11540 4922
rect 11564 4870 11574 4922
rect 11574 4870 11620 4922
rect 11644 4870 11690 4922
rect 11690 4870 11700 4922
rect 11724 4870 11754 4922
rect 11754 4870 11780 4922
rect 11484 4868 11540 4870
rect 11564 4868 11620 4870
rect 11644 4868 11700 4870
rect 11724 4868 11780 4870
rect 11484 3834 11540 3836
rect 11564 3834 11620 3836
rect 11644 3834 11700 3836
rect 11724 3834 11780 3836
rect 11484 3782 11510 3834
rect 11510 3782 11540 3834
rect 11564 3782 11574 3834
rect 11574 3782 11620 3834
rect 11644 3782 11690 3834
rect 11690 3782 11700 3834
rect 11724 3782 11754 3834
rect 11754 3782 11780 3834
rect 11484 3780 11540 3782
rect 11564 3780 11620 3782
rect 11644 3780 11700 3782
rect 11724 3780 11780 3782
rect 8852 2202 8908 2204
rect 8932 2202 8988 2204
rect 9012 2202 9068 2204
rect 9092 2202 9148 2204
rect 8852 2150 8878 2202
rect 8878 2150 8908 2202
rect 8932 2150 8942 2202
rect 8942 2150 8988 2202
rect 9012 2150 9058 2202
rect 9058 2150 9068 2202
rect 9092 2150 9122 2202
rect 9122 2150 9148 2202
rect 8852 2148 8908 2150
rect 8932 2148 8988 2150
rect 9012 2148 9068 2150
rect 9092 2148 9148 2150
rect 11484 2746 11540 2748
rect 11564 2746 11620 2748
rect 11644 2746 11700 2748
rect 11724 2746 11780 2748
rect 11484 2694 11510 2746
rect 11510 2694 11540 2746
rect 11564 2694 11574 2746
rect 11574 2694 11620 2746
rect 11644 2694 11690 2746
rect 11690 2694 11700 2746
rect 11724 2694 11754 2746
rect 11754 2694 11780 2746
rect 11484 2692 11540 2694
rect 11564 2692 11620 2694
rect 11644 2692 11700 2694
rect 11724 2692 11780 2694
rect 13082 9424 13138 9480
rect 12346 7284 12348 7304
rect 12348 7284 12400 7304
rect 12400 7284 12402 7304
rect 12346 7248 12402 7284
rect 14554 15408 14610 15464
rect 13818 14592 13874 14648
rect 14116 14170 14172 14172
rect 14196 14170 14252 14172
rect 14276 14170 14332 14172
rect 14356 14170 14412 14172
rect 14116 14118 14142 14170
rect 14142 14118 14172 14170
rect 14196 14118 14206 14170
rect 14206 14118 14252 14170
rect 14276 14118 14322 14170
rect 14322 14118 14332 14170
rect 14356 14118 14386 14170
rect 14386 14118 14412 14170
rect 14116 14116 14172 14118
rect 14196 14116 14252 14118
rect 14276 14116 14332 14118
rect 14356 14116 14412 14118
rect 13910 13912 13966 13968
rect 13266 9152 13322 9208
rect 14116 13082 14172 13084
rect 14196 13082 14252 13084
rect 14276 13082 14332 13084
rect 14356 13082 14412 13084
rect 14116 13030 14142 13082
rect 14142 13030 14172 13082
rect 14196 13030 14206 13082
rect 14206 13030 14252 13082
rect 14276 13030 14322 13082
rect 14322 13030 14332 13082
rect 14356 13030 14386 13082
rect 14386 13030 14412 13082
rect 14116 13028 14172 13030
rect 14196 13028 14252 13030
rect 14276 13028 14332 13030
rect 14356 13028 14412 13030
rect 14462 12824 14518 12880
rect 14116 11994 14172 11996
rect 14196 11994 14252 11996
rect 14276 11994 14332 11996
rect 14356 11994 14412 11996
rect 14116 11942 14142 11994
rect 14142 11942 14172 11994
rect 14196 11942 14206 11994
rect 14206 11942 14252 11994
rect 14276 11942 14322 11994
rect 14322 11942 14332 11994
rect 14356 11942 14386 11994
rect 14386 11942 14412 11994
rect 14116 11940 14172 11942
rect 14196 11940 14252 11942
rect 14276 11940 14332 11942
rect 14356 11940 14412 11942
rect 14116 10906 14172 10908
rect 14196 10906 14252 10908
rect 14276 10906 14332 10908
rect 14356 10906 14412 10908
rect 14116 10854 14142 10906
rect 14142 10854 14172 10906
rect 14196 10854 14206 10906
rect 14206 10854 14252 10906
rect 14276 10854 14322 10906
rect 14322 10854 14332 10906
rect 14356 10854 14386 10906
rect 14386 10854 14412 10906
rect 14116 10852 14172 10854
rect 14196 10852 14252 10854
rect 14276 10852 14332 10854
rect 14356 10852 14412 10854
rect 13634 9560 13690 9616
rect 13910 10376 13966 10432
rect 12898 7248 12954 7304
rect 13174 7792 13230 7848
rect 14116 9818 14172 9820
rect 14196 9818 14252 9820
rect 14276 9818 14332 9820
rect 14356 9818 14412 9820
rect 14116 9766 14142 9818
rect 14142 9766 14172 9818
rect 14196 9766 14206 9818
rect 14206 9766 14252 9818
rect 14276 9766 14322 9818
rect 14322 9766 14332 9818
rect 14356 9766 14386 9818
rect 14386 9766 14412 9818
rect 14116 9764 14172 9766
rect 14196 9764 14252 9766
rect 14276 9764 14332 9766
rect 14356 9764 14412 9766
rect 16394 16224 16450 16280
rect 16118 13776 16174 13832
rect 15014 12416 15070 12472
rect 14830 12044 14832 12064
rect 14832 12044 14884 12064
rect 14884 12044 14886 12064
rect 14830 12008 14886 12044
rect 15106 12008 15162 12064
rect 14116 8730 14172 8732
rect 14196 8730 14252 8732
rect 14276 8730 14332 8732
rect 14356 8730 14412 8732
rect 14116 8678 14142 8730
rect 14142 8678 14172 8730
rect 14196 8678 14206 8730
rect 14206 8678 14252 8730
rect 14276 8678 14322 8730
rect 14322 8678 14332 8730
rect 14356 8678 14386 8730
rect 14386 8678 14412 8730
rect 14116 8676 14172 8678
rect 14196 8676 14252 8678
rect 14276 8676 14332 8678
rect 14356 8676 14412 8678
rect 14094 8472 14150 8528
rect 14646 9560 14702 9616
rect 14116 7642 14172 7644
rect 14196 7642 14252 7644
rect 14276 7642 14332 7644
rect 14356 7642 14412 7644
rect 14116 7590 14142 7642
rect 14142 7590 14172 7642
rect 14196 7590 14206 7642
rect 14206 7590 14252 7642
rect 14276 7590 14322 7642
rect 14322 7590 14332 7642
rect 14356 7590 14386 7642
rect 14386 7590 14412 7642
rect 14116 7588 14172 7590
rect 14196 7588 14252 7590
rect 14276 7588 14332 7590
rect 14356 7588 14412 7590
rect 14370 7268 14426 7304
rect 14370 7248 14372 7268
rect 14372 7248 14424 7268
rect 14424 7248 14426 7268
rect 14830 11192 14886 11248
rect 15014 10784 15070 10840
rect 15750 11600 15806 11656
rect 15382 9288 15438 9344
rect 15290 9152 15346 9208
rect 14830 8200 14886 8256
rect 14646 7792 14702 7848
rect 14646 7384 14702 7440
rect 14116 6554 14172 6556
rect 14196 6554 14252 6556
rect 14276 6554 14332 6556
rect 14356 6554 14412 6556
rect 14116 6502 14142 6554
rect 14142 6502 14172 6554
rect 14196 6502 14206 6554
rect 14206 6502 14252 6554
rect 14276 6502 14322 6554
rect 14322 6502 14332 6554
rect 14356 6502 14386 6554
rect 14386 6502 14412 6554
rect 14116 6500 14172 6502
rect 14196 6500 14252 6502
rect 14276 6500 14332 6502
rect 14356 6500 14412 6502
rect 14116 5466 14172 5468
rect 14196 5466 14252 5468
rect 14276 5466 14332 5468
rect 14356 5466 14412 5468
rect 14116 5414 14142 5466
rect 14142 5414 14172 5466
rect 14196 5414 14206 5466
rect 14206 5414 14252 5466
rect 14276 5414 14322 5466
rect 14322 5414 14332 5466
rect 14356 5414 14386 5466
rect 14386 5414 14412 5466
rect 14116 5412 14172 5414
rect 14196 5412 14252 5414
rect 14276 5412 14332 5414
rect 14356 5412 14412 5414
rect 14116 4378 14172 4380
rect 14196 4378 14252 4380
rect 14276 4378 14332 4380
rect 14356 4378 14412 4380
rect 14116 4326 14142 4378
rect 14142 4326 14172 4378
rect 14196 4326 14206 4378
rect 14206 4326 14252 4378
rect 14276 4326 14322 4378
rect 14322 4326 14332 4378
rect 14356 4326 14386 4378
rect 14386 4326 14412 4378
rect 14116 4324 14172 4326
rect 14196 4324 14252 4326
rect 14276 4324 14332 4326
rect 14356 4324 14412 4326
rect 15106 5616 15162 5672
rect 15566 9152 15622 9208
rect 14116 3290 14172 3292
rect 14196 3290 14252 3292
rect 14276 3290 14332 3292
rect 14356 3290 14412 3292
rect 14116 3238 14142 3290
rect 14142 3238 14172 3290
rect 14196 3238 14206 3290
rect 14206 3238 14252 3290
rect 14276 3238 14322 3290
rect 14322 3238 14332 3290
rect 14356 3238 14386 3290
rect 14386 3238 14412 3290
rect 14116 3236 14172 3238
rect 14196 3236 14252 3238
rect 14276 3236 14332 3238
rect 14356 3236 14412 3238
rect 14116 2202 14172 2204
rect 14196 2202 14252 2204
rect 14276 2202 14332 2204
rect 14356 2202 14412 2204
rect 14116 2150 14142 2202
rect 14142 2150 14172 2202
rect 14196 2150 14206 2202
rect 14206 2150 14252 2202
rect 14276 2150 14322 2202
rect 14322 2150 14332 2202
rect 14356 2150 14386 2202
rect 14386 2150 14412 2202
rect 14116 2148 14172 2150
rect 14196 2148 14252 2150
rect 14276 2148 14332 2150
rect 14356 2148 14412 2150
rect 15106 3576 15162 3632
rect 16026 9832 16082 9888
rect 15934 9016 15990 9072
rect 16118 6976 16174 7032
rect 16026 6432 16082 6488
rect 16210 6024 16266 6080
rect 14830 1808 14886 1864
rect 14646 1400 14702 1456
rect 14554 584 14610 640
rect 2778 176 2834 232
rect 15106 992 15162 1048
rect 16026 5208 16082 5264
rect 16026 4800 16082 4856
rect 16026 4428 16028 4448
rect 16028 4428 16080 4448
rect 16080 4428 16082 4448
rect 16026 4392 16082 4428
rect 16026 3984 16082 4040
rect 16026 3032 16082 3088
rect 16026 2624 16082 2680
rect 16026 2252 16028 2272
rect 16028 2252 16080 2272
rect 16080 2252 16082 2272
rect 16026 2216 16082 2252
rect 14922 176 14978 232
<< metal3 >>
rect 0 16690 480 16720
rect 4797 16690 4863 16693
rect 0 16688 4863 16690
rect 0 16632 4802 16688
rect 4858 16632 4863 16688
rect 0 16630 4863 16632
rect 0 16600 480 16630
rect 4797 16627 4863 16630
rect 14917 16690 14983 16693
rect 17520 16690 18000 16720
rect 14917 16688 18000 16690
rect 14917 16632 14922 16688
rect 14978 16632 18000 16688
rect 14917 16630 18000 16632
rect 14917 16627 14983 16630
rect 17520 16600 18000 16630
rect 0 16282 480 16312
rect 3049 16282 3115 16285
rect 0 16280 3115 16282
rect 0 16224 3054 16280
rect 3110 16224 3115 16280
rect 0 16222 3115 16224
rect 0 16192 480 16222
rect 3049 16219 3115 16222
rect 16389 16282 16455 16285
rect 17520 16282 18000 16312
rect 16389 16280 18000 16282
rect 16389 16224 16394 16280
rect 16450 16224 18000 16280
rect 16389 16222 18000 16224
rect 16389 16219 16455 16222
rect 17520 16192 18000 16222
rect 0 15874 480 15904
rect 3141 15874 3207 15877
rect 0 15872 3207 15874
rect 0 15816 3146 15872
rect 3202 15816 3207 15872
rect 0 15814 3207 15816
rect 0 15784 480 15814
rect 3141 15811 3207 15814
rect 13169 15874 13235 15877
rect 17520 15874 18000 15904
rect 13169 15872 18000 15874
rect 13169 15816 13174 15872
rect 13230 15816 18000 15872
rect 13169 15814 18000 15816
rect 13169 15811 13235 15814
rect 17520 15784 18000 15814
rect 0 15466 480 15496
rect 3877 15466 3943 15469
rect 0 15464 3943 15466
rect 0 15408 3882 15464
rect 3938 15408 3943 15464
rect 0 15406 3943 15408
rect 0 15376 480 15406
rect 3877 15403 3943 15406
rect 14549 15466 14615 15469
rect 17520 15466 18000 15496
rect 14549 15464 18000 15466
rect 14549 15408 14554 15464
rect 14610 15408 18000 15464
rect 14549 15406 18000 15408
rect 14549 15403 14615 15406
rect 17520 15376 18000 15406
rect 0 15058 480 15088
rect 3509 15058 3575 15061
rect 0 15056 3575 15058
rect 0 15000 3514 15056
rect 3570 15000 3575 15056
rect 0 14998 3575 15000
rect 0 14968 480 14998
rect 3509 14995 3575 14998
rect 10593 15058 10659 15061
rect 17520 15058 18000 15088
rect 10593 15056 18000 15058
rect 10593 15000 10598 15056
rect 10654 15000 18000 15056
rect 10593 14998 18000 15000
rect 10593 14995 10659 14998
rect 17520 14968 18000 14998
rect 6208 14720 6528 14721
rect 0 14650 480 14680
rect 6208 14656 6216 14720
rect 6280 14656 6296 14720
rect 6360 14656 6376 14720
rect 6440 14656 6456 14720
rect 6520 14656 6528 14720
rect 6208 14655 6528 14656
rect 11472 14720 11792 14721
rect 11472 14656 11480 14720
rect 11544 14656 11560 14720
rect 11624 14656 11640 14720
rect 11704 14656 11720 14720
rect 11784 14656 11792 14720
rect 11472 14655 11792 14656
rect 5809 14650 5875 14653
rect 0 14648 5875 14650
rect 0 14592 5814 14648
rect 5870 14592 5875 14648
rect 0 14590 5875 14592
rect 0 14560 480 14590
rect 5809 14587 5875 14590
rect 13813 14650 13879 14653
rect 17520 14650 18000 14680
rect 13813 14648 18000 14650
rect 13813 14592 13818 14648
rect 13874 14592 18000 14648
rect 13813 14590 18000 14592
rect 13813 14587 13879 14590
rect 17520 14560 18000 14590
rect 0 14242 480 14272
rect 2313 14242 2379 14245
rect 17520 14242 18000 14272
rect 0 14240 2379 14242
rect 0 14184 2318 14240
rect 2374 14184 2379 14240
rect 0 14182 2379 14184
rect 0 14152 480 14182
rect 2313 14179 2379 14182
rect 15334 14182 18000 14242
rect 3576 14176 3896 14177
rect 3576 14112 3584 14176
rect 3648 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3896 14176
rect 3576 14111 3896 14112
rect 8840 14176 9160 14177
rect 8840 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9160 14176
rect 8840 14111 9160 14112
rect 14104 14176 14424 14177
rect 14104 14112 14112 14176
rect 14176 14112 14192 14176
rect 14256 14112 14272 14176
rect 14336 14112 14352 14176
rect 14416 14112 14424 14176
rect 14104 14111 14424 14112
rect 13905 13970 13971 13973
rect 15334 13970 15394 14182
rect 17520 14152 18000 14182
rect 13905 13968 15394 13970
rect 13905 13912 13910 13968
rect 13966 13912 15394 13968
rect 13905 13910 15394 13912
rect 13905 13907 13971 13910
rect 0 13834 480 13864
rect 2957 13834 3023 13837
rect 0 13832 3023 13834
rect 0 13776 2962 13832
rect 3018 13776 3023 13832
rect 0 13774 3023 13776
rect 0 13744 480 13774
rect 2957 13771 3023 13774
rect 16113 13834 16179 13837
rect 17520 13834 18000 13864
rect 16113 13832 18000 13834
rect 16113 13776 16118 13832
rect 16174 13776 18000 13832
rect 16113 13774 18000 13776
rect 16113 13771 16179 13774
rect 17520 13744 18000 13774
rect 6208 13632 6528 13633
rect 6208 13568 6216 13632
rect 6280 13568 6296 13632
rect 6360 13568 6376 13632
rect 6440 13568 6456 13632
rect 6520 13568 6528 13632
rect 6208 13567 6528 13568
rect 11472 13632 11792 13633
rect 11472 13568 11480 13632
rect 11544 13568 11560 13632
rect 11624 13568 11640 13632
rect 11704 13568 11720 13632
rect 11784 13568 11792 13632
rect 11472 13567 11792 13568
rect 0 13290 480 13320
rect 4153 13290 4219 13293
rect 0 13288 4219 13290
rect 0 13232 4158 13288
rect 4214 13232 4219 13288
rect 0 13230 4219 13232
rect 0 13200 480 13230
rect 4153 13227 4219 13230
rect 13077 13290 13143 13293
rect 17520 13290 18000 13320
rect 13077 13288 18000 13290
rect 13077 13232 13082 13288
rect 13138 13232 18000 13288
rect 13077 13230 18000 13232
rect 13077 13227 13143 13230
rect 17520 13200 18000 13230
rect 3576 13088 3896 13089
rect 3576 13024 3584 13088
rect 3648 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3896 13088
rect 3576 13023 3896 13024
rect 8840 13088 9160 13089
rect 8840 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9160 13088
rect 8840 13023 9160 13024
rect 14104 13088 14424 13089
rect 14104 13024 14112 13088
rect 14176 13024 14192 13088
rect 14256 13024 14272 13088
rect 14336 13024 14352 13088
rect 14416 13024 14424 13088
rect 14104 13023 14424 13024
rect 0 12882 480 12912
rect 3509 12882 3575 12885
rect 0 12880 3575 12882
rect 0 12824 3514 12880
rect 3570 12824 3575 12880
rect 0 12822 3575 12824
rect 0 12792 480 12822
rect 3509 12819 3575 12822
rect 14457 12882 14523 12885
rect 17520 12882 18000 12912
rect 14457 12880 18000 12882
rect 14457 12824 14462 12880
rect 14518 12824 18000 12880
rect 14457 12822 18000 12824
rect 14457 12819 14523 12822
rect 17520 12792 18000 12822
rect 6208 12544 6528 12545
rect 0 12474 480 12504
rect 6208 12480 6216 12544
rect 6280 12480 6296 12544
rect 6360 12480 6376 12544
rect 6440 12480 6456 12544
rect 6520 12480 6528 12544
rect 6208 12479 6528 12480
rect 11472 12544 11792 12545
rect 11472 12480 11480 12544
rect 11544 12480 11560 12544
rect 11624 12480 11640 12544
rect 11704 12480 11720 12544
rect 11784 12480 11792 12544
rect 11472 12479 11792 12480
rect 4061 12474 4127 12477
rect 0 12472 4127 12474
rect 0 12416 4066 12472
rect 4122 12416 4127 12472
rect 0 12414 4127 12416
rect 0 12384 480 12414
rect 4061 12411 4127 12414
rect 15009 12474 15075 12477
rect 17520 12474 18000 12504
rect 15009 12472 18000 12474
rect 15009 12416 15014 12472
rect 15070 12416 18000 12472
rect 15009 12414 18000 12416
rect 15009 12411 15075 12414
rect 17520 12384 18000 12414
rect 4153 12202 4219 12205
rect 8201 12202 8267 12205
rect 4153 12200 8267 12202
rect 4153 12144 4158 12200
rect 4214 12144 8206 12200
rect 8262 12144 8267 12200
rect 4153 12142 8267 12144
rect 4153 12139 4219 12142
rect 8201 12139 8267 12142
rect 0 12066 480 12096
rect 3417 12066 3483 12069
rect 0 12064 3483 12066
rect 0 12008 3422 12064
rect 3478 12008 3483 12064
rect 0 12006 3483 12008
rect 0 11976 480 12006
rect 3417 12003 3483 12006
rect 14825 12066 14891 12069
rect 15101 12066 15167 12069
rect 17520 12066 18000 12096
rect 14825 12064 18000 12066
rect 14825 12008 14830 12064
rect 14886 12008 15106 12064
rect 15162 12008 18000 12064
rect 14825 12006 18000 12008
rect 14825 12003 14891 12006
rect 15101 12003 15167 12006
rect 3576 12000 3896 12001
rect 3576 11936 3584 12000
rect 3648 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3896 12000
rect 3576 11935 3896 11936
rect 8840 12000 9160 12001
rect 8840 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9160 12000
rect 8840 11935 9160 11936
rect 14104 12000 14424 12001
rect 14104 11936 14112 12000
rect 14176 11936 14192 12000
rect 14256 11936 14272 12000
rect 14336 11936 14352 12000
rect 14416 11936 14424 12000
rect 17520 11976 18000 12006
rect 14104 11935 14424 11936
rect 2313 11794 2379 11797
rect 9397 11794 9463 11797
rect 2313 11792 9463 11794
rect 2313 11736 2318 11792
rect 2374 11736 9402 11792
rect 9458 11736 9463 11792
rect 2313 11734 9463 11736
rect 2313 11731 2379 11734
rect 9397 11731 9463 11734
rect 0 11658 480 11688
rect 2865 11658 2931 11661
rect 0 11656 2931 11658
rect 0 11600 2870 11656
rect 2926 11600 2931 11656
rect 0 11598 2931 11600
rect 0 11568 480 11598
rect 2865 11595 2931 11598
rect 15745 11658 15811 11661
rect 17520 11658 18000 11688
rect 15745 11656 18000 11658
rect 15745 11600 15750 11656
rect 15806 11600 18000 11656
rect 15745 11598 18000 11600
rect 15745 11595 15811 11598
rect 17520 11568 18000 11598
rect 7833 11522 7899 11525
rect 8017 11522 8083 11525
rect 7833 11520 8083 11522
rect 7833 11464 7838 11520
rect 7894 11464 8022 11520
rect 8078 11464 8083 11520
rect 7833 11462 8083 11464
rect 7833 11459 7899 11462
rect 8017 11459 8083 11462
rect 6208 11456 6528 11457
rect 6208 11392 6216 11456
rect 6280 11392 6296 11456
rect 6360 11392 6376 11456
rect 6440 11392 6456 11456
rect 6520 11392 6528 11456
rect 6208 11391 6528 11392
rect 11472 11456 11792 11457
rect 11472 11392 11480 11456
rect 11544 11392 11560 11456
rect 11624 11392 11640 11456
rect 11704 11392 11720 11456
rect 11784 11392 11792 11456
rect 11472 11391 11792 11392
rect 0 11250 480 11280
rect 4061 11250 4127 11253
rect 0 11248 4127 11250
rect 0 11192 4066 11248
rect 4122 11192 4127 11248
rect 0 11190 4127 11192
rect 0 11160 480 11190
rect 4061 11187 4127 11190
rect 4981 11250 5047 11253
rect 8293 11250 8359 11253
rect 4981 11248 8359 11250
rect 4981 11192 4986 11248
rect 5042 11192 8298 11248
rect 8354 11192 8359 11248
rect 4981 11190 8359 11192
rect 4981 11187 5047 11190
rect 8293 11187 8359 11190
rect 14825 11250 14891 11253
rect 17520 11250 18000 11280
rect 14825 11248 18000 11250
rect 14825 11192 14830 11248
rect 14886 11192 18000 11248
rect 14825 11190 18000 11192
rect 14825 11187 14891 11190
rect 17520 11160 18000 11190
rect 3576 10912 3896 10913
rect 0 10842 480 10872
rect 3576 10848 3584 10912
rect 3648 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3896 10912
rect 3576 10847 3896 10848
rect 8840 10912 9160 10913
rect 8840 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9160 10912
rect 8840 10847 9160 10848
rect 14104 10912 14424 10913
rect 14104 10848 14112 10912
rect 14176 10848 14192 10912
rect 14256 10848 14272 10912
rect 14336 10848 14352 10912
rect 14416 10848 14424 10912
rect 14104 10847 14424 10848
rect 3141 10842 3207 10845
rect 0 10840 3207 10842
rect 0 10784 3146 10840
rect 3202 10784 3207 10840
rect 0 10782 3207 10784
rect 0 10752 480 10782
rect 3141 10779 3207 10782
rect 15009 10842 15075 10845
rect 17520 10842 18000 10872
rect 15009 10840 18000 10842
rect 15009 10784 15014 10840
rect 15070 10784 18000 10840
rect 15009 10782 18000 10784
rect 15009 10779 15075 10782
rect 17520 10752 18000 10782
rect 2681 10570 2747 10573
rect 9213 10570 9279 10573
rect 2681 10568 9279 10570
rect 2681 10512 2686 10568
rect 2742 10512 9218 10568
rect 9274 10512 9279 10568
rect 2681 10510 9279 10512
rect 2681 10507 2747 10510
rect 9213 10507 9279 10510
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 13905 10434 13971 10437
rect 17520 10434 18000 10464
rect 13905 10432 18000 10434
rect 13905 10376 13910 10432
rect 13966 10376 18000 10432
rect 13905 10374 18000 10376
rect 13905 10371 13971 10374
rect 6208 10368 6528 10369
rect 6208 10304 6216 10368
rect 6280 10304 6296 10368
rect 6360 10304 6376 10368
rect 6440 10304 6456 10368
rect 6520 10304 6528 10368
rect 6208 10303 6528 10304
rect 11472 10368 11792 10369
rect 11472 10304 11480 10368
rect 11544 10304 11560 10368
rect 11624 10304 11640 10368
rect 11704 10304 11720 10368
rect 11784 10304 11792 10368
rect 17520 10344 18000 10374
rect 11472 10303 11792 10304
rect 2957 10298 3023 10301
rect 3325 10298 3391 10301
rect 2957 10296 3391 10298
rect 2957 10240 2962 10296
rect 3018 10240 3330 10296
rect 3386 10240 3391 10296
rect 2957 10238 3391 10240
rect 2957 10235 3023 10238
rect 3325 10235 3391 10238
rect 0 9890 480 9920
rect 2865 9890 2931 9893
rect 0 9888 2931 9890
rect 0 9832 2870 9888
rect 2926 9832 2931 9888
rect 0 9830 2931 9832
rect 0 9800 480 9830
rect 2865 9827 2931 9830
rect 16021 9890 16087 9893
rect 17520 9890 18000 9920
rect 16021 9888 18000 9890
rect 16021 9832 16026 9888
rect 16082 9832 18000 9888
rect 16021 9830 18000 9832
rect 16021 9827 16087 9830
rect 3576 9824 3896 9825
rect 3576 9760 3584 9824
rect 3648 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3896 9824
rect 3576 9759 3896 9760
rect 8840 9824 9160 9825
rect 8840 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9160 9824
rect 8840 9759 9160 9760
rect 14104 9824 14424 9825
rect 14104 9760 14112 9824
rect 14176 9760 14192 9824
rect 14256 9760 14272 9824
rect 14336 9760 14352 9824
rect 14416 9760 14424 9824
rect 17520 9800 18000 9830
rect 14104 9759 14424 9760
rect 10317 9754 10383 9757
rect 11053 9754 11119 9757
rect 10317 9752 11119 9754
rect 10317 9696 10322 9752
rect 10378 9696 11058 9752
rect 11114 9696 11119 9752
rect 10317 9694 11119 9696
rect 10317 9691 10383 9694
rect 11053 9691 11119 9694
rect 3509 9618 3575 9621
rect 4705 9618 4771 9621
rect 3509 9616 4771 9618
rect 3509 9560 3514 9616
rect 3570 9560 4710 9616
rect 4766 9560 4771 9616
rect 3509 9558 4771 9560
rect 3509 9555 3575 9558
rect 4705 9555 4771 9558
rect 10409 9618 10475 9621
rect 13629 9618 13695 9621
rect 10409 9616 13695 9618
rect 10409 9560 10414 9616
rect 10470 9560 13634 9616
rect 13690 9560 13695 9616
rect 10409 9558 13695 9560
rect 10409 9555 10475 9558
rect 13629 9555 13695 9558
rect 14641 9618 14707 9621
rect 14774 9618 14780 9620
rect 14641 9616 14780 9618
rect 14641 9560 14646 9616
rect 14702 9560 14780 9616
rect 14641 9558 14780 9560
rect 14641 9555 14707 9558
rect 14774 9556 14780 9558
rect 14844 9556 14850 9620
rect 0 9482 480 9512
rect 8569 9482 8635 9485
rect 9121 9482 9187 9485
rect 0 9480 9187 9482
rect 0 9424 8574 9480
rect 8630 9424 9126 9480
rect 9182 9424 9187 9480
rect 0 9422 9187 9424
rect 0 9392 480 9422
rect 8569 9419 8635 9422
rect 9121 9419 9187 9422
rect 10685 9482 10751 9485
rect 13077 9482 13143 9485
rect 17520 9482 18000 9512
rect 10685 9480 12634 9482
rect 10685 9424 10690 9480
rect 10746 9424 12634 9480
rect 10685 9422 12634 9424
rect 10685 9419 10751 9422
rect 12574 9346 12634 9422
rect 13077 9480 18000 9482
rect 13077 9424 13082 9480
rect 13138 9424 18000 9480
rect 13077 9422 18000 9424
rect 13077 9419 13143 9422
rect 17520 9392 18000 9422
rect 15377 9346 15443 9349
rect 12574 9344 15443 9346
rect 12574 9288 15382 9344
rect 15438 9288 15443 9344
rect 12574 9286 15443 9288
rect 15377 9283 15443 9286
rect 6208 9280 6528 9281
rect 6208 9216 6216 9280
rect 6280 9216 6296 9280
rect 6360 9216 6376 9280
rect 6440 9216 6456 9280
rect 6520 9216 6528 9280
rect 6208 9215 6528 9216
rect 11472 9280 11792 9281
rect 11472 9216 11480 9280
rect 11544 9216 11560 9280
rect 11624 9216 11640 9280
rect 11704 9216 11720 9280
rect 11784 9216 11792 9280
rect 11472 9215 11792 9216
rect 13261 9210 13327 9213
rect 15285 9210 15351 9213
rect 15561 9210 15627 9213
rect 13261 9208 15627 9210
rect 13261 9152 13266 9208
rect 13322 9152 15290 9208
rect 15346 9152 15566 9208
rect 15622 9152 15627 9208
rect 13261 9150 15627 9152
rect 13261 9147 13327 9150
rect 15285 9147 15351 9150
rect 15561 9147 15627 9150
rect 0 9074 480 9104
rect 2405 9074 2471 9077
rect 7741 9074 7807 9077
rect 0 9014 1778 9074
rect 0 8984 480 9014
rect 1718 8938 1778 9014
rect 2405 9072 7807 9074
rect 2405 9016 2410 9072
rect 2466 9016 7746 9072
rect 7802 9016 7807 9072
rect 2405 9014 7807 9016
rect 2405 9011 2471 9014
rect 7741 9011 7807 9014
rect 10593 9074 10659 9077
rect 15929 9074 15995 9077
rect 17520 9074 18000 9104
rect 10593 9072 18000 9074
rect 10593 9016 10598 9072
rect 10654 9016 15934 9072
rect 15990 9016 18000 9072
rect 10593 9014 18000 9016
rect 10593 9011 10659 9014
rect 15929 9011 15995 9014
rect 17520 8984 18000 9014
rect 2497 8938 2563 8941
rect 4521 8938 4587 8941
rect 7373 8938 7439 8941
rect 1718 8936 7439 8938
rect 1718 8880 2502 8936
rect 2558 8880 4526 8936
rect 4582 8880 7378 8936
rect 7434 8880 7439 8936
rect 1718 8878 7439 8880
rect 2497 8875 2563 8878
rect 4521 8875 4587 8878
rect 7373 8875 7439 8878
rect 3576 8736 3896 8737
rect 0 8666 480 8696
rect 3576 8672 3584 8736
rect 3648 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3896 8736
rect 3576 8671 3896 8672
rect 8840 8736 9160 8737
rect 8840 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9160 8736
rect 8840 8671 9160 8672
rect 14104 8736 14424 8737
rect 14104 8672 14112 8736
rect 14176 8672 14192 8736
rect 14256 8672 14272 8736
rect 14336 8672 14352 8736
rect 14416 8672 14424 8736
rect 14104 8671 14424 8672
rect 17520 8666 18000 8696
rect 0 8606 3434 8666
rect 0 8576 480 8606
rect 2773 8530 2839 8533
rect 2638 8528 2839 8530
rect 2638 8472 2778 8528
rect 2834 8472 2839 8528
rect 2638 8470 2839 8472
rect 3374 8530 3434 8606
rect 14598 8606 18000 8666
rect 8293 8530 8359 8533
rect 3374 8528 8359 8530
rect 3374 8472 8298 8528
rect 8354 8472 8359 8528
rect 3374 8470 8359 8472
rect 0 8258 480 8288
rect 2638 8258 2698 8470
rect 2773 8467 2839 8470
rect 8293 8467 8359 8470
rect 9857 8530 9923 8533
rect 11513 8530 11579 8533
rect 9857 8528 11579 8530
rect 9857 8472 9862 8528
rect 9918 8472 11518 8528
rect 11574 8472 11579 8528
rect 9857 8470 11579 8472
rect 9857 8467 9923 8470
rect 11513 8467 11579 8470
rect 14089 8530 14155 8533
rect 14598 8530 14658 8606
rect 17520 8576 18000 8606
rect 14089 8528 14658 8530
rect 14089 8472 14094 8528
rect 14150 8472 14658 8528
rect 14089 8470 14658 8472
rect 14089 8467 14155 8470
rect 0 8198 2698 8258
rect 14825 8258 14891 8261
rect 17520 8258 18000 8288
rect 14825 8256 18000 8258
rect 14825 8200 14830 8256
rect 14886 8200 18000 8256
rect 14825 8198 18000 8200
rect 0 8168 480 8198
rect 14825 8195 14891 8198
rect 6208 8192 6528 8193
rect 6208 8128 6216 8192
rect 6280 8128 6296 8192
rect 6360 8128 6376 8192
rect 6440 8128 6456 8192
rect 6520 8128 6528 8192
rect 6208 8127 6528 8128
rect 11472 8192 11792 8193
rect 11472 8128 11480 8192
rect 11544 8128 11560 8192
rect 11624 8128 11640 8192
rect 11704 8128 11720 8192
rect 11784 8128 11792 8192
rect 17520 8168 18000 8198
rect 11472 8127 11792 8128
rect 0 7850 480 7880
rect 3969 7850 4035 7853
rect 0 7848 4035 7850
rect 0 7792 3974 7848
rect 4030 7792 4035 7848
rect 0 7790 4035 7792
rect 0 7760 480 7790
rect 3969 7787 4035 7790
rect 11513 7850 11579 7853
rect 13169 7850 13235 7853
rect 11513 7848 13235 7850
rect 11513 7792 11518 7848
rect 11574 7792 13174 7848
rect 13230 7792 13235 7848
rect 11513 7790 13235 7792
rect 11513 7787 11579 7790
rect 13169 7787 13235 7790
rect 14641 7850 14707 7853
rect 17520 7850 18000 7880
rect 14641 7848 18000 7850
rect 14641 7792 14646 7848
rect 14702 7792 18000 7848
rect 14641 7790 18000 7792
rect 14641 7787 14707 7790
rect 17520 7760 18000 7790
rect 3576 7648 3896 7649
rect 3576 7584 3584 7648
rect 3648 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3896 7648
rect 3576 7583 3896 7584
rect 8840 7648 9160 7649
rect 8840 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9160 7648
rect 8840 7583 9160 7584
rect 14104 7648 14424 7649
rect 14104 7584 14112 7648
rect 14176 7584 14192 7648
rect 14256 7584 14272 7648
rect 14336 7584 14352 7648
rect 14416 7584 14424 7648
rect 14104 7583 14424 7584
rect 0 7442 480 7472
rect 4061 7442 4127 7445
rect 0 7440 4127 7442
rect 0 7384 4066 7440
rect 4122 7384 4127 7440
rect 0 7382 4127 7384
rect 0 7352 480 7382
rect 4061 7379 4127 7382
rect 14641 7442 14707 7445
rect 17520 7442 18000 7472
rect 14641 7440 18000 7442
rect 14641 7384 14646 7440
rect 14702 7384 18000 7440
rect 14641 7382 18000 7384
rect 14641 7379 14707 7382
rect 17520 7352 18000 7382
rect 12341 7306 12407 7309
rect 12893 7306 12959 7309
rect 12341 7304 12959 7306
rect 12341 7248 12346 7304
rect 12402 7248 12898 7304
rect 12954 7248 12959 7304
rect 12341 7246 12959 7248
rect 12341 7243 12407 7246
rect 12893 7243 12959 7246
rect 14365 7306 14431 7309
rect 14774 7306 14780 7308
rect 14365 7304 14780 7306
rect 14365 7248 14370 7304
rect 14426 7248 14780 7304
rect 14365 7246 14780 7248
rect 14365 7243 14431 7246
rect 14774 7244 14780 7246
rect 14844 7244 14850 7308
rect 4061 7170 4127 7173
rect 1350 7168 4127 7170
rect 1350 7112 4066 7168
rect 4122 7112 4127 7168
rect 1350 7110 4127 7112
rect 0 7034 480 7064
rect 1350 7034 1410 7110
rect 4061 7107 4127 7110
rect 6208 7104 6528 7105
rect 6208 7040 6216 7104
rect 6280 7040 6296 7104
rect 6360 7040 6376 7104
rect 6440 7040 6456 7104
rect 6520 7040 6528 7104
rect 6208 7039 6528 7040
rect 11472 7104 11792 7105
rect 11472 7040 11480 7104
rect 11544 7040 11560 7104
rect 11624 7040 11640 7104
rect 11704 7040 11720 7104
rect 11784 7040 11792 7104
rect 11472 7039 11792 7040
rect 0 6974 1410 7034
rect 16113 7034 16179 7037
rect 17520 7034 18000 7064
rect 16113 7032 18000 7034
rect 16113 6976 16118 7032
rect 16174 6976 18000 7032
rect 16113 6974 18000 6976
rect 0 6944 480 6974
rect 16113 6971 16179 6974
rect 17520 6944 18000 6974
rect 8201 6762 8267 6765
rect 9305 6762 9371 6765
rect 8201 6760 9371 6762
rect 8201 6704 8206 6760
rect 8262 6704 9310 6760
rect 9366 6704 9371 6760
rect 8201 6702 9371 6704
rect 8201 6699 8267 6702
rect 9305 6699 9371 6702
rect 3576 6560 3896 6561
rect 0 6490 480 6520
rect 3576 6496 3584 6560
rect 3648 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3896 6560
rect 3576 6495 3896 6496
rect 8840 6560 9160 6561
rect 8840 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9160 6560
rect 8840 6495 9160 6496
rect 14104 6560 14424 6561
rect 14104 6496 14112 6560
rect 14176 6496 14192 6560
rect 14256 6496 14272 6560
rect 14336 6496 14352 6560
rect 14416 6496 14424 6560
rect 14104 6495 14424 6496
rect 2957 6490 3023 6493
rect 0 6488 3023 6490
rect 0 6432 2962 6488
rect 3018 6432 3023 6488
rect 0 6430 3023 6432
rect 0 6400 480 6430
rect 2957 6427 3023 6430
rect 16021 6490 16087 6493
rect 17520 6490 18000 6520
rect 16021 6488 18000 6490
rect 16021 6432 16026 6488
rect 16082 6432 18000 6488
rect 16021 6430 18000 6432
rect 16021 6427 16087 6430
rect 17520 6400 18000 6430
rect 3417 6218 3483 6221
rect 1350 6216 3483 6218
rect 1350 6160 3422 6216
rect 3478 6160 3483 6216
rect 1350 6158 3483 6160
rect 0 6082 480 6112
rect 1350 6082 1410 6158
rect 3417 6155 3483 6158
rect 0 6022 1410 6082
rect 16205 6082 16271 6085
rect 17520 6082 18000 6112
rect 16205 6080 18000 6082
rect 16205 6024 16210 6080
rect 16266 6024 18000 6080
rect 16205 6022 18000 6024
rect 0 5992 480 6022
rect 16205 6019 16271 6022
rect 6208 6016 6528 6017
rect 6208 5952 6216 6016
rect 6280 5952 6296 6016
rect 6360 5952 6376 6016
rect 6440 5952 6456 6016
rect 6520 5952 6528 6016
rect 6208 5951 6528 5952
rect 11472 6016 11792 6017
rect 11472 5952 11480 6016
rect 11544 5952 11560 6016
rect 11624 5952 11640 6016
rect 11704 5952 11720 6016
rect 11784 5952 11792 6016
rect 17520 5992 18000 6022
rect 11472 5951 11792 5952
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 15101 5674 15167 5677
rect 17520 5674 18000 5704
rect 15101 5672 18000 5674
rect 15101 5616 15106 5672
rect 15162 5616 18000 5672
rect 15101 5614 18000 5616
rect 15101 5611 15167 5614
rect 17520 5584 18000 5614
rect 3576 5472 3896 5473
rect 3576 5408 3584 5472
rect 3648 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3896 5472
rect 3576 5407 3896 5408
rect 8840 5472 9160 5473
rect 8840 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9160 5472
rect 8840 5407 9160 5408
rect 14104 5472 14424 5473
rect 14104 5408 14112 5472
rect 14176 5408 14192 5472
rect 14256 5408 14272 5472
rect 14336 5408 14352 5472
rect 14416 5408 14424 5472
rect 14104 5407 14424 5408
rect 0 5266 480 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 480 5206
rect 4061 5203 4127 5206
rect 16021 5266 16087 5269
rect 17520 5266 18000 5296
rect 16021 5264 18000 5266
rect 16021 5208 16026 5264
rect 16082 5208 18000 5264
rect 16021 5206 18000 5208
rect 16021 5203 16087 5206
rect 17520 5176 18000 5206
rect 6208 4928 6528 4929
rect 0 4858 480 4888
rect 6208 4864 6216 4928
rect 6280 4864 6296 4928
rect 6360 4864 6376 4928
rect 6440 4864 6456 4928
rect 6520 4864 6528 4928
rect 6208 4863 6528 4864
rect 11472 4928 11792 4929
rect 11472 4864 11480 4928
rect 11544 4864 11560 4928
rect 11624 4864 11640 4928
rect 11704 4864 11720 4928
rect 11784 4864 11792 4928
rect 11472 4863 11792 4864
rect 2865 4858 2931 4861
rect 0 4856 2931 4858
rect 0 4800 2870 4856
rect 2926 4800 2931 4856
rect 0 4798 2931 4800
rect 0 4768 480 4798
rect 2865 4795 2931 4798
rect 16021 4858 16087 4861
rect 17520 4858 18000 4888
rect 16021 4856 18000 4858
rect 16021 4800 16026 4856
rect 16082 4800 18000 4856
rect 16021 4798 18000 4800
rect 16021 4795 16087 4798
rect 17520 4768 18000 4798
rect 0 4450 480 4480
rect 2773 4450 2839 4453
rect 0 4448 2839 4450
rect 0 4392 2778 4448
rect 2834 4392 2839 4448
rect 0 4390 2839 4392
rect 0 4360 480 4390
rect 2773 4387 2839 4390
rect 16021 4450 16087 4453
rect 17520 4450 18000 4480
rect 16021 4448 18000 4450
rect 16021 4392 16026 4448
rect 16082 4392 18000 4448
rect 16021 4390 18000 4392
rect 16021 4387 16087 4390
rect 3576 4384 3896 4385
rect 3576 4320 3584 4384
rect 3648 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3896 4384
rect 3576 4319 3896 4320
rect 8840 4384 9160 4385
rect 8840 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9160 4384
rect 8840 4319 9160 4320
rect 14104 4384 14424 4385
rect 14104 4320 14112 4384
rect 14176 4320 14192 4384
rect 14256 4320 14272 4384
rect 14336 4320 14352 4384
rect 14416 4320 14424 4384
rect 17520 4360 18000 4390
rect 14104 4319 14424 4320
rect 0 4042 480 4072
rect 4061 4042 4127 4045
rect 0 4040 4127 4042
rect 0 3984 4066 4040
rect 4122 3984 4127 4040
rect 0 3982 4127 3984
rect 0 3952 480 3982
rect 4061 3979 4127 3982
rect 16021 4042 16087 4045
rect 17520 4042 18000 4072
rect 16021 4040 18000 4042
rect 16021 3984 16026 4040
rect 16082 3984 18000 4040
rect 16021 3982 18000 3984
rect 16021 3979 16087 3982
rect 17520 3952 18000 3982
rect 6208 3840 6528 3841
rect 6208 3776 6216 3840
rect 6280 3776 6296 3840
rect 6360 3776 6376 3840
rect 6440 3776 6456 3840
rect 6520 3776 6528 3840
rect 6208 3775 6528 3776
rect 11472 3840 11792 3841
rect 11472 3776 11480 3840
rect 11544 3776 11560 3840
rect 11624 3776 11640 3840
rect 11704 3776 11720 3840
rect 11784 3776 11792 3840
rect 11472 3775 11792 3776
rect 0 3634 480 3664
rect 1577 3634 1643 3637
rect 0 3632 1643 3634
rect 0 3576 1582 3632
rect 1638 3576 1643 3632
rect 0 3574 1643 3576
rect 0 3544 480 3574
rect 1577 3571 1643 3574
rect 15101 3634 15167 3637
rect 17520 3634 18000 3664
rect 15101 3632 18000 3634
rect 15101 3576 15106 3632
rect 15162 3576 18000 3632
rect 15101 3574 18000 3576
rect 15101 3571 15167 3574
rect 17520 3544 18000 3574
rect 3576 3296 3896 3297
rect 3576 3232 3584 3296
rect 3648 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3896 3296
rect 3576 3231 3896 3232
rect 8840 3296 9160 3297
rect 8840 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9160 3296
rect 8840 3231 9160 3232
rect 14104 3296 14424 3297
rect 14104 3232 14112 3296
rect 14176 3232 14192 3296
rect 14256 3232 14272 3296
rect 14336 3232 14352 3296
rect 14416 3232 14424 3296
rect 14104 3231 14424 3232
rect 0 3090 480 3120
rect 3417 3090 3483 3093
rect 0 3088 3483 3090
rect 0 3032 3422 3088
rect 3478 3032 3483 3088
rect 0 3030 3483 3032
rect 0 3000 480 3030
rect 3417 3027 3483 3030
rect 16021 3090 16087 3093
rect 17520 3090 18000 3120
rect 16021 3088 18000 3090
rect 16021 3032 16026 3088
rect 16082 3032 18000 3088
rect 16021 3030 18000 3032
rect 16021 3027 16087 3030
rect 17520 3000 18000 3030
rect 6208 2752 6528 2753
rect 0 2682 480 2712
rect 6208 2688 6216 2752
rect 6280 2688 6296 2752
rect 6360 2688 6376 2752
rect 6440 2688 6456 2752
rect 6520 2688 6528 2752
rect 6208 2687 6528 2688
rect 11472 2752 11792 2753
rect 11472 2688 11480 2752
rect 11544 2688 11560 2752
rect 11624 2688 11640 2752
rect 11704 2688 11720 2752
rect 11784 2688 11792 2752
rect 11472 2687 11792 2688
rect 3325 2682 3391 2685
rect 0 2680 3391 2682
rect 0 2624 3330 2680
rect 3386 2624 3391 2680
rect 0 2622 3391 2624
rect 0 2592 480 2622
rect 3325 2619 3391 2622
rect 16021 2682 16087 2685
rect 17520 2682 18000 2712
rect 16021 2680 18000 2682
rect 16021 2624 16026 2680
rect 16082 2624 18000 2680
rect 16021 2622 18000 2624
rect 16021 2619 16087 2622
rect 17520 2592 18000 2622
rect 0 2274 480 2304
rect 2865 2274 2931 2277
rect 0 2272 2931 2274
rect 0 2216 2870 2272
rect 2926 2216 2931 2272
rect 0 2214 2931 2216
rect 0 2184 480 2214
rect 2865 2211 2931 2214
rect 16021 2274 16087 2277
rect 17520 2274 18000 2304
rect 16021 2272 18000 2274
rect 16021 2216 16026 2272
rect 16082 2216 18000 2272
rect 16021 2214 18000 2216
rect 16021 2211 16087 2214
rect 3576 2208 3896 2209
rect 3576 2144 3584 2208
rect 3648 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3896 2208
rect 3576 2143 3896 2144
rect 8840 2208 9160 2209
rect 8840 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9160 2208
rect 8840 2143 9160 2144
rect 14104 2208 14424 2209
rect 14104 2144 14112 2208
rect 14176 2144 14192 2208
rect 14256 2144 14272 2208
rect 14336 2144 14352 2208
rect 14416 2144 14424 2208
rect 17520 2184 18000 2214
rect 14104 2143 14424 2144
rect 0 1866 480 1896
rect 2957 1866 3023 1869
rect 0 1864 3023 1866
rect 0 1808 2962 1864
rect 3018 1808 3023 1864
rect 0 1806 3023 1808
rect 0 1776 480 1806
rect 2957 1803 3023 1806
rect 14825 1866 14891 1869
rect 17520 1866 18000 1896
rect 14825 1864 18000 1866
rect 14825 1808 14830 1864
rect 14886 1808 18000 1864
rect 14825 1806 18000 1808
rect 14825 1803 14891 1806
rect 17520 1776 18000 1806
rect 0 1458 480 1488
rect 2129 1458 2195 1461
rect 0 1456 2195 1458
rect 0 1400 2134 1456
rect 2190 1400 2195 1456
rect 0 1398 2195 1400
rect 0 1368 480 1398
rect 2129 1395 2195 1398
rect 14641 1458 14707 1461
rect 17520 1458 18000 1488
rect 14641 1456 18000 1458
rect 14641 1400 14646 1456
rect 14702 1400 18000 1456
rect 14641 1398 18000 1400
rect 14641 1395 14707 1398
rect 17520 1368 18000 1398
rect 0 1050 480 1080
rect 3049 1050 3115 1053
rect 0 1048 3115 1050
rect 0 992 3054 1048
rect 3110 992 3115 1048
rect 0 990 3115 992
rect 0 960 480 990
rect 3049 987 3115 990
rect 15101 1050 15167 1053
rect 17520 1050 18000 1080
rect 15101 1048 18000 1050
rect 15101 992 15106 1048
rect 15162 992 18000 1048
rect 15101 990 18000 992
rect 15101 987 15167 990
rect 17520 960 18000 990
rect 0 642 480 672
rect 3141 642 3207 645
rect 0 640 3207 642
rect 0 584 3146 640
rect 3202 584 3207 640
rect 0 582 3207 584
rect 0 552 480 582
rect 3141 579 3207 582
rect 14549 642 14615 645
rect 17520 642 18000 672
rect 14549 640 18000 642
rect 14549 584 14554 640
rect 14610 584 18000 640
rect 14549 582 18000 584
rect 14549 579 14615 582
rect 17520 552 18000 582
rect 0 234 480 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 480 174
rect 2773 171 2839 174
rect 14917 234 14983 237
rect 17520 234 18000 264
rect 14917 232 18000 234
rect 14917 176 14922 232
rect 14978 176 18000 232
rect 14917 174 18000 176
rect 14917 171 14983 174
rect 17520 144 18000 174
<< via3 >>
rect 6216 14716 6280 14720
rect 6216 14660 6220 14716
rect 6220 14660 6276 14716
rect 6276 14660 6280 14716
rect 6216 14656 6280 14660
rect 6296 14716 6360 14720
rect 6296 14660 6300 14716
rect 6300 14660 6356 14716
rect 6356 14660 6360 14716
rect 6296 14656 6360 14660
rect 6376 14716 6440 14720
rect 6376 14660 6380 14716
rect 6380 14660 6436 14716
rect 6436 14660 6440 14716
rect 6376 14656 6440 14660
rect 6456 14716 6520 14720
rect 6456 14660 6460 14716
rect 6460 14660 6516 14716
rect 6516 14660 6520 14716
rect 6456 14656 6520 14660
rect 11480 14716 11544 14720
rect 11480 14660 11484 14716
rect 11484 14660 11540 14716
rect 11540 14660 11544 14716
rect 11480 14656 11544 14660
rect 11560 14716 11624 14720
rect 11560 14660 11564 14716
rect 11564 14660 11620 14716
rect 11620 14660 11624 14716
rect 11560 14656 11624 14660
rect 11640 14716 11704 14720
rect 11640 14660 11644 14716
rect 11644 14660 11700 14716
rect 11700 14660 11704 14716
rect 11640 14656 11704 14660
rect 11720 14716 11784 14720
rect 11720 14660 11724 14716
rect 11724 14660 11780 14716
rect 11780 14660 11784 14716
rect 11720 14656 11784 14660
rect 3584 14172 3648 14176
rect 3584 14116 3588 14172
rect 3588 14116 3644 14172
rect 3644 14116 3648 14172
rect 3584 14112 3648 14116
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 8848 14172 8912 14176
rect 8848 14116 8852 14172
rect 8852 14116 8908 14172
rect 8908 14116 8912 14172
rect 8848 14112 8912 14116
rect 8928 14172 8992 14176
rect 8928 14116 8932 14172
rect 8932 14116 8988 14172
rect 8988 14116 8992 14172
rect 8928 14112 8992 14116
rect 9008 14172 9072 14176
rect 9008 14116 9012 14172
rect 9012 14116 9068 14172
rect 9068 14116 9072 14172
rect 9008 14112 9072 14116
rect 9088 14172 9152 14176
rect 9088 14116 9092 14172
rect 9092 14116 9148 14172
rect 9148 14116 9152 14172
rect 9088 14112 9152 14116
rect 14112 14172 14176 14176
rect 14112 14116 14116 14172
rect 14116 14116 14172 14172
rect 14172 14116 14176 14172
rect 14112 14112 14176 14116
rect 14192 14172 14256 14176
rect 14192 14116 14196 14172
rect 14196 14116 14252 14172
rect 14252 14116 14256 14172
rect 14192 14112 14256 14116
rect 14272 14172 14336 14176
rect 14272 14116 14276 14172
rect 14276 14116 14332 14172
rect 14332 14116 14336 14172
rect 14272 14112 14336 14116
rect 14352 14172 14416 14176
rect 14352 14116 14356 14172
rect 14356 14116 14412 14172
rect 14412 14116 14416 14172
rect 14352 14112 14416 14116
rect 6216 13628 6280 13632
rect 6216 13572 6220 13628
rect 6220 13572 6276 13628
rect 6276 13572 6280 13628
rect 6216 13568 6280 13572
rect 6296 13628 6360 13632
rect 6296 13572 6300 13628
rect 6300 13572 6356 13628
rect 6356 13572 6360 13628
rect 6296 13568 6360 13572
rect 6376 13628 6440 13632
rect 6376 13572 6380 13628
rect 6380 13572 6436 13628
rect 6436 13572 6440 13628
rect 6376 13568 6440 13572
rect 6456 13628 6520 13632
rect 6456 13572 6460 13628
rect 6460 13572 6516 13628
rect 6516 13572 6520 13628
rect 6456 13568 6520 13572
rect 11480 13628 11544 13632
rect 11480 13572 11484 13628
rect 11484 13572 11540 13628
rect 11540 13572 11544 13628
rect 11480 13568 11544 13572
rect 11560 13628 11624 13632
rect 11560 13572 11564 13628
rect 11564 13572 11620 13628
rect 11620 13572 11624 13628
rect 11560 13568 11624 13572
rect 11640 13628 11704 13632
rect 11640 13572 11644 13628
rect 11644 13572 11700 13628
rect 11700 13572 11704 13628
rect 11640 13568 11704 13572
rect 11720 13628 11784 13632
rect 11720 13572 11724 13628
rect 11724 13572 11780 13628
rect 11780 13572 11784 13628
rect 11720 13568 11784 13572
rect 3584 13084 3648 13088
rect 3584 13028 3588 13084
rect 3588 13028 3644 13084
rect 3644 13028 3648 13084
rect 3584 13024 3648 13028
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 8848 13084 8912 13088
rect 8848 13028 8852 13084
rect 8852 13028 8908 13084
rect 8908 13028 8912 13084
rect 8848 13024 8912 13028
rect 8928 13084 8992 13088
rect 8928 13028 8932 13084
rect 8932 13028 8988 13084
rect 8988 13028 8992 13084
rect 8928 13024 8992 13028
rect 9008 13084 9072 13088
rect 9008 13028 9012 13084
rect 9012 13028 9068 13084
rect 9068 13028 9072 13084
rect 9008 13024 9072 13028
rect 9088 13084 9152 13088
rect 9088 13028 9092 13084
rect 9092 13028 9148 13084
rect 9148 13028 9152 13084
rect 9088 13024 9152 13028
rect 14112 13084 14176 13088
rect 14112 13028 14116 13084
rect 14116 13028 14172 13084
rect 14172 13028 14176 13084
rect 14112 13024 14176 13028
rect 14192 13084 14256 13088
rect 14192 13028 14196 13084
rect 14196 13028 14252 13084
rect 14252 13028 14256 13084
rect 14192 13024 14256 13028
rect 14272 13084 14336 13088
rect 14272 13028 14276 13084
rect 14276 13028 14332 13084
rect 14332 13028 14336 13084
rect 14272 13024 14336 13028
rect 14352 13084 14416 13088
rect 14352 13028 14356 13084
rect 14356 13028 14412 13084
rect 14412 13028 14416 13084
rect 14352 13024 14416 13028
rect 6216 12540 6280 12544
rect 6216 12484 6220 12540
rect 6220 12484 6276 12540
rect 6276 12484 6280 12540
rect 6216 12480 6280 12484
rect 6296 12540 6360 12544
rect 6296 12484 6300 12540
rect 6300 12484 6356 12540
rect 6356 12484 6360 12540
rect 6296 12480 6360 12484
rect 6376 12540 6440 12544
rect 6376 12484 6380 12540
rect 6380 12484 6436 12540
rect 6436 12484 6440 12540
rect 6376 12480 6440 12484
rect 6456 12540 6520 12544
rect 6456 12484 6460 12540
rect 6460 12484 6516 12540
rect 6516 12484 6520 12540
rect 6456 12480 6520 12484
rect 11480 12540 11544 12544
rect 11480 12484 11484 12540
rect 11484 12484 11540 12540
rect 11540 12484 11544 12540
rect 11480 12480 11544 12484
rect 11560 12540 11624 12544
rect 11560 12484 11564 12540
rect 11564 12484 11620 12540
rect 11620 12484 11624 12540
rect 11560 12480 11624 12484
rect 11640 12540 11704 12544
rect 11640 12484 11644 12540
rect 11644 12484 11700 12540
rect 11700 12484 11704 12540
rect 11640 12480 11704 12484
rect 11720 12540 11784 12544
rect 11720 12484 11724 12540
rect 11724 12484 11780 12540
rect 11780 12484 11784 12540
rect 11720 12480 11784 12484
rect 3584 11996 3648 12000
rect 3584 11940 3588 11996
rect 3588 11940 3644 11996
rect 3644 11940 3648 11996
rect 3584 11936 3648 11940
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 8848 11996 8912 12000
rect 8848 11940 8852 11996
rect 8852 11940 8908 11996
rect 8908 11940 8912 11996
rect 8848 11936 8912 11940
rect 8928 11996 8992 12000
rect 8928 11940 8932 11996
rect 8932 11940 8988 11996
rect 8988 11940 8992 11996
rect 8928 11936 8992 11940
rect 9008 11996 9072 12000
rect 9008 11940 9012 11996
rect 9012 11940 9068 11996
rect 9068 11940 9072 11996
rect 9008 11936 9072 11940
rect 9088 11996 9152 12000
rect 9088 11940 9092 11996
rect 9092 11940 9148 11996
rect 9148 11940 9152 11996
rect 9088 11936 9152 11940
rect 14112 11996 14176 12000
rect 14112 11940 14116 11996
rect 14116 11940 14172 11996
rect 14172 11940 14176 11996
rect 14112 11936 14176 11940
rect 14192 11996 14256 12000
rect 14192 11940 14196 11996
rect 14196 11940 14252 11996
rect 14252 11940 14256 11996
rect 14192 11936 14256 11940
rect 14272 11996 14336 12000
rect 14272 11940 14276 11996
rect 14276 11940 14332 11996
rect 14332 11940 14336 11996
rect 14272 11936 14336 11940
rect 14352 11996 14416 12000
rect 14352 11940 14356 11996
rect 14356 11940 14412 11996
rect 14412 11940 14416 11996
rect 14352 11936 14416 11940
rect 6216 11452 6280 11456
rect 6216 11396 6220 11452
rect 6220 11396 6276 11452
rect 6276 11396 6280 11452
rect 6216 11392 6280 11396
rect 6296 11452 6360 11456
rect 6296 11396 6300 11452
rect 6300 11396 6356 11452
rect 6356 11396 6360 11452
rect 6296 11392 6360 11396
rect 6376 11452 6440 11456
rect 6376 11396 6380 11452
rect 6380 11396 6436 11452
rect 6436 11396 6440 11452
rect 6376 11392 6440 11396
rect 6456 11452 6520 11456
rect 6456 11396 6460 11452
rect 6460 11396 6516 11452
rect 6516 11396 6520 11452
rect 6456 11392 6520 11396
rect 11480 11452 11544 11456
rect 11480 11396 11484 11452
rect 11484 11396 11540 11452
rect 11540 11396 11544 11452
rect 11480 11392 11544 11396
rect 11560 11452 11624 11456
rect 11560 11396 11564 11452
rect 11564 11396 11620 11452
rect 11620 11396 11624 11452
rect 11560 11392 11624 11396
rect 11640 11452 11704 11456
rect 11640 11396 11644 11452
rect 11644 11396 11700 11452
rect 11700 11396 11704 11452
rect 11640 11392 11704 11396
rect 11720 11452 11784 11456
rect 11720 11396 11724 11452
rect 11724 11396 11780 11452
rect 11780 11396 11784 11452
rect 11720 11392 11784 11396
rect 3584 10908 3648 10912
rect 3584 10852 3588 10908
rect 3588 10852 3644 10908
rect 3644 10852 3648 10908
rect 3584 10848 3648 10852
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 8848 10908 8912 10912
rect 8848 10852 8852 10908
rect 8852 10852 8908 10908
rect 8908 10852 8912 10908
rect 8848 10848 8912 10852
rect 8928 10908 8992 10912
rect 8928 10852 8932 10908
rect 8932 10852 8988 10908
rect 8988 10852 8992 10908
rect 8928 10848 8992 10852
rect 9008 10908 9072 10912
rect 9008 10852 9012 10908
rect 9012 10852 9068 10908
rect 9068 10852 9072 10908
rect 9008 10848 9072 10852
rect 9088 10908 9152 10912
rect 9088 10852 9092 10908
rect 9092 10852 9148 10908
rect 9148 10852 9152 10908
rect 9088 10848 9152 10852
rect 14112 10908 14176 10912
rect 14112 10852 14116 10908
rect 14116 10852 14172 10908
rect 14172 10852 14176 10908
rect 14112 10848 14176 10852
rect 14192 10908 14256 10912
rect 14192 10852 14196 10908
rect 14196 10852 14252 10908
rect 14252 10852 14256 10908
rect 14192 10848 14256 10852
rect 14272 10908 14336 10912
rect 14272 10852 14276 10908
rect 14276 10852 14332 10908
rect 14332 10852 14336 10908
rect 14272 10848 14336 10852
rect 14352 10908 14416 10912
rect 14352 10852 14356 10908
rect 14356 10852 14412 10908
rect 14412 10852 14416 10908
rect 14352 10848 14416 10852
rect 6216 10364 6280 10368
rect 6216 10308 6220 10364
rect 6220 10308 6276 10364
rect 6276 10308 6280 10364
rect 6216 10304 6280 10308
rect 6296 10364 6360 10368
rect 6296 10308 6300 10364
rect 6300 10308 6356 10364
rect 6356 10308 6360 10364
rect 6296 10304 6360 10308
rect 6376 10364 6440 10368
rect 6376 10308 6380 10364
rect 6380 10308 6436 10364
rect 6436 10308 6440 10364
rect 6376 10304 6440 10308
rect 6456 10364 6520 10368
rect 6456 10308 6460 10364
rect 6460 10308 6516 10364
rect 6516 10308 6520 10364
rect 6456 10304 6520 10308
rect 11480 10364 11544 10368
rect 11480 10308 11484 10364
rect 11484 10308 11540 10364
rect 11540 10308 11544 10364
rect 11480 10304 11544 10308
rect 11560 10364 11624 10368
rect 11560 10308 11564 10364
rect 11564 10308 11620 10364
rect 11620 10308 11624 10364
rect 11560 10304 11624 10308
rect 11640 10364 11704 10368
rect 11640 10308 11644 10364
rect 11644 10308 11700 10364
rect 11700 10308 11704 10364
rect 11640 10304 11704 10308
rect 11720 10364 11784 10368
rect 11720 10308 11724 10364
rect 11724 10308 11780 10364
rect 11780 10308 11784 10364
rect 11720 10304 11784 10308
rect 3584 9820 3648 9824
rect 3584 9764 3588 9820
rect 3588 9764 3644 9820
rect 3644 9764 3648 9820
rect 3584 9760 3648 9764
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 8848 9820 8912 9824
rect 8848 9764 8852 9820
rect 8852 9764 8908 9820
rect 8908 9764 8912 9820
rect 8848 9760 8912 9764
rect 8928 9820 8992 9824
rect 8928 9764 8932 9820
rect 8932 9764 8988 9820
rect 8988 9764 8992 9820
rect 8928 9760 8992 9764
rect 9008 9820 9072 9824
rect 9008 9764 9012 9820
rect 9012 9764 9068 9820
rect 9068 9764 9072 9820
rect 9008 9760 9072 9764
rect 9088 9820 9152 9824
rect 9088 9764 9092 9820
rect 9092 9764 9148 9820
rect 9148 9764 9152 9820
rect 9088 9760 9152 9764
rect 14112 9820 14176 9824
rect 14112 9764 14116 9820
rect 14116 9764 14172 9820
rect 14172 9764 14176 9820
rect 14112 9760 14176 9764
rect 14192 9820 14256 9824
rect 14192 9764 14196 9820
rect 14196 9764 14252 9820
rect 14252 9764 14256 9820
rect 14192 9760 14256 9764
rect 14272 9820 14336 9824
rect 14272 9764 14276 9820
rect 14276 9764 14332 9820
rect 14332 9764 14336 9820
rect 14272 9760 14336 9764
rect 14352 9820 14416 9824
rect 14352 9764 14356 9820
rect 14356 9764 14412 9820
rect 14412 9764 14416 9820
rect 14352 9760 14416 9764
rect 14780 9556 14844 9620
rect 6216 9276 6280 9280
rect 6216 9220 6220 9276
rect 6220 9220 6276 9276
rect 6276 9220 6280 9276
rect 6216 9216 6280 9220
rect 6296 9276 6360 9280
rect 6296 9220 6300 9276
rect 6300 9220 6356 9276
rect 6356 9220 6360 9276
rect 6296 9216 6360 9220
rect 6376 9276 6440 9280
rect 6376 9220 6380 9276
rect 6380 9220 6436 9276
rect 6436 9220 6440 9276
rect 6376 9216 6440 9220
rect 6456 9276 6520 9280
rect 6456 9220 6460 9276
rect 6460 9220 6516 9276
rect 6516 9220 6520 9276
rect 6456 9216 6520 9220
rect 11480 9276 11544 9280
rect 11480 9220 11484 9276
rect 11484 9220 11540 9276
rect 11540 9220 11544 9276
rect 11480 9216 11544 9220
rect 11560 9276 11624 9280
rect 11560 9220 11564 9276
rect 11564 9220 11620 9276
rect 11620 9220 11624 9276
rect 11560 9216 11624 9220
rect 11640 9276 11704 9280
rect 11640 9220 11644 9276
rect 11644 9220 11700 9276
rect 11700 9220 11704 9276
rect 11640 9216 11704 9220
rect 11720 9276 11784 9280
rect 11720 9220 11724 9276
rect 11724 9220 11780 9276
rect 11780 9220 11784 9276
rect 11720 9216 11784 9220
rect 3584 8732 3648 8736
rect 3584 8676 3588 8732
rect 3588 8676 3644 8732
rect 3644 8676 3648 8732
rect 3584 8672 3648 8676
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 8848 8732 8912 8736
rect 8848 8676 8852 8732
rect 8852 8676 8908 8732
rect 8908 8676 8912 8732
rect 8848 8672 8912 8676
rect 8928 8732 8992 8736
rect 8928 8676 8932 8732
rect 8932 8676 8988 8732
rect 8988 8676 8992 8732
rect 8928 8672 8992 8676
rect 9008 8732 9072 8736
rect 9008 8676 9012 8732
rect 9012 8676 9068 8732
rect 9068 8676 9072 8732
rect 9008 8672 9072 8676
rect 9088 8732 9152 8736
rect 9088 8676 9092 8732
rect 9092 8676 9148 8732
rect 9148 8676 9152 8732
rect 9088 8672 9152 8676
rect 14112 8732 14176 8736
rect 14112 8676 14116 8732
rect 14116 8676 14172 8732
rect 14172 8676 14176 8732
rect 14112 8672 14176 8676
rect 14192 8732 14256 8736
rect 14192 8676 14196 8732
rect 14196 8676 14252 8732
rect 14252 8676 14256 8732
rect 14192 8672 14256 8676
rect 14272 8732 14336 8736
rect 14272 8676 14276 8732
rect 14276 8676 14332 8732
rect 14332 8676 14336 8732
rect 14272 8672 14336 8676
rect 14352 8732 14416 8736
rect 14352 8676 14356 8732
rect 14356 8676 14412 8732
rect 14412 8676 14416 8732
rect 14352 8672 14416 8676
rect 6216 8188 6280 8192
rect 6216 8132 6220 8188
rect 6220 8132 6276 8188
rect 6276 8132 6280 8188
rect 6216 8128 6280 8132
rect 6296 8188 6360 8192
rect 6296 8132 6300 8188
rect 6300 8132 6356 8188
rect 6356 8132 6360 8188
rect 6296 8128 6360 8132
rect 6376 8188 6440 8192
rect 6376 8132 6380 8188
rect 6380 8132 6436 8188
rect 6436 8132 6440 8188
rect 6376 8128 6440 8132
rect 6456 8188 6520 8192
rect 6456 8132 6460 8188
rect 6460 8132 6516 8188
rect 6516 8132 6520 8188
rect 6456 8128 6520 8132
rect 11480 8188 11544 8192
rect 11480 8132 11484 8188
rect 11484 8132 11540 8188
rect 11540 8132 11544 8188
rect 11480 8128 11544 8132
rect 11560 8188 11624 8192
rect 11560 8132 11564 8188
rect 11564 8132 11620 8188
rect 11620 8132 11624 8188
rect 11560 8128 11624 8132
rect 11640 8188 11704 8192
rect 11640 8132 11644 8188
rect 11644 8132 11700 8188
rect 11700 8132 11704 8188
rect 11640 8128 11704 8132
rect 11720 8188 11784 8192
rect 11720 8132 11724 8188
rect 11724 8132 11780 8188
rect 11780 8132 11784 8188
rect 11720 8128 11784 8132
rect 3584 7644 3648 7648
rect 3584 7588 3588 7644
rect 3588 7588 3644 7644
rect 3644 7588 3648 7644
rect 3584 7584 3648 7588
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 8848 7644 8912 7648
rect 8848 7588 8852 7644
rect 8852 7588 8908 7644
rect 8908 7588 8912 7644
rect 8848 7584 8912 7588
rect 8928 7644 8992 7648
rect 8928 7588 8932 7644
rect 8932 7588 8988 7644
rect 8988 7588 8992 7644
rect 8928 7584 8992 7588
rect 9008 7644 9072 7648
rect 9008 7588 9012 7644
rect 9012 7588 9068 7644
rect 9068 7588 9072 7644
rect 9008 7584 9072 7588
rect 9088 7644 9152 7648
rect 9088 7588 9092 7644
rect 9092 7588 9148 7644
rect 9148 7588 9152 7644
rect 9088 7584 9152 7588
rect 14112 7644 14176 7648
rect 14112 7588 14116 7644
rect 14116 7588 14172 7644
rect 14172 7588 14176 7644
rect 14112 7584 14176 7588
rect 14192 7644 14256 7648
rect 14192 7588 14196 7644
rect 14196 7588 14252 7644
rect 14252 7588 14256 7644
rect 14192 7584 14256 7588
rect 14272 7644 14336 7648
rect 14272 7588 14276 7644
rect 14276 7588 14332 7644
rect 14332 7588 14336 7644
rect 14272 7584 14336 7588
rect 14352 7644 14416 7648
rect 14352 7588 14356 7644
rect 14356 7588 14412 7644
rect 14412 7588 14416 7644
rect 14352 7584 14416 7588
rect 14780 7244 14844 7308
rect 6216 7100 6280 7104
rect 6216 7044 6220 7100
rect 6220 7044 6276 7100
rect 6276 7044 6280 7100
rect 6216 7040 6280 7044
rect 6296 7100 6360 7104
rect 6296 7044 6300 7100
rect 6300 7044 6356 7100
rect 6356 7044 6360 7100
rect 6296 7040 6360 7044
rect 6376 7100 6440 7104
rect 6376 7044 6380 7100
rect 6380 7044 6436 7100
rect 6436 7044 6440 7100
rect 6376 7040 6440 7044
rect 6456 7100 6520 7104
rect 6456 7044 6460 7100
rect 6460 7044 6516 7100
rect 6516 7044 6520 7100
rect 6456 7040 6520 7044
rect 11480 7100 11544 7104
rect 11480 7044 11484 7100
rect 11484 7044 11540 7100
rect 11540 7044 11544 7100
rect 11480 7040 11544 7044
rect 11560 7100 11624 7104
rect 11560 7044 11564 7100
rect 11564 7044 11620 7100
rect 11620 7044 11624 7100
rect 11560 7040 11624 7044
rect 11640 7100 11704 7104
rect 11640 7044 11644 7100
rect 11644 7044 11700 7100
rect 11700 7044 11704 7100
rect 11640 7040 11704 7044
rect 11720 7100 11784 7104
rect 11720 7044 11724 7100
rect 11724 7044 11780 7100
rect 11780 7044 11784 7100
rect 11720 7040 11784 7044
rect 3584 6556 3648 6560
rect 3584 6500 3588 6556
rect 3588 6500 3644 6556
rect 3644 6500 3648 6556
rect 3584 6496 3648 6500
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 8848 6556 8912 6560
rect 8848 6500 8852 6556
rect 8852 6500 8908 6556
rect 8908 6500 8912 6556
rect 8848 6496 8912 6500
rect 8928 6556 8992 6560
rect 8928 6500 8932 6556
rect 8932 6500 8988 6556
rect 8988 6500 8992 6556
rect 8928 6496 8992 6500
rect 9008 6556 9072 6560
rect 9008 6500 9012 6556
rect 9012 6500 9068 6556
rect 9068 6500 9072 6556
rect 9008 6496 9072 6500
rect 9088 6556 9152 6560
rect 9088 6500 9092 6556
rect 9092 6500 9148 6556
rect 9148 6500 9152 6556
rect 9088 6496 9152 6500
rect 14112 6556 14176 6560
rect 14112 6500 14116 6556
rect 14116 6500 14172 6556
rect 14172 6500 14176 6556
rect 14112 6496 14176 6500
rect 14192 6556 14256 6560
rect 14192 6500 14196 6556
rect 14196 6500 14252 6556
rect 14252 6500 14256 6556
rect 14192 6496 14256 6500
rect 14272 6556 14336 6560
rect 14272 6500 14276 6556
rect 14276 6500 14332 6556
rect 14332 6500 14336 6556
rect 14272 6496 14336 6500
rect 14352 6556 14416 6560
rect 14352 6500 14356 6556
rect 14356 6500 14412 6556
rect 14412 6500 14416 6556
rect 14352 6496 14416 6500
rect 6216 6012 6280 6016
rect 6216 5956 6220 6012
rect 6220 5956 6276 6012
rect 6276 5956 6280 6012
rect 6216 5952 6280 5956
rect 6296 6012 6360 6016
rect 6296 5956 6300 6012
rect 6300 5956 6356 6012
rect 6356 5956 6360 6012
rect 6296 5952 6360 5956
rect 6376 6012 6440 6016
rect 6376 5956 6380 6012
rect 6380 5956 6436 6012
rect 6436 5956 6440 6012
rect 6376 5952 6440 5956
rect 6456 6012 6520 6016
rect 6456 5956 6460 6012
rect 6460 5956 6516 6012
rect 6516 5956 6520 6012
rect 6456 5952 6520 5956
rect 11480 6012 11544 6016
rect 11480 5956 11484 6012
rect 11484 5956 11540 6012
rect 11540 5956 11544 6012
rect 11480 5952 11544 5956
rect 11560 6012 11624 6016
rect 11560 5956 11564 6012
rect 11564 5956 11620 6012
rect 11620 5956 11624 6012
rect 11560 5952 11624 5956
rect 11640 6012 11704 6016
rect 11640 5956 11644 6012
rect 11644 5956 11700 6012
rect 11700 5956 11704 6012
rect 11640 5952 11704 5956
rect 11720 6012 11784 6016
rect 11720 5956 11724 6012
rect 11724 5956 11780 6012
rect 11780 5956 11784 6012
rect 11720 5952 11784 5956
rect 3584 5468 3648 5472
rect 3584 5412 3588 5468
rect 3588 5412 3644 5468
rect 3644 5412 3648 5468
rect 3584 5408 3648 5412
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 8848 5468 8912 5472
rect 8848 5412 8852 5468
rect 8852 5412 8908 5468
rect 8908 5412 8912 5468
rect 8848 5408 8912 5412
rect 8928 5468 8992 5472
rect 8928 5412 8932 5468
rect 8932 5412 8988 5468
rect 8988 5412 8992 5468
rect 8928 5408 8992 5412
rect 9008 5468 9072 5472
rect 9008 5412 9012 5468
rect 9012 5412 9068 5468
rect 9068 5412 9072 5468
rect 9008 5408 9072 5412
rect 9088 5468 9152 5472
rect 9088 5412 9092 5468
rect 9092 5412 9148 5468
rect 9148 5412 9152 5468
rect 9088 5408 9152 5412
rect 14112 5468 14176 5472
rect 14112 5412 14116 5468
rect 14116 5412 14172 5468
rect 14172 5412 14176 5468
rect 14112 5408 14176 5412
rect 14192 5468 14256 5472
rect 14192 5412 14196 5468
rect 14196 5412 14252 5468
rect 14252 5412 14256 5468
rect 14192 5408 14256 5412
rect 14272 5468 14336 5472
rect 14272 5412 14276 5468
rect 14276 5412 14332 5468
rect 14332 5412 14336 5468
rect 14272 5408 14336 5412
rect 14352 5468 14416 5472
rect 14352 5412 14356 5468
rect 14356 5412 14412 5468
rect 14412 5412 14416 5468
rect 14352 5408 14416 5412
rect 6216 4924 6280 4928
rect 6216 4868 6220 4924
rect 6220 4868 6276 4924
rect 6276 4868 6280 4924
rect 6216 4864 6280 4868
rect 6296 4924 6360 4928
rect 6296 4868 6300 4924
rect 6300 4868 6356 4924
rect 6356 4868 6360 4924
rect 6296 4864 6360 4868
rect 6376 4924 6440 4928
rect 6376 4868 6380 4924
rect 6380 4868 6436 4924
rect 6436 4868 6440 4924
rect 6376 4864 6440 4868
rect 6456 4924 6520 4928
rect 6456 4868 6460 4924
rect 6460 4868 6516 4924
rect 6516 4868 6520 4924
rect 6456 4864 6520 4868
rect 11480 4924 11544 4928
rect 11480 4868 11484 4924
rect 11484 4868 11540 4924
rect 11540 4868 11544 4924
rect 11480 4864 11544 4868
rect 11560 4924 11624 4928
rect 11560 4868 11564 4924
rect 11564 4868 11620 4924
rect 11620 4868 11624 4924
rect 11560 4864 11624 4868
rect 11640 4924 11704 4928
rect 11640 4868 11644 4924
rect 11644 4868 11700 4924
rect 11700 4868 11704 4924
rect 11640 4864 11704 4868
rect 11720 4924 11784 4928
rect 11720 4868 11724 4924
rect 11724 4868 11780 4924
rect 11780 4868 11784 4924
rect 11720 4864 11784 4868
rect 3584 4380 3648 4384
rect 3584 4324 3588 4380
rect 3588 4324 3644 4380
rect 3644 4324 3648 4380
rect 3584 4320 3648 4324
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 8848 4380 8912 4384
rect 8848 4324 8852 4380
rect 8852 4324 8908 4380
rect 8908 4324 8912 4380
rect 8848 4320 8912 4324
rect 8928 4380 8992 4384
rect 8928 4324 8932 4380
rect 8932 4324 8988 4380
rect 8988 4324 8992 4380
rect 8928 4320 8992 4324
rect 9008 4380 9072 4384
rect 9008 4324 9012 4380
rect 9012 4324 9068 4380
rect 9068 4324 9072 4380
rect 9008 4320 9072 4324
rect 9088 4380 9152 4384
rect 9088 4324 9092 4380
rect 9092 4324 9148 4380
rect 9148 4324 9152 4380
rect 9088 4320 9152 4324
rect 14112 4380 14176 4384
rect 14112 4324 14116 4380
rect 14116 4324 14172 4380
rect 14172 4324 14176 4380
rect 14112 4320 14176 4324
rect 14192 4380 14256 4384
rect 14192 4324 14196 4380
rect 14196 4324 14252 4380
rect 14252 4324 14256 4380
rect 14192 4320 14256 4324
rect 14272 4380 14336 4384
rect 14272 4324 14276 4380
rect 14276 4324 14332 4380
rect 14332 4324 14336 4380
rect 14272 4320 14336 4324
rect 14352 4380 14416 4384
rect 14352 4324 14356 4380
rect 14356 4324 14412 4380
rect 14412 4324 14416 4380
rect 14352 4320 14416 4324
rect 6216 3836 6280 3840
rect 6216 3780 6220 3836
rect 6220 3780 6276 3836
rect 6276 3780 6280 3836
rect 6216 3776 6280 3780
rect 6296 3836 6360 3840
rect 6296 3780 6300 3836
rect 6300 3780 6356 3836
rect 6356 3780 6360 3836
rect 6296 3776 6360 3780
rect 6376 3836 6440 3840
rect 6376 3780 6380 3836
rect 6380 3780 6436 3836
rect 6436 3780 6440 3836
rect 6376 3776 6440 3780
rect 6456 3836 6520 3840
rect 6456 3780 6460 3836
rect 6460 3780 6516 3836
rect 6516 3780 6520 3836
rect 6456 3776 6520 3780
rect 11480 3836 11544 3840
rect 11480 3780 11484 3836
rect 11484 3780 11540 3836
rect 11540 3780 11544 3836
rect 11480 3776 11544 3780
rect 11560 3836 11624 3840
rect 11560 3780 11564 3836
rect 11564 3780 11620 3836
rect 11620 3780 11624 3836
rect 11560 3776 11624 3780
rect 11640 3836 11704 3840
rect 11640 3780 11644 3836
rect 11644 3780 11700 3836
rect 11700 3780 11704 3836
rect 11640 3776 11704 3780
rect 11720 3836 11784 3840
rect 11720 3780 11724 3836
rect 11724 3780 11780 3836
rect 11780 3780 11784 3836
rect 11720 3776 11784 3780
rect 3584 3292 3648 3296
rect 3584 3236 3588 3292
rect 3588 3236 3644 3292
rect 3644 3236 3648 3292
rect 3584 3232 3648 3236
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 8848 3292 8912 3296
rect 8848 3236 8852 3292
rect 8852 3236 8908 3292
rect 8908 3236 8912 3292
rect 8848 3232 8912 3236
rect 8928 3292 8992 3296
rect 8928 3236 8932 3292
rect 8932 3236 8988 3292
rect 8988 3236 8992 3292
rect 8928 3232 8992 3236
rect 9008 3292 9072 3296
rect 9008 3236 9012 3292
rect 9012 3236 9068 3292
rect 9068 3236 9072 3292
rect 9008 3232 9072 3236
rect 9088 3292 9152 3296
rect 9088 3236 9092 3292
rect 9092 3236 9148 3292
rect 9148 3236 9152 3292
rect 9088 3232 9152 3236
rect 14112 3292 14176 3296
rect 14112 3236 14116 3292
rect 14116 3236 14172 3292
rect 14172 3236 14176 3292
rect 14112 3232 14176 3236
rect 14192 3292 14256 3296
rect 14192 3236 14196 3292
rect 14196 3236 14252 3292
rect 14252 3236 14256 3292
rect 14192 3232 14256 3236
rect 14272 3292 14336 3296
rect 14272 3236 14276 3292
rect 14276 3236 14332 3292
rect 14332 3236 14336 3292
rect 14272 3232 14336 3236
rect 14352 3292 14416 3296
rect 14352 3236 14356 3292
rect 14356 3236 14412 3292
rect 14412 3236 14416 3292
rect 14352 3232 14416 3236
rect 6216 2748 6280 2752
rect 6216 2692 6220 2748
rect 6220 2692 6276 2748
rect 6276 2692 6280 2748
rect 6216 2688 6280 2692
rect 6296 2748 6360 2752
rect 6296 2692 6300 2748
rect 6300 2692 6356 2748
rect 6356 2692 6360 2748
rect 6296 2688 6360 2692
rect 6376 2748 6440 2752
rect 6376 2692 6380 2748
rect 6380 2692 6436 2748
rect 6436 2692 6440 2748
rect 6376 2688 6440 2692
rect 6456 2748 6520 2752
rect 6456 2692 6460 2748
rect 6460 2692 6516 2748
rect 6516 2692 6520 2748
rect 6456 2688 6520 2692
rect 11480 2748 11544 2752
rect 11480 2692 11484 2748
rect 11484 2692 11540 2748
rect 11540 2692 11544 2748
rect 11480 2688 11544 2692
rect 11560 2748 11624 2752
rect 11560 2692 11564 2748
rect 11564 2692 11620 2748
rect 11620 2692 11624 2748
rect 11560 2688 11624 2692
rect 11640 2748 11704 2752
rect 11640 2692 11644 2748
rect 11644 2692 11700 2748
rect 11700 2692 11704 2748
rect 11640 2688 11704 2692
rect 11720 2748 11784 2752
rect 11720 2692 11724 2748
rect 11724 2692 11780 2748
rect 11780 2692 11784 2748
rect 11720 2688 11784 2692
rect 3584 2204 3648 2208
rect 3584 2148 3588 2204
rect 3588 2148 3644 2204
rect 3644 2148 3648 2204
rect 3584 2144 3648 2148
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 8848 2204 8912 2208
rect 8848 2148 8852 2204
rect 8852 2148 8908 2204
rect 8908 2148 8912 2204
rect 8848 2144 8912 2148
rect 8928 2204 8992 2208
rect 8928 2148 8932 2204
rect 8932 2148 8988 2204
rect 8988 2148 8992 2204
rect 8928 2144 8992 2148
rect 9008 2204 9072 2208
rect 9008 2148 9012 2204
rect 9012 2148 9068 2204
rect 9068 2148 9072 2204
rect 9008 2144 9072 2148
rect 9088 2204 9152 2208
rect 9088 2148 9092 2204
rect 9092 2148 9148 2204
rect 9148 2148 9152 2204
rect 9088 2144 9152 2148
rect 14112 2204 14176 2208
rect 14112 2148 14116 2204
rect 14116 2148 14172 2204
rect 14172 2148 14176 2204
rect 14112 2144 14176 2148
rect 14192 2204 14256 2208
rect 14192 2148 14196 2204
rect 14196 2148 14252 2204
rect 14252 2148 14256 2204
rect 14192 2144 14256 2148
rect 14272 2204 14336 2208
rect 14272 2148 14276 2204
rect 14276 2148 14332 2204
rect 14332 2148 14336 2204
rect 14272 2144 14336 2148
rect 14352 2204 14416 2208
rect 14352 2148 14356 2204
rect 14356 2148 14412 2204
rect 14412 2148 14416 2204
rect 14352 2144 14416 2148
<< metal4 >>
rect 3576 14176 3896 14736
rect 3576 14112 3584 14176
rect 3648 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3896 14176
rect 3576 13088 3896 14112
rect 3576 13024 3584 13088
rect 3648 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3896 13088
rect 3576 12000 3896 13024
rect 3576 11936 3584 12000
rect 3648 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3896 12000
rect 3576 10912 3896 11936
rect 3576 10848 3584 10912
rect 3648 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3896 10912
rect 3576 9824 3896 10848
rect 3576 9760 3584 9824
rect 3648 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3896 9824
rect 3576 8736 3896 9760
rect 3576 8672 3584 8736
rect 3648 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3896 8736
rect 3576 7648 3896 8672
rect 3576 7584 3584 7648
rect 3648 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3896 7648
rect 3576 6560 3896 7584
rect 3576 6496 3584 6560
rect 3648 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3896 6560
rect 3576 5472 3896 6496
rect 3576 5408 3584 5472
rect 3648 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3896 5472
rect 3576 4384 3896 5408
rect 3576 4320 3584 4384
rect 3648 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3896 4384
rect 3576 3296 3896 4320
rect 3576 3232 3584 3296
rect 3648 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3896 3296
rect 3576 2208 3896 3232
rect 3576 2144 3584 2208
rect 3648 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3896 2208
rect 3576 2128 3896 2144
rect 6208 14720 6528 14736
rect 6208 14656 6216 14720
rect 6280 14656 6296 14720
rect 6360 14656 6376 14720
rect 6440 14656 6456 14720
rect 6520 14656 6528 14720
rect 6208 13632 6528 14656
rect 6208 13568 6216 13632
rect 6280 13568 6296 13632
rect 6360 13568 6376 13632
rect 6440 13568 6456 13632
rect 6520 13568 6528 13632
rect 6208 12544 6528 13568
rect 6208 12480 6216 12544
rect 6280 12480 6296 12544
rect 6360 12480 6376 12544
rect 6440 12480 6456 12544
rect 6520 12480 6528 12544
rect 6208 11456 6528 12480
rect 6208 11392 6216 11456
rect 6280 11392 6296 11456
rect 6360 11392 6376 11456
rect 6440 11392 6456 11456
rect 6520 11392 6528 11456
rect 6208 10368 6528 11392
rect 6208 10304 6216 10368
rect 6280 10304 6296 10368
rect 6360 10304 6376 10368
rect 6440 10304 6456 10368
rect 6520 10304 6528 10368
rect 6208 9280 6528 10304
rect 6208 9216 6216 9280
rect 6280 9216 6296 9280
rect 6360 9216 6376 9280
rect 6440 9216 6456 9280
rect 6520 9216 6528 9280
rect 6208 8192 6528 9216
rect 6208 8128 6216 8192
rect 6280 8128 6296 8192
rect 6360 8128 6376 8192
rect 6440 8128 6456 8192
rect 6520 8128 6528 8192
rect 6208 7104 6528 8128
rect 6208 7040 6216 7104
rect 6280 7040 6296 7104
rect 6360 7040 6376 7104
rect 6440 7040 6456 7104
rect 6520 7040 6528 7104
rect 6208 6016 6528 7040
rect 6208 5952 6216 6016
rect 6280 5952 6296 6016
rect 6360 5952 6376 6016
rect 6440 5952 6456 6016
rect 6520 5952 6528 6016
rect 6208 4928 6528 5952
rect 6208 4864 6216 4928
rect 6280 4864 6296 4928
rect 6360 4864 6376 4928
rect 6440 4864 6456 4928
rect 6520 4864 6528 4928
rect 6208 3840 6528 4864
rect 6208 3776 6216 3840
rect 6280 3776 6296 3840
rect 6360 3776 6376 3840
rect 6440 3776 6456 3840
rect 6520 3776 6528 3840
rect 6208 2752 6528 3776
rect 6208 2688 6216 2752
rect 6280 2688 6296 2752
rect 6360 2688 6376 2752
rect 6440 2688 6456 2752
rect 6520 2688 6528 2752
rect 6208 2128 6528 2688
rect 8840 14176 9160 14736
rect 8840 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9160 14176
rect 8840 13088 9160 14112
rect 8840 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9160 13088
rect 8840 12000 9160 13024
rect 8840 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9160 12000
rect 8840 10912 9160 11936
rect 8840 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9160 10912
rect 8840 9824 9160 10848
rect 8840 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9160 9824
rect 8840 8736 9160 9760
rect 8840 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9160 8736
rect 8840 7648 9160 8672
rect 8840 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9160 7648
rect 8840 6560 9160 7584
rect 8840 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9160 6560
rect 8840 5472 9160 6496
rect 8840 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9160 5472
rect 8840 4384 9160 5408
rect 8840 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9160 4384
rect 8840 3296 9160 4320
rect 8840 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9160 3296
rect 8840 2208 9160 3232
rect 8840 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9160 2208
rect 8840 2128 9160 2144
rect 11472 14720 11792 14736
rect 11472 14656 11480 14720
rect 11544 14656 11560 14720
rect 11624 14656 11640 14720
rect 11704 14656 11720 14720
rect 11784 14656 11792 14720
rect 11472 13632 11792 14656
rect 11472 13568 11480 13632
rect 11544 13568 11560 13632
rect 11624 13568 11640 13632
rect 11704 13568 11720 13632
rect 11784 13568 11792 13632
rect 11472 12544 11792 13568
rect 11472 12480 11480 12544
rect 11544 12480 11560 12544
rect 11624 12480 11640 12544
rect 11704 12480 11720 12544
rect 11784 12480 11792 12544
rect 11472 11456 11792 12480
rect 11472 11392 11480 11456
rect 11544 11392 11560 11456
rect 11624 11392 11640 11456
rect 11704 11392 11720 11456
rect 11784 11392 11792 11456
rect 11472 10368 11792 11392
rect 11472 10304 11480 10368
rect 11544 10304 11560 10368
rect 11624 10304 11640 10368
rect 11704 10304 11720 10368
rect 11784 10304 11792 10368
rect 11472 9280 11792 10304
rect 11472 9216 11480 9280
rect 11544 9216 11560 9280
rect 11624 9216 11640 9280
rect 11704 9216 11720 9280
rect 11784 9216 11792 9280
rect 11472 8192 11792 9216
rect 11472 8128 11480 8192
rect 11544 8128 11560 8192
rect 11624 8128 11640 8192
rect 11704 8128 11720 8192
rect 11784 8128 11792 8192
rect 11472 7104 11792 8128
rect 11472 7040 11480 7104
rect 11544 7040 11560 7104
rect 11624 7040 11640 7104
rect 11704 7040 11720 7104
rect 11784 7040 11792 7104
rect 11472 6016 11792 7040
rect 11472 5952 11480 6016
rect 11544 5952 11560 6016
rect 11624 5952 11640 6016
rect 11704 5952 11720 6016
rect 11784 5952 11792 6016
rect 11472 4928 11792 5952
rect 11472 4864 11480 4928
rect 11544 4864 11560 4928
rect 11624 4864 11640 4928
rect 11704 4864 11720 4928
rect 11784 4864 11792 4928
rect 11472 3840 11792 4864
rect 11472 3776 11480 3840
rect 11544 3776 11560 3840
rect 11624 3776 11640 3840
rect 11704 3776 11720 3840
rect 11784 3776 11792 3840
rect 11472 2752 11792 3776
rect 11472 2688 11480 2752
rect 11544 2688 11560 2752
rect 11624 2688 11640 2752
rect 11704 2688 11720 2752
rect 11784 2688 11792 2752
rect 11472 2128 11792 2688
rect 14104 14176 14424 14736
rect 14104 14112 14112 14176
rect 14176 14112 14192 14176
rect 14256 14112 14272 14176
rect 14336 14112 14352 14176
rect 14416 14112 14424 14176
rect 14104 13088 14424 14112
rect 14104 13024 14112 13088
rect 14176 13024 14192 13088
rect 14256 13024 14272 13088
rect 14336 13024 14352 13088
rect 14416 13024 14424 13088
rect 14104 12000 14424 13024
rect 14104 11936 14112 12000
rect 14176 11936 14192 12000
rect 14256 11936 14272 12000
rect 14336 11936 14352 12000
rect 14416 11936 14424 12000
rect 14104 10912 14424 11936
rect 14104 10848 14112 10912
rect 14176 10848 14192 10912
rect 14256 10848 14272 10912
rect 14336 10848 14352 10912
rect 14416 10848 14424 10912
rect 14104 9824 14424 10848
rect 14104 9760 14112 9824
rect 14176 9760 14192 9824
rect 14256 9760 14272 9824
rect 14336 9760 14352 9824
rect 14416 9760 14424 9824
rect 14104 8736 14424 9760
rect 14779 9620 14845 9621
rect 14779 9556 14780 9620
rect 14844 9556 14845 9620
rect 14779 9555 14845 9556
rect 14104 8672 14112 8736
rect 14176 8672 14192 8736
rect 14256 8672 14272 8736
rect 14336 8672 14352 8736
rect 14416 8672 14424 8736
rect 14104 7648 14424 8672
rect 14104 7584 14112 7648
rect 14176 7584 14192 7648
rect 14256 7584 14272 7648
rect 14336 7584 14352 7648
rect 14416 7584 14424 7648
rect 14104 6560 14424 7584
rect 14782 7309 14842 9555
rect 14779 7308 14845 7309
rect 14779 7244 14780 7308
rect 14844 7244 14845 7308
rect 14779 7243 14845 7244
rect 14104 6496 14112 6560
rect 14176 6496 14192 6560
rect 14256 6496 14272 6560
rect 14336 6496 14352 6560
rect 14416 6496 14424 6560
rect 14104 5472 14424 6496
rect 14104 5408 14112 5472
rect 14176 5408 14192 5472
rect 14256 5408 14272 5472
rect 14336 5408 14352 5472
rect 14416 5408 14424 5472
rect 14104 4384 14424 5408
rect 14104 4320 14112 4384
rect 14176 4320 14192 4384
rect 14256 4320 14272 4384
rect 14336 4320 14352 4384
rect 14416 4320 14424 4384
rect 14104 3296 14424 4320
rect 14104 3232 14112 3296
rect 14176 3232 14192 3296
rect 14256 3232 14272 3296
rect 14336 3232 14352 3296
rect 14416 3232 14424 3296
rect 14104 2208 14424 3232
rect 14104 2144 14112 2208
rect 14176 2144 14192 2208
rect 14256 2144 14272 2208
rect 14336 2144 14352 2208
rect 14416 2144 14424 2208
rect 14104 2128 14424 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _29_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1605641404
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1605641404
transform 1 0 2300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1605641404
transform 1 0 1932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1605641404
transform 1 0 2668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_19 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3772 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21
timestamp 1605641404
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1605641404
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_35
timestamp 1605641404
transform 1 0 4324 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_45
timestamp 1605641404
transform 1 0 5244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1605641404
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 8188 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7636 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6992 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_80
timestamp 1605641404
transform 1 0 8464 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1605641404
transform 1 0 7820 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10028 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1605641404
transform 1 0 9660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1605641404
transform 1 0 10580 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110
timestamp 1605641404
transform 1 0 11224 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106
timestamp 1605641404
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11316 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10948 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_116
timestamp 1605641404
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1605641404
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117
timestamp 1605641404
transform 1 0 11868 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1605641404
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137
timestamp 1605641404
transform 1 0 13708 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1605641404
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_133
timestamp 1605641404
transform 1 0 13340 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_141
timestamp 1605641404
transform 1 0 14076 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_146
timestamp 1605641404
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1605641404
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1605641404
transform 1 0 14904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1605641404
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_154
timestamp 1605641404
transform 1 0 15272 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1605641404
transform 1 0 16192 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1605641404
transform 1 0 16192 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1605641404
transform 1 0 15824 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1605641404
transform 1 0 15824 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 16836 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 16836 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1605641404
transform 1 0 2392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_10
timestamp 1605641404
transform 1 0 2024 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_18
timestamp 1605641404
transform 1 0 2760 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1605641404
transform 1 0 3128 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_26
timestamp 1605641404
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1605641404
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_36
timestamp 1605641404
transform 1 0 4416 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5428 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_44
timestamp 1605641404
transform 1 0 5152 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8280 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_63
timestamp 1605641404
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_75
timestamp 1605641404
transform 1 0 8004 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1605641404
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1605641404
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1605641404
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_115
timestamp 1605641404
transform 1 0 11684 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1605641404
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_127
timestamp 1605641404
transform 1 0 12788 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_139
timestamp 1605641404
transform 1 0 13892 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1605641404
transform 1 0 15824 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1605641404
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_154
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1605641404
transform 1 0 16192 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 16836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1605641404
transform 1 0 1564 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2944 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_9
timestamp 1605641404
transform 1 0 1932 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_17
timestamp 1605641404
transform 1 0 2668 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4140 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1605641404
transform 1 0 3772 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_49
timestamp 1605641404
transform 1 0 5612 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_62
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8648 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 7452 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp 1605641404
transform 1 0 7360 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1605641404
transform 1 0 8280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _15_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10488 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1605641404
transform 1 0 10120 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11132 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_105
timestamp 1605641404
transform 1 0 10764 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1605641404
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1605641404
transform 1 0 14352 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_132
timestamp 1605641404
transform 1 0 13248 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1605641404
transform 1 0 15824 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1605641404
transform 1 0 15088 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_148
timestamp 1605641404
transform 1 0 14720 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1605641404
transform 1 0 15456 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1605641404
transform 1 0 16192 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 16836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2116 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1605641404
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_36
timestamp 1605641404
transform 1 0 4416 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5152 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1605641404
transform 1 0 5980 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7728 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_66
timestamp 1605641404
transform 1 0 7176 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_81
timestamp 1605641404
transform 1 0 8556 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1605641404
transform 1 0 9936 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1605641404
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 11132 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12512 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_105
timestamp 1605641404
transform 1 0 10764 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_118
timestamp 1605641404
transform 1 0 11960 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_133
timestamp 1605641404
transform 1 0 13340 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1605641404
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1605641404
transform 1 0 15824 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_154
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1605641404
transform 1 0 16192 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 16836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1932 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_18
timestamp 1605641404
transform 1 0 2760 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4324 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3128 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 1605641404
transform 1 0 3956 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 5520 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1605641404
transform 1 0 5152 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1605641404
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8648 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1605641404
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1605641404
transform 1 0 10488 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12512 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_111
timestamp 1605641404
transform 1 0 11316 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1605641404
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_123
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13708 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_133
timestamp 1605641404
transform 1 0 13340 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1605641404
transform 1 0 15824 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_146
timestamp 1605641404
transform 1 0 14536 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1605641404
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1605641404
transform 1 0 16192 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 16836 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1656 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1564 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1605641404
transform 1 0 2208 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1605641404
transform 1 0 2392 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 2760 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2576 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4416 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4416 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_32
timestamp 1605641404
transform 1 0 4048 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 6348 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_45
timestamp 1605641404
transform 1 0 5244 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_52
timestamp 1605641404
transform 1 0 5888 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1605641404
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _09_
timestamp 1605641404
transform 1 0 7544 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 8740 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8372 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1605641404
transform 1 0 7176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_73
timestamp 1605641404
transform 1 0 7820 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_71
timestamp 1605641404
transform 1 0 7636 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9936 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1605641404
transform 1 0 10120 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1605641404
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1605641404
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_92
timestamp 1605641404
transform 1 0 9568 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11776 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_107
timestamp 1605641404
transform 1 0 10948 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_115
timestamp 1605641404
transform 1 0 11684 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_112
timestamp 1605641404
transform 1 0 11408 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp 1605641404
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 13616 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13984 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_132
timestamp 1605641404
transform 1 0 13248 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1605641404
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1605641404
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1605641404
transform 1 0 15824 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1605641404
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1605641404
transform 1 0 16192 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_152
timestamp 1605641404
transform 1 0 15088 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1605641404
transform 1 0 16192 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 16836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 16836 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2116 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1605641404
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 4784 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 1605641404
transform 1 0 4416 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6256 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5060 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_52
timestamp 1605641404
transform 1 0 5888 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8096 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_72
timestamp 1605641404
transform 1 0 7728 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _14_
timestamp 1605641404
transform 1 0 10120 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1605641404
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 1605641404
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_101
timestamp 1605641404
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10764 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_121
timestamp 1605641404
transform 1 0 12236 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1605641404
transform 1 0 14444 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1605641404
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_140
timestamp 1605641404
transform 1 0 13984 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_144
timestamp 1605641404
transform 1 0 14352 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1605641404
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1605641404
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 16836 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_167
timestamp 1605641404
transform 1 0 16468 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1605641404
transform 1 0 1564 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2484 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_9
timestamp 1605641404
transform 1 0 1932 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_24
timestamp 1605641404
transform 1 0 3312 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1605641404
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1605641404
transform 1 0 6072 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_50
timestamp 1605641404
transform 1 0 5704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1605641404
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 8096 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_9_71
timestamp 1605641404
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_75
timestamp 1605641404
transform 1 0 8004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9936 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11408 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1605641404
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1605641404
transform 1 0 14260 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1605641404
transform 1 0 13892 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1605641404
transform 1 0 15824 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_152
timestamp 1605641404
transform 1 0 15088 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1605641404
transform 1 0 16192 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 16836 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1605641404
transform 1 0 2760 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1564 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1605641404
transform 1 0 2392 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1605641404
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1605641404
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1605641404
transform 1 0 5704 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 6716 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 6440 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1605641404
transform 1 0 5336 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_54
timestamp 1605641404
transform 1 0 6072 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8372 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_70
timestamp 1605641404
transform 1 0 7544 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_78
timestamp 1605641404
transform 1 0 8280 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9752 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1605641404
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1605641404
transform 1 0 10580 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10948 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12144 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_116
timestamp 1605641404
transform 1 0 11776 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13340 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_129
timestamp 1605641404
transform 1 0 12972 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_142
timestamp 1605641404
transform 1 0 14168 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1605641404
transform 1 0 14536 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1605641404
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1605641404
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 16836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_167
timestamp 1605641404
transform 1 0 16468 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2116 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1605641404
transform 1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 3956 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1605641404
transform 1 0 3588 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1605641404
transform 1 0 5796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_47
timestamp 1605641404
transform 1 0 5428 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_55
timestamp 1605641404
transform 1 0 6164 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8004 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1605641404
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9844 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1605641404
transform 1 0 9476 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_104
timestamp 1605641404
transform 1 0 10672 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11040 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1605641404
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1605641404
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13984 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12788 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 1605641404
transform 1 0 13616 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1605641404
transform 1 0 15824 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_156
timestamp 1605641404
transform 1 0 15456 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1605641404
transform 1 0 16192 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 16836 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2024 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1605641404
transform 1 0 1656 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_19
timestamp 1605641404
transform 1 0 2852 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1605641404
transform 1 0 3220 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1605641404
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_36
timestamp 1605641404
transform 1 0 4416 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5060 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_42
timestamp 1605641404
transform 1 0 4968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_59
timestamp 1605641404
transform 1 0 6532 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6900 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8096 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_72
timestamp 1605641404
transform 1 0 7728 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9936 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1605641404
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1605641404
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_93
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11132 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_105
timestamp 1605641404
transform 1 0 10764 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_125
timestamp 1605641404
transform 1 0 12604 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1605641404
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12972 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_12_138
timestamp 1605641404
transform 1 0 13800 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_144
timestamp 1605641404
transform 1 0 14352 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1605641404
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1605641404
transform 1 0 16100 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1605641404
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1605641404
transform 1 0 1932 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1605641404
transform 1 0 1932 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1605641404
transform 1 0 1564 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_19
timestamp 1605641404
transform 1 0 2852 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1605641404
transform 1 0 2300 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2024 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3312 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4600 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_23
timestamp 1605641404
transform 1 0 3220 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_40
timestamp 1605641404
transform 1 0 4784 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_22
timestamp 1605641404
transform 1 0 3128 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1605641404
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5520 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 5152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_47
timestamp 1605641404
transform 1 0 5428 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1605641404
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1605641404
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8648 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 8372 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7176 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1605641404
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_75
timestamp 1605641404
transform 1 0 8004 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9752 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10212 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_91
timestamp 1605641404
transform 1 0 9476 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1605641404
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1605641404
transform 1 0 11776 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 11408 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1605641404
transform 1 0 11040 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_115
timestamp 1605641404
transform 1 0 11684 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1605641404
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_110
timestamp 1605641404
transform 1 0 11224 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_125
timestamp 1605641404
transform 1 0 12604 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1605641404
transform 1 0 13340 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13984 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_139
timestamp 1605641404
transform 1 0 13892 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1605641404
transform 1 0 13616 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1605641404
transform 1 0 14628 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15364 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15364 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1605641404
transform 1 0 14996 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1605641404
transform 1 0 16192 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1605641404
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1605641404
transform 1 0 16192 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 16836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2852 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1656 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1605641404
transform 1 0 2484 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1605641404
transform 1 0 4692 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_35
timestamp 1605641404
transform 1 0 4324 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_48
timestamp 1605641404
transform 1 0 5520 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1605641404
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8648 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7268 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1605641404
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_76
timestamp 1605641404
transform 1 0 8096 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10488 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_98
timestamp 1605641404
transform 1 0 10120 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1605641404
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14168 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12880 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1605641404
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_137
timestamp 1605641404
transform 1 0 13708 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_141
timestamp 1605641404
transform 1 0 14076 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1605641404
transform 1 0 15640 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1605641404
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 16836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1932 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 4508 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_25
timestamp 1605641404
transform 1 0 3404 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1605641404
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5796 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_46
timestamp 1605641404
transform 1 0 5336 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_50
timestamp 1605641404
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 7728 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1605641404
transform 1 0 7268 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_71
timestamp 1605641404
transform 1 0 7636 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1605641404
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1605641404
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_117
timestamp 1605641404
transform 1 0 11868 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_125
timestamp 1605641404
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12880 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_144
timestamp 1605641404
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1605641404
transform 1 0 15364 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1605641404
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_164
timestamp 1605641404
transform 1 0 16192 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 16836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1932 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_18
timestamp 1605641404
transform 1 0 2760 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1605641404
transform 1 0 3128 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 3956 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_26
timestamp 1605641404
transform 1 0 3496 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_30
timestamp 1605641404
transform 1 0 3864 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_40
timestamp 1605641404
transform 1 0 4784 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _12_
timestamp 1605641404
transform 1 0 5152 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_47
timestamp 1605641404
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 7360 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8556 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_77
timestamp 1605641404
transform 1 0 8188 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_90
timestamp 1605641404
transform 1 0 9384 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_102
timestamp 1605641404
transform 1 0 10488 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_114
timestamp 1605641404
transform 1 0 11592 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_132
timestamp 1605641404
transform 1 0 13248 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_144
timestamp 1605641404
transform 1 0 14352 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 14904 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1605641404
transform 1 0 15732 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 16836 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1605641404
transform 1 0 16468 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1656 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1605641404
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1605641404
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1605641404
transform 1 0 4876 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 6256 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_53
timestamp 1605641404
transform 1 0 5980 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _13_
timestamp 1605641404
transform 1 0 8648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 7452 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_65
timestamp 1605641404
transform 1 0 7084 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_78
timestamp 1605641404
transform 1 0 8280 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1605641404
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1605641404
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1605641404
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1605641404
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1605641404
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1605641404
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1605641404
transform 1 0 15824 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_154
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_164
timestamp 1605641404
transform 1 0 16192 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 16836 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1605641404
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1605641404
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1605641404
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1605641404
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1605641404
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1605641404
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1605641404
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1605641404
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1605641404
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1605641404
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1605641404
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1605641404
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1605641404
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1605641404
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1605641404
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1605641404
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1605641404
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1605641404
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1605641404
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1605641404
transform 1 0 15732 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1605641404
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 16836 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1605641404
transform 1 0 16468 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1605641404
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1605641404
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1605641404
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1605641404
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1605641404
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1605641404
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1605641404
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1605641404
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1605641404
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1605641404
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1605641404
transform 1 0 15732 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 16836 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1605641404
transform 1 0 16468 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1605641404
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1605641404
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1605641404
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1605641404
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1605641404
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1605641404
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1605641404
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1605641404
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1605641404
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1605641404
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1605641404
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1605641404
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1605641404
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1605641404
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 16836 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 754 0 810 480 6 bottom_grid_pin_0_
port 0 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 bottom_grid_pin_10_
port 1 nsew default tristate
rlabel metal2 s 9770 0 9826 480 6 bottom_grid_pin_12_
port 2 nsew default tristate
rlabel metal2 s 11242 0 11298 480 6 bottom_grid_pin_14_
port 3 nsew default tristate
rlabel metal2 s 12714 0 12770 480 6 bottom_grid_pin_16_
port 4 nsew default tristate
rlabel metal2 s 2226 0 2282 480 6 bottom_grid_pin_2_
port 5 nsew default tristate
rlabel metal2 s 3698 0 3754 480 6 bottom_grid_pin_4_
port 6 nsew default tristate
rlabel metal2 s 5262 0 5318 480 6 bottom_grid_pin_6_
port 7 nsew default tristate
rlabel metal2 s 6734 0 6790 480 6 bottom_grid_pin_8_
port 8 nsew default tristate
rlabel metal2 s 14278 0 14334 480 6 ccff_head
port 9 nsew default input
rlabel metal2 s 15750 0 15806 480 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 14152 480 14272 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 144 480 264 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 5176 480 5296 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 5992 480 6112 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 6400 480 6520 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 6944 480 7064 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 7760 480 7880 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 8168 480 8288 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 552 480 672 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 960 480 1080 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 1776 480 1896 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 3544 480 3664 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal3 s 17520 8576 18000 8696 6 chanx_right_in[0]
port 51 nsew default input
rlabel metal3 s 17520 12792 18000 12912 6 chanx_right_in[10]
port 52 nsew default input
rlabel metal3 s 17520 13200 18000 13320 6 chanx_right_in[11]
port 53 nsew default input
rlabel metal3 s 17520 13744 18000 13864 6 chanx_right_in[12]
port 54 nsew default input
rlabel metal3 s 17520 14152 18000 14272 6 chanx_right_in[13]
port 55 nsew default input
rlabel metal3 s 17520 14560 18000 14680 6 chanx_right_in[14]
port 56 nsew default input
rlabel metal3 s 17520 14968 18000 15088 6 chanx_right_in[15]
port 57 nsew default input
rlabel metal3 s 17520 15376 18000 15496 6 chanx_right_in[16]
port 58 nsew default input
rlabel metal3 s 17520 15784 18000 15904 6 chanx_right_in[17]
port 59 nsew default input
rlabel metal3 s 17520 16192 18000 16312 6 chanx_right_in[18]
port 60 nsew default input
rlabel metal3 s 17520 16600 18000 16720 6 chanx_right_in[19]
port 61 nsew default input
rlabel metal3 s 17520 8984 18000 9104 6 chanx_right_in[1]
port 62 nsew default input
rlabel metal3 s 17520 9392 18000 9512 6 chanx_right_in[2]
port 63 nsew default input
rlabel metal3 s 17520 9800 18000 9920 6 chanx_right_in[3]
port 64 nsew default input
rlabel metal3 s 17520 10344 18000 10464 6 chanx_right_in[4]
port 65 nsew default input
rlabel metal3 s 17520 10752 18000 10872 6 chanx_right_in[5]
port 66 nsew default input
rlabel metal3 s 17520 11160 18000 11280 6 chanx_right_in[6]
port 67 nsew default input
rlabel metal3 s 17520 11568 18000 11688 6 chanx_right_in[7]
port 68 nsew default input
rlabel metal3 s 17520 11976 18000 12096 6 chanx_right_in[8]
port 69 nsew default input
rlabel metal3 s 17520 12384 18000 12504 6 chanx_right_in[9]
port 70 nsew default input
rlabel metal3 s 17520 144 18000 264 6 chanx_right_out[0]
port 71 nsew default tristate
rlabel metal3 s 17520 4360 18000 4480 6 chanx_right_out[10]
port 72 nsew default tristate
rlabel metal3 s 17520 4768 18000 4888 6 chanx_right_out[11]
port 73 nsew default tristate
rlabel metal3 s 17520 5176 18000 5296 6 chanx_right_out[12]
port 74 nsew default tristate
rlabel metal3 s 17520 5584 18000 5704 6 chanx_right_out[13]
port 75 nsew default tristate
rlabel metal3 s 17520 5992 18000 6112 6 chanx_right_out[14]
port 76 nsew default tristate
rlabel metal3 s 17520 6400 18000 6520 6 chanx_right_out[15]
port 77 nsew default tristate
rlabel metal3 s 17520 6944 18000 7064 6 chanx_right_out[16]
port 78 nsew default tristate
rlabel metal3 s 17520 7352 18000 7472 6 chanx_right_out[17]
port 79 nsew default tristate
rlabel metal3 s 17520 7760 18000 7880 6 chanx_right_out[18]
port 80 nsew default tristate
rlabel metal3 s 17520 8168 18000 8288 6 chanx_right_out[19]
port 81 nsew default tristate
rlabel metal3 s 17520 552 18000 672 6 chanx_right_out[1]
port 82 nsew default tristate
rlabel metal3 s 17520 960 18000 1080 6 chanx_right_out[2]
port 83 nsew default tristate
rlabel metal3 s 17520 1368 18000 1488 6 chanx_right_out[3]
port 84 nsew default tristate
rlabel metal3 s 17520 1776 18000 1896 6 chanx_right_out[4]
port 85 nsew default tristate
rlabel metal3 s 17520 2184 18000 2304 6 chanx_right_out[5]
port 86 nsew default tristate
rlabel metal3 s 17520 2592 18000 2712 6 chanx_right_out[6]
port 87 nsew default tristate
rlabel metal3 s 17520 3000 18000 3120 6 chanx_right_out[7]
port 88 nsew default tristate
rlabel metal3 s 17520 3544 18000 3664 6 chanx_right_out[8]
port 89 nsew default tristate
rlabel metal3 s 17520 3952 18000 4072 6 chanx_right_out[9]
port 90 nsew default tristate
rlabel metal2 s 17222 0 17278 480 6 prog_clk
port 91 nsew default input
rlabel metal4 s 3576 2128 3896 14736 6 VPWR
port 92 nsew default input
rlabel metal4 s 6208 2128 6528 14736 6 VGND
port 93 nsew default input
<< properties >>
string FIXED_BBOX 0 0 18000 16720
<< end >>
